`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dnggK926ZO8IcqDoMNn+02G/VftJbxi0F35zAh8yZfVxgvLF2b9aq4w4oUnKHq1lHa2cMYZaw85x
LCwpXay1TA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fNzeM8DWHmNDwcUo6c5l9AxoHKSaL7c/3jnlfXX4MgZWXzpwiBCrJ+UlRxrtebikqwNHjIj0BVFb
eZzTL+Nck01cnRQytXx4bE5DiOcgGM46HcWWq1+WNbBhhh8wjiboABJ5Ns+MiyeVzpRsmBA+DTYy
c+mm/OjcjxFm34kX54c=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RkMb7zse1PBAWAvneoYBnbNlOe7unHd0UcjwFZDPkI//0l3t18dSfFuJ2AyTKpwvezEwVfSYRg3o
5+zQEyt7OoGwOGmwuZNPEISxdETPjGiil7p49FM/V9Zz5RHLLjBfTHb/9p8diL0/rptYvIcMPUJC
sdHa5DXZq1PDofchPNzFv/4XFsWwBx0JyWD+uEgBlwypBWHDXSMltZgKPw+DI6/bv+/bs0/jet0G
08DVjR28jGc4/nvG1ka0w8kPoX4mOmUHesCw0t1UM2f7wMYKPvP2v4kUN83QLfxu8oFhVkBvpTZ+
ZgR3m5c98hnLqR1ELNl3leXUXGeOhZOd7Jtd8A==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QMpmYn52STXtmI441q0X39y9uJo4exAhQ3jx+SNYPflkVOl1MveRn1gXPzqdob54xfXhwhCF68PK
ZQrfJoncfQ2fYiWgrK9Mlir+6WafwY7iZYhM1s2tbcuecSjZ0+LDhRFXLINDDfgdFAer/LSCPwm1
51RQSi1IcaQm+JBZxoLM5kHYps06S9EtDDR4loRqs2tKUvZ3hpRx5e7oopOvJGp6NHUN9kgxjulG
uwJem/YUHaRAOLD3/T66P7EmVL/SQhf5pMVEVykKdBEhkwTBL6z5cuIaoWGNWk5vxCJDvnKO/yHt
TtZZbWtCAumd2RegAsh/3W4fwTg5hdCybcWeFw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CCDLl4cjWbLLcg11gegPc0SGUcgD3JPkyZAuyEptVv9XiPNtW5F/O4GcBzSzCoN6pyyXv59XuObw
i1OUF/+HaFwvF5VmRSx77zwSb2+J5wiUyHQ0z+iy4bAkcwPXm9BVVyMgUdbPbDDiwy21uG0SkXXZ
IMxe4ECqHhj2SNNrQOg=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bBvfOsxVjqQTTUggJgqnrIOMWiwIzWZm9Nihn5GUxU3VJ1/nNbalfLlJuiKrjB/Nz5lhAdMOqfTR
j4cGiPAOwS505ay+Ndorz5qP8Iycz/eOGawswkyfhFvF1ThSZi4fG0olLXse0OH881O15jB9P1EL
aj+Io7JkWusXBUvJbt9fesa8/BQaps+T3z+h77lYf1Hj0jKb7GR0Tvw6PI0HKxsp+H6nz4xXHOhR
nsH3hCDi+NYH8BosNl8MVb9J1AzsSwWKG7Mao11u8tWEXUFbV5arLIn/KFB0G0+a/9fWEVpegZFG
7fazSwNtOUVPwr7b1lBno7BufrkBEZ4jqVRGEw==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1QtT/UxSbh7J2IbT6pU2xP/X69UpEsBQVMSThGJZsmmMjz/xFRkDtv1MU+OV+AZo6h0HriEmBt9y
xlAbTNnMs473sHd7vy8KVbaFQbhZTgGDAQQTdWI8YZj/HZBm87QBxymMNfiSDEY7XNicK3Et2/yg
LKhXtLjTkAZk45jpQUOW79WZOHd8DIP3gVN+WKLlr/zGgzbiZTmThT7wNfoN/k5NTMvpIJNjzZBM
yPJFHrsxLCwtBOKCysJb/0HoKfn2xSPUjFPyYg5sqYbVY2zDoWkEeC4QvSLORykugz4zCa3yp+Qo
4r7LA3iUaNm4Xg0z8QABRzqSHz4FFw2sk9OjOw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kPBKsVI7qsOjWj0HTggE0xmdxIkfJDa4wXhEV4AVVS3YT6Tl/1vmJj0BlvvbiOc4nQnsOSoKksEw
9h6xCQOeuo1KrjK989GOmEl1TpXJS9VIFCl57z5Wj4DBKr5SK3u/CsrASXOPPPDZsNbGWiuil+xt
F57TThhVuUpTCLoDQuk8KbFpHTD7ZZVCtDHV62ZJLg46oeMYNOkDyC1SnCwwdotw49yEY0aKSPdS
5lzyGSKgU+vPVh9lWu4hpXxd2MQu0KidKXVenKkrMxSbFSenQ12Qwczt3v6mOzMDt1uJ/fCPz4E8
pSxKrrBWIhwwkYYKB8nnOrlZ6hgNdal+DKOX7Q==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UR6lAh2Q7tK/eUnnykUjcFUUsFV6R/XxvauK/Zyq6yFXdOd9auB69qwEkBZYf70DtbQnZaW5uGPm
q6KHj6roRBdl/xA+zyufOcTVcJitoX8Yydx6YQXY6dpDZsQCbO6nCNDnhDVr1buG3jW5bsCL0L6h
jYUepOy62qbeU0HUkjTdCryRbHYaqTPRoNfXf4pwSYKliycHbuG7YVqMSp4iNkZkzIawYv2b7Qlr
+wR+XdDMIkZXewLl4sbofiFWshI84MSj0fHwgXL+1ORvqfB73sit3KNfYhxViYqukM/mnHq2MxhF
BKuMq+AFI+yrfdhF09KyzrTiAmfNCQfg6n9U8A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1817872)
`protect data_block
uyKRM+FkuNi3lfCsYUlZAV2fHNw2pS9hmB2uvMG49SJnqxB2oAUUAkiHXcoQgyEkpd4EvFiAy8u5
dNYelPo5eax+sy6FDWJPDlTvjWVu2ag3i8mkm+4EurMLe2zwYAGw0X2Rfslytf6Qz+ipoUFb7nXf
j8dR6zTlpsdY8usmrTvy99Z/MniHiCC9WZdNu6ItKt4fyv8IH09cf1Pw0aOloeQ/OINRa4kLyEOP
cPzSbqmLK9JDZwwmd6NoAkLJRFywP4HajZrSzFh/6vcqtmE5l/kCYhA2D/XDmnjEZohiU0+8wJNR
pDygnsbrsWx44q98HFFgLrkqkdPzlKl35BfVHqPJoEtePElVxhsVAlZEDjLKrV4xF2RtrtI8HR7D
gcR2P2Ti93nvHhZkVca+alFR36J/3zeprzedgfJlI/cXT55vlh5949PGClVGgSN4jIqYH0lUyhgM
iwM4Je8jHmYKcJiZscy1RvxdXHK1sTkuk6jfXXipSbfEctqIh72dmJ1ElJA1hp7W9fzi3YoNpZ8Z
In8j4g5MkVOATt4RTfDoQaNvFJhwv6C3NhWWQ3XJCBRq4iqtBf7qDRJPA4+wuJwDLcQEJJvy0cXw
j1k+mKqhuyxk2shcWw0Dok6tjyHHxSbMK+2Tqd4NSv5J0U1Bm65OttOVpBs5IVoaCKRRdrUkiv5n
SFPQpc99ZfnRsRUbik9fUXJha1ZLzXVmA2jXQpAHWdxYqy4Ubc9Cw7l2MxfQ/2cjWyuNoqQ3lHEy
iEvoFbQGih8zY7BS6MgjaNHiYpJ1/FqwBHguDdeRYjkU4iXzfn/0kAONAbtEdECotnzLyaHY26/A
vpM1OAi2kYufmF2CU/a/7XeS4ngw+I6pynSpFteb3KCtFjiGfOgLMLXr0DhkA1piFfj2TX18kFVY
PP8wU7b1oKutMZbrTRMRa/5qef9szmuNoRCsF5RXBW+WZr05Z9grLE6XnC8B09hS8lfgFUsKmw3s
AAQw1RKgmIkCXCLG1RKC6k1PkzUqZgW3x/lZC7tj/qO7wh2mjjLgGkG7YbXw52x82yQuDGasWVov
MRo+k37KHwxLPMa9aNKP1i8GcNVdU3wpJe6zvGgLq6O+LYZDxtVfAnaGC0IGT3OXyxGloIn8J3XK
DUV4Fd610OAJwasdfQmF8NgCuFHqG/SX0aX7J36V4ly+lc4V6p+X2EKLFOZJKFUfSKLmHVaiWCa/
5qgTdDmHjjeen6wyTvUasCYVZR5hwRAVxtZ8pyb9ZtkmJICY0gR9JhA6OyQCHtslg1qGiKYKlEnJ
n8K1m2vHBihSScMB6dIB97X0VqxfFmtQF79hkrrweiFg5w5n8u/2JmcBuCMFNkdZp5B3wQYQ+YeU
MFIUquW4ZdyixavLEb2RsbXmWjxNpha987NCFJaWxZNlFX1IEXfg9VERXRqrsoOZT30Y87PZAezl
SJjYKgf7+G/CwtdKMZY48yk7W1+JDuf/14W6nTh9qUQbcyVJ425C10cgGh63jbXqvilKMNbP28pe
ggf3TimUkLh1v1h0K2azUvDjPmUiLpkNRM4El+K6iMzOCZbrcnasiYWOoYoxCRcHeWzB3b0Q54Tt
DljGqx/BcDEEanBnXafKIkG22h6zERZzM3xkw15NZ5//Kk/C7rJMmizvnkHlZe9S5J5h4UjoSUOJ
cLPAFwmDkiiIi3CPXNRsJOTOs2pcMynNkcssjbcYwNMEdk6MufhcpMOiLSx4q7p07KOrlWuHvzpw
QF7cBfr314zIyi4JxSXZGdBUuAjYiCU5dD85CY8knVJQLsQKLfCdOZF8sxpqRbpVAFoeEr+Pp9Ek
4PylHQnHEdUssySgMFd7gbKJUR1kI19Xc8ZvH1qibF6B1MWmG+zxeh2CuJqtL9ddoOaQAemtl+lb
sIl3mIMUu2hzEAr5jqTwtRqXR9CgeWCpAHpcHJzqfShzcDLVoRIb+MGS0+BQan0WUBYUH0/vDNyV
Kmj4eh++rZuGdf3mH/6LTxh8tiDudnP56D5t/opphLQ9pKT+kwUN4bJP0OHF4oGAbzlTeXzprNen
xp/zHNGPEejPooEkKpiaHR26WFtl36TIXQQvcE47dH+c9IE3so9s86o9xWIDDm7bnuckkdfD6RP4
sDo9TPk+ezaoZ8ymaT0ADjkFVtuycLw1Zifyg/p3LMAbtnJ9hHVGB9dETTEG+DkAwE7W4QnWF9X1
UjoB2Owb88AoVK75Tc5y+Dgrcxz5HWuxplICJb26INSVldPJkKiujiSQuszfdHOm5BBLWd/efQe6
RfrTrTlRWBRnOiDVSUkalTng3cr96aBc6RKzz1U91paB+HaxCeHdOfypidgQNcPjDFCkX+RjvFwL
ZrWrt9jfwDNAb2pjqlE2GiubWsOnt7rluTpf3xWfZZz7IdR+BEqkYkZWOufA/eB5AOr/zujdcyHO
H+nj+uE6pJ3Lom4TgIb+hln11y81SkhMcgnyqi6K1EhnPo/ppFIJ9WUHcukIyM0Dy2zSRgG3qgxV
dAmEcg8D+xOSSlj6Vy9WYz6Kr/8JVQC5UrrUpc+r579+E7/APA3iaadLHBo0vprmcZSyoWPj+IPW
35XkGuTv4w59eSeBE/0yFrz2f+8yceURKW/dryRkDuporHlnFD1QkW9zuTkP2Yx4ijLQgJJ34jRG
IJ6GjO0G8NE6Csit+9du8aeua91gXrZ0UDXRmgxmNUOhFwVNxt8qPbRTm7BEIRLGkmR4rQK86unl
LfDKMfpj6ZvXVP196J79xuQKprhjT2rw4MWXjR/QTJQKW21inLXlXkDTYs8vI5js4YKmFmkfur3S
Kkvgyln/w2LHvEdnCmAGpvyH6dFnSQd5yr2ibQtJh59S77DUqkfGHWaa2OeYdjZq00G3HsoQGKMx
esOSwQlmdS9n0YgyGbwJUqqka5QgUY4bdonLl5IDUlFhv2ZeOpPuyRzQJ9zy8KojDGqVgY7VVf/m
16RSfECEzoY54P67NmByXVYh+lXhTkQWobcEagJne+xwxzS7qeon3AvYm3JRkOXOppJ1fwe766Py
t2nJYPOAdF+vOVNtp+AnBzmEMUb1tHRJ+IaeOzYUCETHx9Px8koUWgfn4qdkh3OijhdI5Hd6OHw8
lj4zCtIDGwBPNCsnTJAPmKw9meS/cYdHQUiGGMSmppS8g3ShlP3KxMT/4Y7wyS6PkAYQsEV8dhQK
MaqxnhM70LAD6GYaITDhV1iEX07Am2gpIKQD+LxI8BVMilJHNf6sOgHGj/vX+2SjQ/madBkXbZJm
0Fy/4D93rYzI8guTXiId4A1AsXgArvliwJi0r9Q/IdlzacSyc5evAvDHW6VEsDSAXg8GEXWOotbI
wgcGRAhvF50xQd9mUXSo1XARXauN14Rf8L+xTDnpbdTznW40YznVWZhS0Glku+HycNs+mDc5nn1W
vgGW3CJKBaMviX4Y25uff3EMVStULRQcgS03gLO1251ujXJTmW/KTdpHFNAlFxcRKdOep7OzRLWE
dsbWbBEbE0f/l9C2WkvZKZt+8MEp2aQ/XB3z8dYwFAdi9J7HUJyflmELHS35U/bQzS16CiLvJj7F
/24U9+l2fvKMzlVMQzSAe+SUZm8pIBRjOm8i5WPf8XkxhCDUvW+GQuJKN3LcfZsCD5mWxoO62pza
BgmzhxS34GfDNVnT4Df/0aJOF7irbvco5Zgc0kJKH/t2HxFd+fPxaRHLre2TBo007vb9IKUBo5zg
z4FTtX7USwUcXOIB4DSmijwoI9Ss7rDMr0ztS4zKuRLfqusDtjHmuwXyl6bRxIdUuKGkxJn2pTAn
Il7ap1Y6aUZKEnAoBo571RbvdCxZDdNRqXcrX1OBHLzIuMt0WggiAP9H+VHLHI05oG3cLupKpQYO
PUZUIL4oyj2kex4ID6rj/0bwuWet74b4RpfVkJSQzlTpgpJB9vptb0iCwYkThMzDo/v33W54k6EB
xjTTlRINH2R5Xxr6uGBPwl8YeqCyazIcPe3siE3P0ONpGAkU6YofAN5ZE39EUWyB7Vq/s6AGk8lL
+wRDF8pMmHu4OCyrjKgY6C98gVXkFY39rFd6yyv3vnno54Uuyr1hDTrFaVg0MwuFKaW+CAGZV8FN
Mpnbch1IYdrGmflXyIUnfKymlw79jFO/7qoiU/VRuEROlv/6UT74eMRpdaG1s9gZNkEw1HOuHHmB
tpUwhKepy9TdwqcDPdHJ/7BHFZAGLxO79/3z4y46C7mrFjyXPj1zMgBW6iYUb/SmN2wqMu0nM/A8
SXiDqyZwZEOq+jK7tnsFUB8rfRK9tw9/mk0T/5LgtNQvG+tbXxIFFrirp/RMuOKjuyBJz2TtJHs7
QLnHvUlGDmzb90z3inYmdbW08gnNzI1ojYSWJcbOZcOafPggQaea09zNx3e1BK+f/O1IfqHJYzql
rkdRoP4CuV49ho3GiQgxIonHqTk1t8zqqUPnOxJNJyvyt1yLqpv0N2BWSpbTcWFg+NkAjdlF1OyY
fmRurC7cgzy4SZFgw1sFPYTsnXMikBwmqAVdXaktPbVCDaa0+dp/rm5rI+UybJcK+p1qSbXSUj9l
PinWTq6NjkB4Ax8bFAhpMrAdpzHq+9+y6jHxMneRn/4y7wRUz1vCYNeEOiu9Czu/imYi/TMRvwQg
/zRAExor+99YrQstEvE5+/CMoeFf5LSJ07DMz+TB7IZGueoOUe0QJ02F9FCLbf8NocVkxa5tF41L
UGL1dr0M4z6IizCBQ0niK2ctYb/hw1FUr+mSaEOAsA7GNPlgBIv2p1kJQYYuUKFaTCZRLe/fsU8t
65JrMNPbd/HWlPYhvneX5rJvLoMycLPa4OtWggrSgiAGcwiXSIGAB2tEYPnyNkuOq7bLP5GYXJ2W
wJWn5KStd7XXU+RYHxHp+a7c7QpqGD5/ZxNIpgiDsy4xgc5hRX493kgdwogaytO1V2oD1b9uWg6y
9KcgMEZBJcagguIs5UJ1kTPA5HVzGiTZQlrWPjIFI606Dm/E+NpnqW+z3GWeSWI87EY91JYKxBdK
pyTncLDTXt++V6/epBPawrQx9fg+4HS4sTOEhaQO8eMjTb2HkxK3GLum6I8AyZ6uJRJGPnNar9l5
nfQMWdjhDOFAH2DpJLQYPKr001DtrfPRH3zbsx3s8pDe+WjeH7RxqCW5QZQ7h1t/HA3IqgF1IGPJ
OfCxTRYrMIxq6uLVxeZTYet4gg8pxFw/7luy18VDoLSCgFqvHalua6BjaQ+ty19Juj9a9RLqUa5r
P+ey03lmQpE3hY3kuf+xjgVO5KsJG422I+WkC8ICUP0QWObx7odt275VSDarWEhQzQOd4yLqtyhr
i3Bx/zltKcVR2nHKlabf61PHQujNPjoDSdhkEdsk9D2pfzbbTsQtXpYIKbQUdb5UJoxZUR2QI5j4
aLB48o8p5iR4LinOo67GFfuWQ4+eM+yLwz4Ba0T6ZiBpfNq2E2nkOlIprG7eoSnqVDToeCMOGOPB
6WgWR1A/cdmOPISPuKYy9QSXwqTmuggue8i1iJ5QrV3n02b9P73BKeO904m9twyiq7i1tIfRSEUy
CH6J2XzvRPH27dcC9tmaM/+GVgX4sxT39tkVAMeg8mXTPiixgZS8sCHifpgFZlQjwUR3DIyyJRlN
u7nOkSocONC0eJ+WMys4FvqhlUj/kYq3vlYbpiiwnBanV03I2S60SEavVSSZ2Qd/bsYKcVJ8tE1L
Vl20eOWavpQcMsUvVs8ewWQaKgM0wO7wdiDong19QTN8BYuE2Z45o8nJkjKr0j+DgA+o50nCRm2a
F9muRnH8MMSUNrU3zXBPRF+KW/dxEVXzQAA/Z6AssoTb7NY+BaaAf0GQtTjTN9a4ZnZiPuYt6tq/
h//C3HJubZEJtD6qpjoZ2iRWVno+hjwkMpniNwJXHJnR9fcWGTkdwI/wNqXCgXCsZ3Jq9LMAglK+
uFH17E83KyS/MDn+GiCgLVTkireuXDrHwKtVjcmipJmRuZK7aNG13s5CKbfgBniKmXCgV11hqSyE
76tgfyCKsy5sjB+FLrgR07m9DcJ2zNdO9eLTZ7QFWtMVV3xps3JHA6SqDLgRMMDMUDhZK+FR/0P0
+yssDF/D8aMILOaeM+pkyB1EhKDfUIDhYM4haJ0rj/YcvgGsx3B+XBe4Kiy7tdeurPe4gvzc4G+g
Dg2WdJNEZ024u40nBAcaDQ8dmrFs8DtQvGMtzqp6cQ6blEbJYVW/y0WybeUuH6tWTWue0dLUfXIS
qyG9v9gGIUGvz4GExZD40FkLPIoGZkA9INKKt1oa9Gold2rImxIWFS7a17JeOezcZdIhB8OLlEWo
cbpYlWvNCxlK+ENCP8jGnMeCqbqSV7WKDrKLkn7b53w4X4R2k/cE+pP2swXjj3yDbzSjt23EGsEv
hY/pytgZo//E3C98B4P2G9kEPnGvBhfc1j1G9DCe8yPYQJPPc0v0Pa5X4gQ7sIqIF6e03HKMhKVH
BRkjsMOkt4JpRnH9yNXwipgcbOJ5z9KS5+85aZzeTdex05nOKUcU5B8pdlLcxHymFxovXH3PYjc6
3gxYnPkHeg+Y4X+8hFhQ5mRndDPeePPKkNPj9ch5o9KsgHEzWjfqfNanpM4Jec+HKnTcA/3zRASd
BPJVXEUUUSBjeZb3w4t5b2pZ/RcRbTlHB6kVO4NqedDGvuMjx3xszR6T2wkI8hM0h7S8ccn7BRP8
AO7VeVgQWO/+hqBCrQ71eazG3E4d9tpOo5/AZnVhZUHp+E4ECwGH1DQRQbRfVWI5jc/k8e6isY6i
Mi8lGvIuNkwr/zLnYRmBQue93OpluxpTd9gZvBNIzc7gWrqRADVp7gwULA5qb1Z4Kjgzh2E3EkPs
vZXyjUa3HPtEP5tqqVQJEMb/dby03kaO4SOOydqF9ej6QOITGqyoMqpyDEh6/YTsGZLYz9xQpfRJ
iWWnfqHpfY6+egpI1jaH6HI6PSppDoJbL/wYcQ6uXSoWP+V0Hqni6O5e1du/suL6z/nwtJYooBM5
8LYP8GCEUYCVG4yrY5VoGLg2OVTVGgmKcZGyAFosAZbpCY9XnlhyjAmtZdnpTSRAl0rbYkFHAbFv
EUh8lVez+l2vy/2d5QScwnpeaup7KkKSvVCOUBiIOTT4dp0QW9dc6XvKwiiM+fqbVgWgZcI1Y25o
nXCw7roCwzG74gqQgObQjkQiUalLiFR3Hh2iiSXAHTijYtcGKI1w4VbIaE8LgijkjlgRaAJVllvW
Ls9MmC1Remed14jWC39byNM2X47FYmOcUEJSZOkdm25J/MK0yihP92vE6YhHwy3qtuqc6hmZhoDH
lJwOOoq4xJaOUeurnkWY5792rfCGg3uffhnPrffpkFZ55TIz7tVu01qfCXbVxjdfiNJCDI2ZyHg9
Bfdh8JV/gX41O3FheGOnvbDu7DhdzM0PploMudUmXxUHn4Br88QoBoGPhF3xQ5sCuVZtru5brF4B
pJkbWL3Rm0rJZQ0tO0d3Z9qObgevh7jUMJxnnLHkP28usC9fYaOTbqAPT7jybqwx8dmwZRPiTVUs
syuqFgH2ZzbX/l+b+ZcklPdR/vyrIHsMw2gbimRZ5r2r+xf/BWdEwoIXfh/rSmnXVMNelCbgJNCs
eGVoRIy9iWabpXfJaTyNvz2XMZ4wYH17qqW1g1JKiG0LCI51oRj99fmXuHVNBTHOe58zYENYHxfu
T0wg/ZstiTJQvzoEh4qzwdcU6T8r0Bc/tVqz/HMsnoe/dByaf6ZzLdw40DqtVq+2HXdHjz+nmq8Q
KNvXgkUpF0ny/vtWea5IRLZ0lnVXrNB5fgogLbqeUr8Glqly1UHQRywKZPFnTdLevVGdu0QNV+jX
f/Sgql4u7J4/+fA3ICdnInkywxs301jDXRWfjLX0kusPg8BDSwHX9u7kXYiw5TN+Huw6AuhLRPja
3XG/O+24R81uMrl6nJeMBcr7Uyr6xUj7a9PHS4zCexNqcSVa2FzSRO4X9WkMSuKYOZtOJ2qFQYko
wKr2HW5q6z0akttUhBPPGl15Nvgc0Zyj7orlFssN74lpJPHjmbNRbmbAKDFjR+/I7sKh5KRUsvKa
+u+dxLG1U9CnqwsAcwUdcqVvs5aD+xrehfEbVa/0ro9b8qDd0+x9O0wHy7nJQMhlFSjEpzN6fVcr
jgMszWoUyGC9ReSB1ytJEDReQzEUqL4ZyqYuDZvlD2mcu1aqHdtBFa6NcnArdDERxJ5nudXoEH6M
+jrDw7Z8JdW1hUJUOOQDIQGab+UE4/PtSAIaD6Bvi+GvrN/zeUFAdE7IY0PZtQBlgXhQ5toMGtaJ
HtYxj0B2R9anobMSWSOwwXSPxktVLjOEMMCCK0gDvm6jWm9+sjSqBd80JePEnssZrT+XKiKstXsx
efNgcPRpcEpnlTRc1OfESdTig53MWtdH6x1DU2JeNAlHjpXzz2z1H/eDm6KdQPUr3O1i73Eqp2Gt
EH4hjEAyUYFHZjlehADf4/BeQzY/xFEXLvUN+sT75GApmD/5xOVM0rGp7C3PbmAbkcLAzoWd8HL+
QwNMATTSdFJw+h5OcYWiSa6b+hx13p5o/A3eipO4PNmhlPUhEECAKsEfAhkzk9uiNxegyu5+hQZh
jCcwXeJF1U4M4Jqf2fE7ry531Z4HJBY6/+9hW1z+fS3sKe7to14pTloi11sQQwRm3rBMW9l9/H2G
2S57c+RVThl8iAeasSI6lgDccPT9XKsqW9e+E2fAfaVpmdijNWh4ZVNGizbJbTVsIQFtR3B274YX
e3Q19GeINBryQMnveAl+8b6sRtzpE1B44CmJ7zZVQlG5nyIsPk7MwZUeeZZTcuTrmDeGgVlQAdaR
G6fFoyeP2hAWT8yeIVBALGrcYgIhjBEVhlYk6gCATvsdAoO5RT10WkSIT7pgTd+od16R4HZDozG9
Rk3n4r0qjwekPSebciU1YIw1YiSiAE9pmawjlr++/ZiPkfniZQej3rCtd9xLwMfOZa0BIwfP0Qm8
MdgZGyCjEToFHx7g95owUeJaMiafH4O4p46Oyq5Xx7F3Ydwbo0bKymKELNxZGAB31s59kNoZ7Vvc
iqxgOzw2ix85b9/g6AWiYdonVwn0psccxiWLchWC8mp5fhX5sFvsUlw/zmxEU4+ELebYmVzH2SLw
xWeDgUBUV+77P+hN7M8YcPYmUqAumN8nrefvvXVOP4xkRDgqhEqGca6na5qjiHCU9q0dfUKD3mop
fa5HjX3FjbicimhJYNTdXeBQAPqwFt1L6UhJnYY8FRDZg/SlhUEDgfhCAR6RNjtaTyr7Lz+MJhuH
uSpV5NOK0tktX5mX+BlLCZFz7D/DrfixTzQTJf/wXxoqMpBL/g4/3ygjCaJzKuYc+F50s4L+68jF
FRZr+CUrMZCDKc2T/AuyMwl3pKANLo6uLuvegR8Rsg/MJRNbFu4bxfk9gV3neYabfv9uJjfuRPDv
1Nk97WSb/HAZqMD7laaNXknj6wU4w7TUg9jlZiE11qMI0hYguWVESsGIIaYpJY36hTHLVrowmaOm
po2RUw+djwSxTs8CFaIvLF6EHb42sYmIcSZ5u9f9EqI3XSJN6/bz5OV/99ref0HeinUghcKa0d71
qDlFs8BpMQt6VShDFbSxbQJHp7jGeJHB4rRkrTf9i6nZGq7t5C/e0ZI8rLkt/hjunYxzEdEmmLOV
4fInFF04O00Dl+XgFj7WBrPVwapCVkYi7HHu12pS5Cgmv1JqQ6Kq7YD6K5vn89hGdgWj2qm4HiWs
h5hbnJ9Vbq8gzFSrS6gzHeB07sxGul7s77f23sKLFDVjza4s+B1KQWUnA27PXBcWXuzlId17Y3nd
Ir8sVCvqBmv+5q43u/6oIyzo42+1U9Zf9LIQy+heP9hSuKoNCzZA/CdIsZLemkKd05ZNSpS+JE3Z
SpxN327JAopaOZmKrFku5D1pdfp73biHOzfAkZN+qtFW6ZZai7fX+OI7Axo/b7cWX/hmxznby6LR
3bLfFUynuPMxXxgZK1J2KkS5e+f2zzL0MFvzLWXTz9T5kXhHkJNUMUgcb2u8NROzBRzgFhtyNz97
LDTt2PURSQnltQ0Ce1GwjrKXifVWejebGnqjYPVJag3WTKE2q2YJ9oz0iefQoT96Qvt1Sq4KolKw
5HgNrzOGqS3sI28XPgw0xFjQ15olkh1ltYcNBcsHsEFQCLRYl8GpPqe/PVthMqXT7Geidzp8CK4S
i7v2dSfVjq6jsQkGjmIXkRR7bmVw4avh0b/cRc9hs1qbmBDJP3+mrb5Tq65ID1YMF8piOXhvyQHX
pgEWCKZOx+vA/J14mwR5UAOpWKAduOKuke7BNFESmXMBJ35YycWeho5kobawweLIdig83UoJqGTe
Q6KhKHdIX45axRkFcpEQK9/v92hf1riXCL2PS1mrr4TXlUxyy3N8kIcFyXnXk2J7/qh9lFzuS2w4
CeMlR9rguhH6IVGavc75nInrm6XfmN76RPbheeGCILE9nC1HejgxANcUpRhlw3xvNduWQmBdEOLi
jE7toJfzKM3YLSzIGpBj37KcuHhDHbXJ00XklBJIinuLIneTv6tqKgAL1ccjWbknYVH1YeVmkZSQ
ZazBhpr22xF373lmK8VChZvNs2SJqkoNSR8GSAVJVxsdaIAhiEDMWtwq5GwJk2KPG/8vbQd6MWpz
6tTMChMiMlXSNBHTlMah+vT2xo6Z1kpd5ORjdbfXn9VRTNluxFN5YskmIy3IsRcoQQxFCKEjkOdr
n6nZrT/JsPGZzfwm4CxqB55rufHo4YQH8D0XhuXAtNve//lsHGRceNJctn+b0WXoT+utqxn0S6aO
Am2MXdDdIs3mLbt1JfxuWGtigkOSxz9tFps5cuCC0tfZWeVnAjQyigo+opePkPnNirbViB4iftCv
CiajBso/8vYFFYEJizY9sD0PbWIar1KDzxMUTz4ivGisQvJ0YaBaknaq8Nwem/yv1wglKqsL3eFM
64vy+UyaOOqeWxbDAsAt7CXEvSJCopUXmHVGcZMRAdwPtlIUKn9sHBrI8UyFkO1O73cbwNZt0pJ7
FUmJoc3XgddudnXIfwymHGeyxHwJzCBYPrAK5LCDEewyVniac/BFcVO8bTgpmjlXA27miNZlyg7V
3DwHDeV6C1IeY+E70LmrzT70Xat2N1DXVKq5IXSTT12EgRCO+uCQHO8KpHyH7CRlcIFGt4dP+/+N
H+sD/1ZDDdNDAjfn5UrSPycvGUtZA0A78kD8W9H8gqm2bXI5/xeLPnidEJPpig/gjTM6eCJuUKsP
qCJYRUDrKByDp+xlLIKyCdoB7shVCAP+LO1wkt2y3cJouH+uThrcNlT1UGajHo9oBa9/fg/1HxFX
+WAS5q9hdi1qjE3pS1manw5c63stk/JwrzZEXIxna/phipGrUyoWBiXpjD0AkAR+K0lJOWLacc7A
dj5PbO5fJExBGEKvAUa5UlYgryrk1++p7lvUCtn1WhzyVSpYMCfRuuH0rajMlY/Mv+8HoruC+QBh
faoR2uohQ6QPkmWaN8Aj9z0FqNzDmD2JFxIhCIEttcccTgl6ROz0274MHI6nxYE93PRlhJrsJUP+
mMC8HRYcpmpZS09dR39zkgNKFqDIPp+sCxIEyTQCo+/JrIVSFEj90Vvjsyu1VHqoL0ft9e/eiqpQ
SOwIx3i3yB/Gfv6WkUIXyaJIu505n39FVawq7J/3iXv4xJ4eBSCEy1g6pslOCBLgaRvVWqzO9+Jv
1MS9ER4Nbpy1m6Jaa5rpaqKeB6Zc7xk1/zIZYTIe++6FP2AiviSmfSkUUF56f9Bf1IzyEEPLHVNK
x26lQAc29F1fo89nMysYKkr2HSK198eIsk+0wf8CurmnAb1mxCE7hsEh9I8qRihG9PjmfeuMW+4B
uLsgxw1kw1kpcSxSCq4gOjYLl66mTWiQ7OmD6RCEmisvt1C6jwQ3TLuazjV3SzGZJW4JTH7aWUiN
8Qchy37OSv7QHa8KF6X3kd8ZvzD6/3kgTEvrVgyRtSJ0eIEx3PUObmKBr5sFfKADRc+ne0Njz/tW
JGHP8mIFp6Ih9bu8RsNm4G5tsWwKw5MXbHxvm2txY4bE4w2zxyZuqbkViG4Y7RUVN1qlpFsuF7Tt
JlXdZsRuwV9ks+G5Ka1iIhJos5DFaeJE/enoJm0U3c+yJwelM/m+ZkaPCv4sabN6Y+uGXJbayNsj
UQUOkgZ6eAcRe19GZjGO/6MmfVmlrbAmSBD3RFCdVZ2IqMsgLiNEeNV7RGWszPXmV2nRg2c2OFlz
8hdLxMGEzYEuHlYv/uzq4ISSVBr8pSfzlJft1h9Z8XNennD7GyOvnXuilAzrFlJRMzcMxHNDeC+I
p2jUS+UFi6SjuK+HVDfqGfDvIn4I5RYtXjpC8oiFMrkbuCcezHuKTqQwe2xkUgvW4wSo+zvUdOll
dyapWdVCWox5OTdk9E8BEQ/ESsk2Ldb67BinFbkkAJvg0actIzP62cjXaG43/5L6CJkPZR+2Xjqt
qLCIUzoWiQMKVg0uM2KNt6b2W6sBo5MG9snl33dc6h7mo8cmvdgY6T2C5WjcUmOEvmRe5F068YPP
ZyASehjhkmVg2dh6/k1S6/w1sdiRLUXccSQtdQqCMOIxckO1cSfRqOOX0mbKmW/rSgQFIumQPYLh
xV9KbSNDdSjb2HTj+kfeS9UpqhpnQ3vkN2eSipuf3yt5kt2iFsYWWK1eVqiIuYVT5JfMmqkX6/ys
qI/yHaWVchU/pAo8t9w3n6ys0XqHxhaaAf76oFTTXGti/B2AWMvOcarUPfqKYN155qb3KwygoZkH
tBneoqSaljqSD3C/aJ91L7QtHuU0sjnOhxNEG5H6h50ZgyVHLHmYhpliTKBnzN18KvvI196ynl+v
kJ80I+AXAK304u0eaRP425etaCgBqmOghnuhyLJki+tlffRsJIkIhFw4P0l+MwCzn5W/P19luIw/
Dzv+tPNAYSnrgYRCoT16Uxj/NFbXVjDRp72D/s34PjAq6UVowrEWQlOhpBNRz1K94JPQMz935A1h
nUgBOsymi/v2PA+0X0SPjzacTNbFHka/OCBF/aEtFzXqbJqF6n8pS9pp0vIvB/xMs/dtDMY0ndZB
GCjdeVWlA7Q2Ey/dWkrTEuw7n0oL3gbZhuRsviWe6ZQU/NTp7t+vjC1vTNahMFIBp5Gdxn1KDJVf
LjriqbKj3EKQFoX5aA5+ToQM37xmH/4twXOPEHljlRArFMlvoVEOMxH9LQzghxxxdudh0g3enEIE
ixZ/gWMOdziCxw3IBrCymAZBCPQ53hDnKYCpHZh9Mb9DdC3wLrxRPKFX7/ez/DuArSE4WDQfxZog
cwDdomLUmqc22iChmHR9hn+9Euyvr1KuSMIADQXTt14OALo3hJuyvOaoIfJEv7NhI5Qg2SUBuqI9
dPYXYCQL6q8BwF/PY56UYutHaew8b3VTATS9Rq57kgJzXtTg6mBXWa7hWQAYcpoQ72GzsVGsGDvc
diFa/Tqr1QksT+3STrBt+ptKpwVGu6CvBtpnMRvIY6qsUnkUli7aJHHMss+sQtFMnF61sZdyXRia
L7t5I9SWtvWxGHkq5H34K2MPZ98FxFszg7j4Mtfe3UlSew9lfn32pW9HwV5LGMmmEZqLZYEH7fGS
0Izay74CYtDHZ47in0B7yU1GLgTC2OTtcmjW6wKojsayuRmoicJ3psYea5v6894oYEBmaCJhy/+4
2fgizPzZ3oLXjtejKKuQa2Srh6ZZYQUmQ+6rncbSwMMAAwtIENrPZ1kd2BqTv87PUm39h1oAi1Zt
5r3tylBxEJmK+VdLBSPb+WHUy5R4JbopCWILtPslw3G8QCbAzG8F5MIYP5Kc+U3cBui0qWCISnYN
ZUl+gbAg4rtARFNBWPWkl4kmwufwJGQd6aWtjxMBQXv38NpqLh9iRozA5vuHapn+trE28TX3knhz
NYi7e4pmF2B4HWxjCxfqpo2Rxc1jkLeOvdodh+dKoUz462n94JkkfmOikRW6dHIzuomw95J1NhT4
RTkRFbDqg1WoF/7/x+Cf+82XttSp8v2q3wdlL+HDJra+qzE5XHlqbja2HlKzYQxjoOPIFSyi66Bn
jWXuzcgKZ3p66A6FkOEbK8SMbo1RU/9ycvJdpdpP56OqGawQve28tzaksK0V/K2MyYx3wD0QbgxW
55HARUbx0ej7tmlhzsKpmvvKCWoCfpvM/OLi+bgBNx9Nzi04EEMwXWCQ4+yJ2sGwXFaRD4DuGvSR
+Y5s6TFOp959h3IiiQlDDfaWaBl5h2cq07Px/5lQ1G/Hb99S3W23CH3for0QUo0IF+HN8hCNhzVY
Nsy50jeCcEZyeBVXXv1Y+NqdmA3K3wlzhvk/2VcDNu0yLn83RgVaj2S9iG5fjzrAJ4u9U61ZtM1W
KCZlZYgjGJm51iz3/7VA2ZapNP3SM0ExH4nFL99bfS+hFE9rsHjzBhuXH43sbENiPC4whpsBKa/I
vuBL7PGoz5CH/dja/jmlB5GQ/E80Ccx2XXbsra9AU09zlTtDBa1VIPQNTk4BSd63yO3u5/xvTyY6
QO8seym3BqXkdFievoO8j61FatFb2X/UTa1E2jkLIAXyg8D/+6SwwAl5+r2hPKbjBccm/CMggmgs
CMqoS/qlcuQNEVJ7n8+9UlxuURjxnYhLPuMPrfJptb0N19UI6sbgaeqGXJkReuSezNeqgTKCfKec
TtDFilK61/3/+NNMv9WGM7OpsNgUf9mRaJl6urVULd61JEa0hNUzD7dPntw1RQKEFImzU4tD/yMQ
IKbAHDGjy/oIVVA2G+2DDf/Lfed1SU6xbxhRYh3Fe8Z4UChm7o/EOxfyrrMHpc0gKvSwvbVh0EdI
Bdoif/CqqZ1yfs0RkIM4+/ExUmTOxm5mWZFBoqEABATVfPq/79HXxl2McPns9MEV0WWOL8BiuB2v
v4G+0yG9aOEfDCR2X9B4yOk754vqEuKm0ynNLYfDWcCNAziLe0D5BY87mY0x5cSvkSxA2F8kPk6U
K3qE0VVTuf7/ERNYqBt4GhwytFTHeIPSbSS7EcPANH91BDwDeUFRo6Wa5vtnwJ7AZD1mSt4g3ayM
0QFwM+6oloMEfAHmeDowS9LrbGdAQCmdsW7NbEJF/v5hPQy+fKX7OyQm1g1LXqd3qdsYgPn89v+/
7R7jEnl+q2Q3duixvBgxe8+s2RJ7lApeH8JPsCf+PIw3YAqWHg14wMUqPeL9gvKoluNHPxooX5x1
aKL2/CgfawqMZe0GV8fTzjKtytO4XA5FRaMBEsr48L1gQQvsfAo8n6xBbx1xY8VMx/YiwxkTeoHp
DUhAMiu9L9w8m/ACfjzhFy0eXqM+V66phEY9Px0bnmO9qoN7T7j+URfWnH356Cvzw/Lc/i7yGI4y
RLFdEdNyqpJXR8d8HrSM7jSiiYc0OvX+KqC7uHOGajyKHc96Hzs7tizldVrOy25OxJ1I1BQwOAbF
4vrTP7uv1JY9gfU/iCQBij808PHooCvBrM+muLjw0kDTgtOThrNTx2X6oOBzHWR+dSf0OBQ2tss2
uaEkFyMVgC6aQxgSuPz4Hp7tLGX90ZGr7mT3WSjjTWmv6Y2s7MqeHS3kVW1FqzMOGUGQ0VLiKgQ1
nq04EQk0lCD7H/7dhSS1+hi6IXpM8mfjFWgtHacKXdNOPCEnpu5c6e85bRf3khyCkVYCJYd/x1sr
XiHHlKYM4c3jbnan5PUciSKwnO7UEc6pcL4GQoZpub2KImCFtJiqsmXIVTVCiweBZGjYJUyEhJFG
9Iv9L2Mk++bNN8NWQ4y/MwkhmFF/OYuBrpyvZWPQroRqW3X2D6bO2bbtwGYbN3AMA8M9u9yz7h5R
NXQBpr+HepF5m/zpfGc8EXbwuABWpGdQ0tnAaPWCVMEFt134R9ci/PDWAgu3lMEEUMUE0YGYZ/uy
QdfY0GAH2Z82fVlTwPy4X5AtMtT8kdXL0emHCKqL55e1bUFCP7Cohc111jzMIMrUhKCH17qHOWct
jabKONs2VDlekJZcPlQNvub6gxVTbP/YnQHLBu3QUoTJv8BltQw4uIqe4EBbiYkBRr9jC9ivbbJy
QYJHxJX79iIH3udin6mz/uLQzV96DYEcFJByYN2EsyItShOv6fK7MDpoWoM12q1QVRhhxEsucQAa
dFQp8O14ALA6b+j1FbS9YPlGvNaaqvoIG1LO15UkIWht5kRzuZcueopv0XThv8AdxEEY3ZrmhF+p
k3BxEXxU/+rhJSpDBava/TrO7ivWDZv9NHE6WjuadNqMM1EqnPI38TD2eLP2mHQMCQpYfyn2ZSKr
1qhc+lDGg9rFhI4NbD/pCet2ZyM58RR8AXPr419MM2NgXp01g9kdW5ncFHKnPWiAF/T9m/E5Gf57
3CVnx+EfW38o/k0b6gHqkPnUJMjlmx13WUx/0Tpsb4Enp2NK8jOEucArJesC5HGLizvvzyS6G8sV
8A/VyIz9vr06lHZZSOVE/YyNlAXUE7l4VvTvMcwfRBsKSF/EkrQNvykGZB+wNX5Wy/89BWGhPw44
eN+GRkH/SJc8OmQi1F/w7V9ZTIJAcS4pWU/PZreK/wcJGelSb5nzCdhnNpyqR9amL0R4UiW+F9OV
M1kh4CYKOkRR2nW+mIRTq+bCuEq80lwdyK1FhCUXeHSMG9HV4pMsgD6eqRvG0eSX7cf5XAwi4F7A
K4jgybQg4fShun/MibJu0lD17X+MIovv4hDW36J1t4M0GBVx6Kg6HoShVqsPcnrBRXPWw750GQbg
/Z7GLcdZOTorQqRdL1yN/HLWMhe0XNlQtJYilZgzOxztsu/jVeleaLgbdlJ/YLm3w1BDmI+ciNxB
cFTlZxybg8I1F3C5jRf6ddXOHUV7xhtD7HBOMhz1SJzbb2Pcx89QnUmip08TJ/qr5JeqsyBtL3Ji
FsCQ/1Pq4yT2rDm26AdPkp+EYI6tj4FGQEOs3bgj0tVVB9E51ZkjrUBDhw8iSLBm36UX36J4XFZw
YkTLsLPcQY6ui4x8ZbJU/qMMkVLiISn8WSWDygTH1b+lEOcRk1LzGyW6GRNCtwmdbUThCgUAgpRP
SqN6ApeJdwnyeDPgQy728uPQpCOpnTUeFo9/yQB7yO3C5bl2oPFjLt3ASjoXDHiiPBgxqsd8Pau+
XSzqcQvn5p8czhjXGA3lxAvNhPyLfp4g8dPhhQeHRG9F/Hgp/KjborNeicA+rsr1XCjbOlbgPqfH
OUmyfWYBnG7OONBxcPd4lPKi0tYoS8LmiorJjFPIRirrfI9ULOqfOYt1WKuHgjAExvfAZzdaN/dF
RQU+t2PVFVfkh2WUzbPjbI7rYBswf/P9J50WGRtXzQGlMYI6Gk98KimZ3iSG6sKR7c3c4muiXNGo
sMu1Qk/vfIJ1HfKhiJcOddujrZ3PVHxW96kqiDB86vCiLbSqwyuiH3tW+YYVd6IMFc9P0xQ8LhxO
d2wfrDKSgMzIZYTYruEzHVS+H3lX7caUAcaVUn2AeJmFjXKf08wPff9ZenlgOMVChNmJaKu7kwTw
UTgYetfRM1tuHmGYkeGxOpweyNDpUAKPmkOGSAUwBHP5JOOfu38DRw6f1OUDVj8jBxM8yWPf68pP
UxC70lIbUb9YQ7nxU02KR7R8eN5Qse8i+u3dVotB6iDegthThXiq1RDsowWSpaygeIBKE1hzTrLY
L+oSLp4BiYdLLNkgNS8eScbk+t27/agWtneViwxHV/HZ1s/rsVHPgF6s3yXR9WwiftYZJSPjLn5X
7cLn8kNUSAqf5A60ljC/OmOJ9GsNKbruglT/HjVqO1k2WO0+hQZOtjs671tFei5Jc29r2XDRVvKD
Yx6FjnU8b3RTcVZS6Wlk4XctSrKh6FJ5nT/niidQf2vV90h7VpGI8Ti+mrZL5Zn/b3kPvozsaFfg
31w632Y55qZMm5fob8051P6d1i+T3H79NRWs0QUNZfrEpQSq9GLMVCvsEMoPkm6MlEf3hhZ3u3Wk
maFqLMDfVoKbeflr8JazMbmqqIXsblL1t9UxgTaY4/ARgzgGMQzeRK3kG8ia/AajITfWXvfr68u4
MrewS8+jI/8jFJzBkto6Li2b+Wsa8f+E0Lm402YusPfqKVWwTqLmzr4EVXZpsv2667X8kgstdeqs
kOkXb5ZcrxdCJfgPCTnlIYXKxovrK7ilKZojdWdQ1hSoE7mQ1nrDubkdmYkOPBqjO28drjNnptFm
rXu+Qrt9cWNN1oObFBSKechjzKjyZKnaOISsYfZ0aPmvMxmqnsIvzNs/vNL75VfCxgOwWl39h608
8DvkDPDJF/O5m1itFoSLmK70Q8gAvvJ4u20kxAHg9c5GKFLxatfTF+DR39MSx7GBeZnPENctxMHk
ug4I68sJhE5JuJB9ouchQodYMZm3EtkJfcUtgBlyN9JnxjJFd9cA6HmwMgPgnmmxqfWAGl9OkjO1
UFd0xRHaVZiqA1TPsQWKEOwGegBeEx+cAYBHyk5TTADR2yeb2bclkJ/7pMrvbxURM19WFengJiwR
7+Rumw0Pg+kBSRQP8/2Uh4ukcMFnjPFtaYKlqXk5E8nBgRacLTqd5/u5ri3FjfxXWOQpGy8SY8m9
hez6ZogDwGJ2asUB17etlCQ4XrZSOlqnJtt4Ka41ms6KTQJ8x3KGHS1jsHU/KwemHcb8HrV5CEPb
OGKvBrQhcWSgq7djPOemB4iOVK55DM8KiCfROjV8ZA3ZqLzEHSKKMH06HH4+zlqsuvHzZdUhscWm
mPWiFeJkH92c0hRv0VAVBM9amPsXFTGajLVfSyA3w0kNtlujJjECfLw4GVMyaTuyqwA8qz7T3meT
5noAhcaKV/ff0QNTB5NJcHsRwVA7GEtytNMURjULk0VGKEHCt/MkncpkdCYVXi8u45Gsg29aAKL1
cA+AkV0tCHY7YjX2PBNUtOvTbyoNTAWi9OB1F51/o0Me7SCOSgSfRMOKM5JQCVqtg29Y6wlFbafH
AaKeqwgdSRAtMTm8MCESzWYdCendsStYcEa0RX9gCGGWH8wBn/izI/C6/IQjnb+ve0ZdeT5+K4sQ
lA3j0vTn1UK/cowYK5BMfI3432YoE6I90T/QaNLaO0YcxRPmtnQ6mS19FULSljDba77PAWkADF6K
Px6Mch5oBHY3/NLevfBs/274gTuMpFoF2trPEWL3+aJG308+t7cqUgdcX2BWjqLPQ/lxMWorJlBP
M1V9D5yglQT0o6hVktt+zFi0Ih0Q6JD1G47A7Gc4/M5qJxT3eN+HvmT/bdU2N4cEG+XKjNO18MjW
HVW65Fl65lDllGtUQDN+fuYDpr9JD0PljbLleNp/J2O7BMLqGiVkDsSX6tOzVJQCdbJvyOQ09m2u
OmmAnFbJdhg9JY/tAwPcbCaeK25D0geiIj8ls+AUPXy4YAyMIBmU5DsxRfv/p+/h2GbRXNvBxoAk
AnE9ZgjwQ+Tbvs785DSyxsSm/xF/ToF0Xpa25EWgVfwiLCEdZGy843dqsw3zuwO80n6fE6Vo8xIM
tbdZoNacdTXZOe2M+C4nJVod+Rz5VYCjWIMFXuhLI6wYOIiHBE2A72qJxpCpz2HVnSppi8LZ9ltj
1JHtrhuUzCnOc5jKjnjnc1Wy9I6jzWl91M+fOBormEaDf9kGA2usHeQxwGd/7nMGe4yaAvGmfCfi
hC5y9bsmAJ7fqI7IYQnZkN/ugUHdbigxRZLTZhYfnFRS1s5DGWBG9fmwhHfkzSJjLGuEupZUwXQu
cn74MdSXgWcwVia4w+1pDSKeeY+xlYSbeLnSlOFaL2bDQxP/oFBdhcZFE46kod2CTV4mFr3iW6Yk
dnK3K3WprwHOmEkMiyCVmKgA3Ez9F1Usw+FzgeseWnWl4+R9NFIH/PusBnITM3vRKY85dtJZrf/G
NFOX7CHycyZVjPZl49UNa+xGhpZxinmpGBvBPoQ+EUI8UJzISk+yrd2A3sx8H/m5ZTuKbZPkstS1
iOPukHk31VzoTyqwlT86Gs++JzRVFJiPNp7LiTdG0eaaYZ59oytQL9wADM3ibufVSpgIT4x6rDQW
7U10W+Uba/BVCAGReNL9+WyKm+GIbKsiVN+e/5/R2K4gKSq1FSvi/kHoptLnxJWo2I6eeZi1YOWr
+rQ+9iPLylfRRSkjE3afK36yeLCKxhHbSS9EgsiM3zz2kK8GMRT0pJ1YsUk3nQ1DRZ+OoIApaODe
BDV2JupLF7mrbysPFfbyUibfQASRgE7p9o16Cxx63nuND0lSGkIVd7YJmDAzQthN0ZnF7FTP/odT
hEIJEv9FLL0JrIaf2telOQZh6IfoKOB7benkWX7rDeIbj+GPXNozAEOf+toQkhUcKspoNU5g/QIz
X8pzhwy4SY94cR7GNHeBvtL2oAkxw2CwArNIqGcVprGjD2NfMU0nAKhsL5qgTs8IFKY6hOKldr61
PlKzIlD86DAZxyLJPoSwEPigNh8f0TzMML8rFY/jTFisYkbaOdWDnzSVUjXZqe4HdyBlHJ/WlWGD
9dOsqlbBJGXd3Kq9dUqv4AXktFsVDTJVdfbs6B4NanEwyHdT0QKojp3p8jcxBc/2iJpcGzdKxHjR
lGMc15Rut0CK+tP7RjpsKiMz0A+Rg1imTcbB2W24Vgb/4GHYV+WBt2H7pEmdxpWhWBnOjimm5dl4
6FlZL28vYFN49686E32nVRG59L5v8loplhC0t+gpUX/dp6vX2zU4Bn+0bY2880mvKG+zYIkF+grC
MjwmL+sGhHH3znylLZmaWjzo6U6boUo6QmwvrVJtCi8xmlldMPRBthZvrRIm5ybcG7dza1t0qJDl
zismpftwGYacifLN0E09yjSu6w9AV1v7cPc6zij0bBTv/sOYdUuywycbDd655Q/d1s5wspuBqa/y
8dfvSX7Yw5doOKM68Ipvq+EHmxESUr6aNWpUIeZvVb6Pt3ob+7A4MV5TR2sgriDH/JoZ5EQrwSpQ
aO17W/r6UVwP0Bf6yUSosDg/tkaeQVrLDTP9gcZS/IP9zHZt/ahhzObOrm5l5M7KxCGFrfJgSJ1J
bIdh6BTAu8cm8HtecTgeKcV95F4M2lHd9MJDGpWaP5ZhTyjYmABRgeiMzEvlzX2rQe/+vl+171yt
00sapKJM3mvwjAq+nXQA1Jkxv+YWq7N/So39wcYh1uz2bgly7eGbaVKGnZctRDuDwss87FbaSFaN
eoTDTyw2pV2isJoVwjLObbrTTwfTcg7gusN6dcBzWjYzvj2o7wt+wJ/JLQ9odDmscCuP7uG7ZxAR
Pcohz7aW3ZJLEi1F1zbw91KrzkojLA+dQ8/cpx9XWGVDjzzN3RNyZr+wUlPlyLDw3CHT8m9NNdTz
jb9dNiUOpk6cnVHExTqWvFqGsl32uoZ/aA3KkYwAYh4zzrPyWqi7hmhAHsJaKjgZYzoQD+92aVnT
imWYGhKMwGVtdqW0DML30bBu/eslVhCvmLpo2htb+tmLxf/6r9+dW8wE35VhC5TsZzRGzYV8Uuat
xAlAYuLQ+2qb09dMFo+BG9gBFr+1lENiqE3GocHXNH6734U647I7CW7e/E6JQxNgfi5nWw79EvZL
flOLAUyrtbkDwRNp4f2LsL/sBCjWAyAN1rePD8KOyMyStKOhlaFMApDFRTYlepqHegjTywM0P4BJ
UfkE4G01JCij4y9oifwmL1p2qki4lMRE2hlZsJGHHjnEyI2aaGizRKfSyDnp+gQPCDrTAVBnMPlT
oQD0jJH+PAHhjC2haDl3Co8Ufk8ePI2o68EzDLZiMkaLembCMmccpMaTHHggreQte3LJJTDYIgPF
h8P0hoqlxd5L5/tHgH/+1P/cBiJzqKSnBeBAxT6nQNG0mJp7YPeG+Au84K/zHcfp5+1laBNXknTZ
YqTntAVrcAg74PFu/iXlD88eCpCXJAvj7OL9XhB8DjHHsB4Y0zvLcvihUERfPGc/8xiVtXHrMMLn
3U8rjEoZJCyL9m6qjS8r9xhMoVZxKSYedVDBryKD5ea7a4vUcb+DJwiVHGU4vH0R3+BramaB0WOn
8RES5nmiu9+7WF1aupxpJD6NAAwGwLSRQWefsgnGK0WiY9OXDrpghQxQdLRUHMiA7L6lV7BNqJ8r
Q6f5bXDP40f7Ti8/CB7aPkW74V68l/lVd2KkIPP/oZ+lT8tuanlICsRr0ix4Us4wnm27Si4NQr3f
UbvkcV96DC96gcquTfeBHTo6MK2G2k4w43WpaYKstTpC3fxlll5Sa4DLhRb2Fgi4Bja2tWeAXlwM
R44umshxQzd2h5jk5VCY0yyyhjHNL2aUAIVBHg4+dKqQSs12YhCTHEmsfwYlSwgsxF05nkQzMkVP
gDwAy8fJEW8ccqPNS6FNA3tNdh6CMZCtweNexvrhyxJnZxqGmeSPZ6xkHFS1pUW/3H8bW9zgrhiJ
1/VOQUsG327nXBFcVpf3xxgL05DdtcfTmIvUqu/Ao8qAf72b/orNC4kH5GZcK8bgAp5Tz4z2BEMR
OPxBtxAVYPEvizicXQsYuWmzYoNrYtcCdF0kW2aIvLM0yaDzqTo6hr0IAwJ0g59dH6E+tOwkc6mY
7vfZyxeK1HPMQUFrnVkAJqdsgUSJT28zXUZM4roC6qEDfTlBoOYRQSPXsPzgfg1PSV8wIKNGlzzS
XSjfexmXZXNhA1lX/SnWkMjonmUbeMYjuTNnHscDteezcUTKZUnfruh+/3hi111hq4R9oEXG6vC9
nOkmu/ulypKLHHCv+clAjQKxxQfltaMgvb7/Ux5PgqB+5oKA12OMXZA++AjZwidkP0KZnPMbLj4P
IyQp2OEdhREjkJ3/C5Peifdmb6r1m3R5CQXv0QdbVlBaqrueVDWkjDDmonLDFNSGR+IOMmGoWEMY
fvQ/F3vbJPYq0gs2OzByByfHtfnbO4tuUB74pWNDtZmPTfCEZXUogdaG/GW8P6+i+24/XPg2ycXu
5EzGmFyJ9ALC2qdtVWHtkbC3Km+MfnGaGqu+M8K14AenN0sBvl03ag7ihPA1/6yHvsghSFRi3w08
32mnqrMY1pPu9bvN0/0G9TzatD3G4uGSJvJMnFTvgZzLX5mmCn+Vjz+6cDUaGbXevA7OnAVFojJL
+ETe2tPHulmVeOgzrzSJV5ZgzZPsY+yf6XgBCAKOdy8EKGeHoc3Yb838oQed3OJLI5/qge4ZwzKu
Ye2wpK3IDLnPey8drYEHcKyR2NwH1A7PtHexMi/Xh2fVi6AUA6X5ooClN1ODaXOi8TWoqOmay+Rr
1zP4RE6hhYmwUAgsKOhvhiy41NvbzLWAJOHrlb6Ld5RhnJ4EE+emxhulqEoZM9AmFwdu39LIF76O
fHA5PYSAvY31t7L3g99NeMDuDMc5ceE5bb7dpdCd9LA7fFY8AExEDdyBHjEBrS4UMkbr4iTvZHO/
vQyf113Ehu5uEpJV6vx3rehlLICzJVpFU3e1HGYh55V+S2mXa6xhyXwGapr1fEf6vo6uJtCGQ7G9
jCTBbIhewlVTuqpPxOOHWR22JqN1b3spvHipn7YfKLaIVsGhCKmoyRoATpIkdLPxzLGcuHmwtpzM
nZTa0+d6y7JymRWfyDWLjrvS9qqjbj6QG9uJBjWn+rzNzXUuCXZ5C5kA3dnrZRaMnGKbWuB50wkT
rVHJrSTT0tAhBbZYbNaaXDpfQIwRm7n/xOcA0pZ10VtFKkMdm5swVzRr5ITroO/VKdfnygxKPFEx
Nyj0eNA0PR0Gsco+tb8sSOoRsv8FuVwxhnphzisZmaJtzgdP/dVNtDqGy/3b22B01t5loWmS62cV
RRFc4IAj6am5hnDpXvGeUxWfrY2QUqgfSxO0h6J01YVieJZLWD2RH9+iMyoVCHCz3PceoO3Yz2KA
g9HtZ/v9iMmla75amgnW5drLQed1gs+YnRYqcZYwqbVxaAZh0/D9moHUQ6BHa4Cus+jtbt21HIv/
2UbDFK3O82avWWWYGAxGeLF25yZHfdmIG4Fi4BSPGgtKk6dFhEPzzsyg4GwMUIc8kegXjmr9Usxh
ddc6ZZBuEihyX/5PlpjPSoO3myXdzjWhHYSxgOQPZ6un5HrtSIP3P+N651rskDC42rG/IVByuF/5
FvugDXZNOxOY4HpfrAKQzatccZqHSYBRZWGn1MJ6sPdaH0EGv+AETiqrQEdvq4wMVbdNIGAijsY9
KKLORa8oTW3IKBPeSnkx8jmfcGMG/XnZSqt3lmqqTkrJ93gTy+I5dIJOzWV0HWct6yh1aDhISOHl
OFFRM8GYMdjXN22LhjkJutiqQlQsyAum1vhIZX9JxZbXuiaCwK4DszbGckQdub1Y0wHVlVc0heNA
Sf4bdfLHIaHXglO7koO9STXuvGblhysaUyLaPBxH7jabCjNhfu69mxeyDt06F4Vuy9g15kmgUJD0
aAt4pqBOo/GPO7tUJZ4Q15zg70wXHJbtYUQAE2e3Fb3gJiH3W7eAgNMmwmJ7ejN1AUYVDkbQIhEy
ugtwHmiI5aKJURPjtCC1CxZ9aErv01Fda/cN7kXQWmkH78B3QcaFd0bu8KNI2dPLDxfpIM2R29p+
a4MrhR2umxHS6ypWeMboPHN8VK/YZBBpm1QTyleStcmZ5REATPIukUa7FBPnjCk49bMBcKNFY6gp
04dzmcdbHboP+jLUkMhPMoyvdEdat5/n8IdZZW2PDgH3tBCsFSESbsamipfLxljajOKt6cTTtqgJ
PJj/3K7ssDX0xP/p//ARyKeV8IVFRUo8lHQD4GZ6V9uCv36nsQbKXToNrGeyvQbkOOpNyi6hz1cc
ApOuVpnARZcaar1t2MjeByU7s8/lRqck+AYDDGLz2JESnT95fYgkDdl6fxZ/GE/pavfbPovKU6oY
VVqmfVo62B8FSN0W+1VBhghO9+58BwG0tT4TjWAKxMMJww+vBOeOl3iD71Ujzh5lkAJylA+Fgf50
zLRxp/cVBAah+9mX5/UDhCpNk758FDTE4hrTTpvpiOMHjIbX2lULWDNX+znIEjR4lndTlqQ8lC4X
64hG5aiofEKcFsVA3pngOwSCeb+WcTURYHjunqhflGflzG5HwQILiIz3B4HmSpMtZxM/VpynyPmy
UDQh/POQqf5nt+jIEimMPvydSQJtXC82YjtXWO0hA2TtQZuM06cfFZ5CV+7dRIep67Anl6WTJnyy
ON1sl5WsRjE0S+quoA8HhnjP/vueU84xgemH9guWrfVhu05tZ1GZQISdeM5IScsK4gnxHHPzJXwN
dLsgLghIJduuFT0qML1juYIW4n7543IT9xokqf5UxNGr8jqhL2nXm0BJ24//J4Uz86oZOuZ6NSeJ
yR5/Hz3xYVa0+ZbPggelVTVnQIuDeffJIpP12ShF5ibr2K7XugQkDXoEQ6/OF1MefBvyi3irtUe+
plVgAoJwRf2ZOdx5dKvv9/IbDUWsKNj/zLtSf/NXPfWEPKNaTP5ekv7i+64+H84HCC2qU40yzOIZ
7YU5fAhukRwCyTGD/ViXKfObgCCf4QY2SpHJzYYztm1BLk7S4XsW5KGa9WyS8ajptItwfXp75HDx
ylIm8Gl5+gk3BaRCpYQCVDGUoOskXC/waXyUEVEY3pMiGm4AwYIMXrHHzOLCaUxyUZsQss7vYXNP
fXgvsfF4VTn5hdITxzd6/DKvimIbZlYRXRKNz5xlJfpyPiucC3p3JERdl1kI6KjHuNW0Re7p7ZhU
x+LLMSdBMTj4L3OjEmhHJH03zTSMkHMw0LAZ4PBGpYW/oWAaghuXqHfbVitm27+bpg7FjZdrNUq2
mTgu/REnSpnaqXl/gjral/lBVYWLm+lniH/phOn0pfBOme5Jkt+6rx4MNEVmy+n1gKBlGidbCjtn
hABj5IoGdQ8WpSF/2smb5Z2iq6FzM7rjPKaTgiYHbLZL5VHBJv6OOPirJcVv3OtUedI0Fdhw5AC5
JoCWlA/9yM9Ns+laRdqRedElJ/anT5CuOv9H56w5QAOg/S99HNxY5uwvPJrLvBpNuetODLwEFE8+
jUA2hsYu9SfmxmlFbSN6zuDNNTx21KOOR5AWbSHsCPkTgSbHsi68kdJoDr9OjRNzaRBEYdhbskSP
73d8DQ5MeRX/m5TITY8fnQe4wQ1oi7hgnbTZafec1io2TTjNXAhL5fDrHBVAFLdwrh+2HsTrhE7S
WkQd2v1YKb7/v7o/OMoIQkoF2/jS0FTOTKrfLbUe+58DLvYCENzvPN/deAO2KiV51WvvbWqVPTgO
fEVroMjJnkd9uXaqn3v1dNqM/TT/kP3Cxbfh3UHUdCY/edhIKR2fAVI3etUTIHb2nva9urvpuKkT
W5Ti4IIew35MMdzIwxPleU8iCVgrH+V+6Mr2KDu7Fz+1om6qPcE/bFg/Ftf3o8S4H1ZqAGxZOFx5
0GBsXV2jsUWKYZx71AkK/W80AdA5eZ7tRKGmW/gChmmlL2kIvO+IxymXjqU0dUul3qvhwVzJ3JGP
pnGeg9Desi4/eWNrT+aCbiNWFu0mTJF/i5CT4a+21Y/sNxzIMUV++iwopKrLta8GxyoNL711gnso
pO+n0zK/mMCcgFTGrbP8A4RKnNjz8VDSS9I4TWeVXF3snOzbjnvAEl3Q+CsyaErqM8h0A+Ef2jOt
aKVYfq3PQbAgZR8dK7nBOG1j5lO/uhfNjTawlX/+AJGbh95zSBOeJxPFGIP5IpYXcbf8Hn1xHU8/
js1/9TAEjqRqc6IeEvSIfrbQUDhObHWHTXl3UFhvBRZDmIMfakvm4BynBdj8yaFitDInJfH/7dLf
an1H2OEiCZsEPKKb9Mr+0DVtC3QtdudzPotlpJsbrMWg3or33ScDFw2fB7+LNb2X1ItKVfHp1k7q
1P17QU8Pe9qdQWptrPfr6mDiqBPYgTK7MHZ2J1tgO6veM+LVjz8vOD/Rk/sZ3memgHCa+ZJLTRVU
uVcQImXVgZSx4Y2r1kQRbgGLTTaOaRl8ooqqewfw4jW0eCQcF0qTvwyn1qCp4mMFX6yfYBa/i6ED
jx81d6Z0lYmnR2arihSsq+bDb8xaRpF3THjv+JlEXxWsWHgLpOVJOXO21y87d5y5YTntV6/PMVzA
OOrzn1ahibLy9sKM/bFV9Q085IUEXZflAgO9bm8QfiITTC8gJTn7pUhumkhnqqz2XdPQxe7CG4+l
21PCYuPsdkGQL8ksmT1T1hz3eKBhTFKESsrBMXq1l0aa1w6LdkeGrsTmIPYxmFG6zlWEXVKFAx0i
RxJtOdwxY2E8w1fSiPv3tANg6O2x37XraG0cxSORON4n/JaLurNjD5JRdogl+WCr4U5UYNaJsDVd
flnnb8IxTtLQEp37k7FMmUo+jwqJ3fK3ua56m/1B9F3XEMqWS8rbzncWQiPw+DdZmg4UOn3IkGkY
mUx1iHrfr/zWwPVSBWHmkO3v4PENyXHKQJh0FBVum4rsegYCHq7RWcgC+QKhC773WFPALpOl/NzH
Er/Ab9+jiG+feDAw8G0hFUUg9WFzuLW0FDcZVLNv8Jru/Fj1nmaO1yiu7xtenaZtDRFyRHTAJF4t
UDNtJVRZViGJIEtVf/YJ+C4EbSU3ITSflW4/mn+UJW8ELYKo/qjCdzS74BS6IQ6npX6J5PjCj1zU
dqIU1UB5fMbHdOuyMO8d2TORBMtprbEbGQILO9QMP2Vrl0LDhbY+iOj+9squPRbQRhBSEtv9UsMg
PEvF+6om5FYATpfoUvS1Kd25HvRBEULDodq5cn49810lpppKQ60OYVJAs4JaSdIo6ZPKeP3QD5SW
gjaEMPYX04FwHZUfgmFSxaWUXf8mp8HTTHEZUa8Wk93BdUJx6481szlUDdLVfDJgQwOEykR8cwlW
eHXZiBWbHfEO6Ht6R1th1EV/duQcPlSYW2t521YwtiQisqJXdq8ZFB9hbl24/BEf5+uLUHuufDGE
a+UMMo//HKJqdvbnlYEfM/WpJ5/oesmAvPuiYfU7IIOeMKpjlgCRn3HGZ+MaqK/qeOYrHBLdOnU0
DZDlQAiAW2MNzClJYu7smSpJKHWi8anaXfdANGebCIw9JTqaHyBta/uC4XzFqoXJ0gFjkEdFjtQp
DUnoX2f54DYuHxYOIXX9YEAAj80OZufWV8KkAFWMn6TU4jMvi38zLIWer2pD+LzeBwb/nTdpwxPD
rPFUfuTKy1ONdvYmgBaLEgPkgx/PSQAj4NpryY6BeaUbwLAjBpmOznDZStwPVf7F4Dz5QzlVlcGm
TWhQcTQNMT5rsoOc3fx6korfc2qVGkWcl4GMgOZ9pYDAQNoP5CicY1WZKu0kX4FCdJK4AE64CO/y
feayXCrTPxZx1RqBX5tVTpiEnk4O6LvoSNRyM9JerHA3lYmaKPoiu01fqNeyiwxSbXh6xFMcmjuY
n9yhjWpYIJxTXEd1wPNDBCD1sjzJbcK+lnNm6HkqeqnqNaMtgnw3GHhU6FVJDueTdIkzbawmM4wY
d+AinhjZxG312a8Co+JR494R4715/t5A9hVMUuBBQwZMlyBdrshYTlG2xmku2K3f5FutEaj8zFJv
e10AUl/YTVdJKCi80qagglOe7McISBc4ppTYF8KV7IJUSsVM9L5cLtfwiIFowQXuxvPhD7JNnmAU
G3fH1EmjZgZmARlY2749NFAEE5bjPK8EFfO9G3PZlaSOWj7jK0u4V4bWPY6T8SP5/q6PQRfV/z9J
82g0s4Qtxo1ELyNBn3AlHuyR++hiymQjE/I3P+pemnx/HWhxnOOeBw6RPY/vEQOSKhNsV5bsn7zh
ogGmmL98LXdhdo21Hj0r2lt1VQVxpkWqSJKD5lDbmIwalyyx7JLhIdb0SYi6MqecXXG8LhlhHaU4
FGg/j+8W+BZy1Vp6PjGRqMwEIrJ//jBiGXxbZArtPvw9hgaMcrm1A+DDoT7oQU2DlV5nJbfhGS/9
bNK4qL/5DtDLSi/m4nzYhoZtcypvUchkaq+wdr5R0PdcEcSzbfRo5K/lcJHZv1xmSHaX7XTo9758
gd3h51KWFcGPaz1s65AdUy/c65o7XfstJQY6OYqcPKF4Bgob1vwj8QvzRnwm4jnW6wdSvDd9P3LZ
ljNRMnRjH5Wye/FZexkivqrw/nAcmep8tMiwzSfdBbWL8VtqKTQ87qtJjoA/cG7djrXX3dAOTRz+
0jTwMcbgiLjSXK/oBJzqGstpnuRmCSLDEhyuUtLoEAl6dwBozJMB/BsQTWEyv1rvHDoPsTeX8Mql
0110DaMCfNzp2jJEjMggIWQe4WtbMrjj4eP+FkGzasSvNbhV3jLNdsuKd9/Ny8EmQdthOjby3DEf
vBrVYXek2/0Ix2kUoy4gyjdpdi0iaJh65CSHNDjkP6MvrM3jmdPd+U8p7cc6+DxZvIdXneVPgSnR
VEr/xVsKANK7D1XmS0LMvLsBiHaWxI1boVV2XbgCUeNhLzHpFYWAdM4mxGjex1CvkZ/V3FdKNyNq
hIKnwnN7qpkhudzOe3Veb8SJPjCzdLlNKgfGA2+DydXhN5Tuu7lLQPzHJ06M9/Hz2/jFdsZ8rBuH
UsFoNwdpA7+fWQcUJ3q+BC2tBRH6p7Ax5xPiwBBtEJoO+QSwQk4PS2iWe8KEi7AKjoFYJwtOa6SQ
1J3IH1SHBN4t/5cXrvy0YK4LeLhIgglQVUfWfKMTsWpB1aOKJBwBKW4EWESIpP6MCfZ+2yll4Ro6
5IULcO2MWADy3DofPLQ1o/jY1j9wvBZ5dYcX5L54xojzZG3dzmBDKUsGDGtCQl+4An+eUMXADai2
NN41buIxUUwBUSeJQ9Vj2Hn1HuyKo5RPAdaJzfMVTU1urt15JJs59cd76aFWe/uESropzf3qdjNr
aUlVqONNXGkB0h9r734GIZ+8wFd0AWLLeYsikvOZUjcNu9zNK++aep24q/cBJiuwZNMW5fQIc0GU
VeFYkwMisz5E2zydHdkEdhBq//XEoXAh5OO/5xglGobrK9j57dgqtCwoODiQcZJHnrf0/afdLPl4
Esrf+650QJebXhzPyntRN+de0b+MAm+fUPtiNsetFIet6ox3eurDaolY6fbclf5E4R9T8QzdX+L1
ggl/e4WK/hTlgrAifkG2eucw9/PVHb+hbVNKUhS/PqnH5hzJWDscgOhNu1wZmp1OrEZbg99F1fn3
xE54nYdxda+OhYwvRADYC2RxHn2fs700KDX2A8aNeMvglcZTV3uJPRvwWQ1YOI5zTJG6rFaMBFim
RimOWY+V2NW5jer2KPnC8e3YFUydhyaN17OfPSUgqeoP8+LpYZQD08z4/KedUdzL81nNd74VQwBT
BQ0GKN9oYdOrqwEnTWXLXGk0uq/dLViyJaU5dT3jYXxKiGp0N0+X2rLvwbGAAMa9U+xgCpnHxoRD
bzvukF/Gy2Jn/G0IF3tFQUJ+U9nkdsRZgwNzHp4E71LnSj40XoLCtjAnMi2wxQiYtTQTfBWprZxa
auPx5iblog4icZT6Fd8gljp3Doh9kntjqEX6N72cMGwlG4cU/0GAnMx8y61Ug5jv8Ybk3OF80sJb
rdazNC61t4E9fCZU1FbmsFtO/3SohGGpch31CO+fUD7roKhUfxkknnYvoD9Z+Z7dRVZxVhqKbqxz
QDeorB21av6lEIlQ9tmDmdUz0MS2ZskIAKd0zlIkzjkWp8xmwOt0pEqttK1WUfZEHbuWTzLYHPrL
b5+RdKla03/smDsIIjj1Ui5vzrUZu3lLatHaZO47xiq67T+RpRTS4jBpDHe5Rls4zvRrCqvQHZ06
KK/fRTLFgEp52TLh2Mm0U2ImVBZIqY7ZO4vNJIcYbNOwLDEBqAAzTtdk25XNa/RRIl+NMSkPoXI3
bX81encrLcA6PDvBxsy7TLDTF6392iomx9MvDW//pLV82xXc7x6HA8IVtfTRdvmBUCDgl3eW5DuL
3uq+NMyE5OMPA67keMN891GAVJx196H1nF2c0RGCxoGP/zEvhTxMhPh0GjDbHuE7kC9i9BuIfbgg
QLY53U2qYsZ2ZH/KcwOlq46mnWVbpPVEhrXHXpMLiHrSm6XOvzMF0DVNVLh6kyQZohT9Wxy8dk8j
WCEr86I3RrAvpuWEwDOf85difHrEfnFIs9gKacE3m9R1n3GcsM+8GRPq2snMKGuwp8e/3ZKtgGkX
5gr/nvB44rAKsO+q+rFUxliiPFKUgD5gM6z+pwAXX4e2f3+nTU/KgQH8bFW/pN0BX0YFG6s6flnL
BFi+ZuraZsqv9JtD+sbHeLhhjBxDSFxfJyQ52iI2XomBPboMO+pPqQNW6KkQPqNT5lunHBKkz/Ir
59DwE/QjJeIvqBU+WDe3EZ1XAbbMmLPJU2SJpYsCwLBePSfBWlJPn6m7D+mpnEbNGL8XY1xUMCcQ
863XvUT2vfd62kw16UJXPvNZ0XqZEsHLkj34z9C8KHPIZ7vBmBW14Ymz4AUoOhLtexFks2Bjiorq
1XhFVcb5i6JgEaLMDJxluGUQ5yCBqZB2zie9UofgOkFLrt+kT3/uzDn0KP5j155rt4ZOEgS1lhTp
DsNf8Oc1EgQBQBXUceWxUD8ErTvHiQIP1OYQljIzEp8K8QWKW9MLpRAQOu0dqZBMdTXirQAhP5lx
qS70qE/eAVE2zAnmozwPhgx1TCp1X71WV2PDSvISYHJRpM6vkPw2K/c2O+GICRIu4MCER+R8D52t
ULNtCcrzWxQrpxgGo9lC/+yV851yhgEsd6Wj0Je2cq6MXryQS3iv8wNI5RYdYc1fKJr8V+iSA1+f
l/lg0qJ5r0dCTEdSlktL1c3NrkT8gvT8aof/lnP7Rr2wAjr8f4sQWfE6Xh9yZWWpYi1wBfOmFB20
NFF6g1hlLOvwyHdtP0XEcaanbjkN/rPdQA7aM/p8AsyEK9vfpSgLiXCSoSZdMzzK/jpFzT/PaCYd
eCwTCc0jvoohZiClSoD0rNZdu17RunrtumKlTonVGGQdTpHP47W7Rts3O5bX1cHdTZTpUDiQET5Q
Y2YNc5j60GFjAVvEU8Z9BdZ5d/LJmnzO0+XQzEvksKgtZeX/7gXMlSTBsUk9KPGpYIdocXkLN7/q
hXmbxLJjqIWGg0xuGBpyxeONml4SE+8/UppsZfPhxQrS1fK8FUYuVneN/OA+ektva2xvYYyL82cA
PBpYl8jnHqXe0P0aD2xSdBk4y5Q2NWjhIOJMnj02/tQyCgmfZ+Vin1/gWaq3sbrD995MyRHmwvzA
zL4wRP95FgLc2L7OiCq9Yt1hXEyP01pkg5fNNc7HwoRn9W009gIg/Z/ATR9MoSD+napIZ2WFlxE8
Xd8aoB27rltS8VowzepeU+d2cVZuUM1VVAl8PEWqP1Csx1bj0FYycGXbaqbO7qfF8IgbHSCY2hyF
EjtPR6MOIOVOz1s+8yHf0r0x4sHPCibEYivfO48E4+WAfub3S+wWnWEoH21E/2QZN1b6nvsPzHtm
kC2BuuRDEn/gY9F6ux3cBT3lThwvsVRzenf4jweLw3eF57kvczUAjknRolQmEPitD9+xdrOslFrr
2wvZ4pmB2lgbSBK78ZjK4897uNwP+PemYc40Sfv2UsJh5vIF/sTu7Zzx1GwreEayb0RJAmaeJRRQ
V/4ZJJxfPoveqM3NnfypSx78KTTL/S+D09nnxbmHzqM/ucY8GgkFu+orORS84p9q5dsxo5KJQgqr
ORiX4CYzPFSC3+ziET9eqHguN16k0XNQINoCfRSw8vyOhmB+vFoqrVEmC6AWz0hTGXTtZQ7NplHU
q44TVMY6ud9I3CNpqOb2KxzRtQvOgkTx+x7hxmN+RbYvXG6DhEsF+PDvFz7Y8Rb8r2gDr2RZNgRq
Ps9vQ7LvPwwpSCew7KdvEMh7QOQxbMraQ72XlZLZEEW71WINnde2iNLFACV/45/vGpqavyoyrD3w
Ejali9zYNXH21mEaCukRnfw9+G/6dcQvIX/TdgCHutHPdZdrykhGShpSm4v3ZHSEu2IzvHNCVdgD
q2iQ6KGOq9h8tqGDKvKjSUsiNr3gf3usCzlpT06mufuVlWwJDsbFJanZHKg+7XB1L42XLKbLjN9a
2FJr9ufKF/cIHIaESQXw+vBaVRX7jhONx3hThi0tZHGYC6l/lduHvKtMYmoI6byWVnKEgHQXBHxU
ksWt6LF1+sgysdGrwgtNm6Tz2DkT53v1eH5BiS4NEeh8sRcCPsoAmdqWRq7egJ0gQvZ6ytQVhrLm
vB/IlIgXdR7PE2jri61caYdEzTtQl+bU3KkjU6E1wdd81gyjjg1Hbj8HXxRszygUrru/IhomwLho
LYHU8yDXzRZgdUcrdJzp6CxXFiT+RB5zKsRIXRBhIl8W3LdzNJyFslZWN8baDcY3vXJAQMcYWRrC
BAZEaHK/pxEsSfxw1Ip6w19IcaDh4GnkfHGot7OUspEWUY071v2tQP4lOeQ6pHtO68Y5XeSLTtYg
+GvzHxpRHA+/4DtzcmMsv57cJU7lIbuAr6GEQ4X1wGUTJ4P3UHrWceGba+grlN/I7A+OFPju1R18
s0Y9V8xAhZP6NwmqhAPeNuLStMiMu4zpf0sz+IT6unaXjv1Bldrpn0+B67pLLQEGvM5BBWm46xEe
7ZibhdxuSpQa6Uxzqd787xWEt22D4ojyoxbsUJT6cR2dAa7cGa4awZhzJubhZJM5rnJ32tsI5dfJ
hR9Yeb2qTLLUIkNhg4wBWrYPau7CJw9SitK5Tteteh8902EheZAf/jH8dzqKeoYtS0xPh69TAQfV
FTL1LzeHSKGf6MtbtMeThCPiO11EUcYbQ6V1N4w4VfjhWYejSu2ds6I5SN1SlUsfmMxq3Ts1zmnE
Deo4pZj+dlkR0hhD2nVHAwBt1g8g9LgTKxH3nXm1cnMmn3O15EqMrMXHevxrYeRTfU0MmvUKC67s
YH3UUJzsULF/yXcBWbaV0TskBdou7Latbk7YRB9uln/E+XUJpMO5u6w6KXABDpMZ7YZ9PRbXcvuz
HQbosbk+hPMDJD0S6LoZHoO15e48lLPZRkpiRwrMSh6y/R/f4kqzlktN7da7piMhUXOp9t8oXHMY
OF7bd8lB4RtP7FvFD2qcKCMoiccaJt5yKZWJkqXlPjQkD9nGfGn0VqeHGWVsMvtjQRxVOEgwzW8k
w7DBR1PwNHEr7RTAhFdysiLXpJtvUo6wlwBT5bPqXsyS5LB+yFBBML+M0l0T3TNiyqhVCP2J9ty7
YcgcXdclG9zChEWO6gl4axQ9s86EtqHq2pWXEHNGKbjKY/mdcDclsP7OA/1BOfIB5wQzaoBVnxIY
67M+gnM5s+NEvI84zmv90I9u9MD8vfDaWUvQleu/Zj9ljOB/yJ9RrOVG+S2/dJm0r+GyjhwB7nRt
wwn2anLHMyIyDFUmAJqVtm+XbeWlWZ1C4CLi764LAaHpVdWl/wp2QPUa/j+ws0BF+Cuw+laXJ0Ff
rg8wgBHsPrKWHIYW2y6xtrx951dAtigE2ElRzf4btZlZngY0ynHlW6szXazgYPFsBQvJRSHreaWl
DUYXPwsI5xl+PbG5Jq2nqbIvPi72rZ2Pcg34Mxl527GeitjpE62weGTO09sjYxpmqYSBtjNg45Os
dw9FFgR74paiw4OGhCC+sNaEENn4B3QQSPAod32/QuqijoC0PnSCiACeKopnmR7AGnrv7NUsxvlo
a1xbJG8pcvkgwr1pENHr9czuJ0tEQpsRJHCoZIymQ95WTwmP4YMCR3HimNbQ78Y+kRxt8l7Sv67+
4N5drMXwYot25AzPA+CJfAlJJsPgiD+HetK1ravbD+3W7smmW6iZppQD0DO4URVrOcb4t01S7nB1
uvj+o+jo2kmRIjCgM9EALDcKJjqQHq9lFPkfL3C0rtKnRGL1irLNvG9Pd3ayIuASBg/PNj7JM3u3
HwD8d0LhK9wvQ1cUzd84zqga+xlM7EVT1BvMe2bnBXFkO5bYBarYkHirhLzCxnGFExzkx8X4aVHt
IYiZc0OPwfl1b5ViCsNKEiovMeQ4dTduxjbincrQmbFQWb+R/jejIGizjiZO3MAiFvxxkOe22RWs
4WKrD0oqADlTfyG7euCAhgk6XI5SZdVTgwQ2516O3g7CZk4FNtQQdxTads4h9PILG7qzgfIHiYQ3
yQHoYpiBkhisYGfg+GyuXEJ1W3p+mHmt2bMop40R5Ug/4sQ1kiiSIWWnI+oApF1XB91sPpQSQDw7
ftC1PiKW/nuz8jOoalISsgdBZB8i8mzcW9KPzf55xtXfCP7DNlSTmN037uCF9Mn/q4z8f1xBMB/4
6qMNKofOOfPQq26N0wgZ3H+5pgH55R/q0xXexJ4Gz6AA4RgAzk7zpZr2yk7Ei/h604I686pHTHsR
5xL/i4cXIFjql0HMUpI26eQd9KP7Isdc5apiWijvVpgA3pnUzGjl0du8J4Plk8wwMuhfgnIMIJY1
+bQokUPdw8/UTTdow+lkMQL1dYhheBnnO/tw/kxlbBLUzMzyBqIPYhbqrlXDQS1TdVXxhAyTPLI1
/xS1pDfpsvh2GscmGLpFWnpEV2kJDn8YVb2diVfHzPMBj/Rzzwv7MN1LS1/4XI3h+nwfjMcvr0wa
+E3HUYstPCDRcypsIcc4ky1cN/a8qxynQhtCSPpb9VF0lLfHXID0tNVjB4MQzgocA3OvvCkICRM+
5LfxkF5dF8F8GCUXEJwcro9wdl/cR+X6yZTNYfwt/f0PW9/21+I4bRrWTH0fG/Mnmxrz55XdYVfm
lA0d5y7xnka4+WQ64poKH4CfV12IC1My5rSqZVwYe+Yw1orDfBNebpIJ8Ey9BGIoGenebOZZrMkn
wu+f78mkAOr+AOgatQudMrszjEv1vFV00qHQ9M41PmGtfdFvXQKYL6EgHHiDBGvyrPL1ncn9PdX+
aKH8qfPRi/UzjeauKWcp1DwWahJGgHefnTJwZqfZ6hBt6wTUM/szi/F6OIxIA4j6jJysgaef5FrV
RRcfqajdn236uM8axncWY7e7Qz3Tfk4Zy13/0i0SLaVmG8rwb1rx0/p3hwRYfmNhNY2+HXZPKPlS
hgY60Mm+tUWs0NHWgOxmAYxoxQvpDRF/SrquZVPOcwDdFapXLERUBTv1/RSGBrFx9266DWpBDCQL
xvWQ05ZtFSUn6V77b1K/9m4cHOisIbiYe2Za3SjKqYRXCkYbwuj24esIlNXKFroao1Mp2U8dhhP1
Qe7kqaxjQDwZi1WUTwQFQceeZ8cRQayE9+Tsrs2Za+HFTFXpgAPiP6hjn7WQk3Nr0iHJMVMny+0+
i0ZUb0NLdEeZQzzfqaT15OJ4IydsP4PRbwVAjHX/u2jaYUXX5cSvCP34JYQCP3n61Fsz4LzrhvtG
TG1zmWGKq0XciWCUhNTkVQRFRONCBk0CPfLkJK6C7n3uC2F6H4FSkrZe5ZhNe9nnlGIcHl71PUDa
wBvfOi6dITAsnntDJzC5ymOpld7d3qVEg4Q7zC2YN3VABfaleEJHPjJ3WjrxT4mN0AcfoP1Hpygn
dhN9QA+GFARXLGTGjKmAFt1QfADqF+Zp+ofV+3N/fbtfvX5m8TeovAJHUDiFnRkv1q+0PYt/CuSL
58yobfT0p1Zq6Id6VruFGpxuhmgjyn5064V+O6w0e1rjyC5tS1ZBWVriv9ak7ZKVGYZBSqJTok8T
WX7Gzc5kpZoZwwhxrkkqw8W12209RDkgHCx9cu4NxLqmWMDcYSFLUGwCnhGTK1cmZqG1f7o92MKe
jo9fe7MnkXmkimJC7pE3FM2JQj4tK6zq0z92EuWK0RiACLIaSMcASUbjVsjM4sa4h88RyFujdRBk
HM6Sgu+yA7fs8hPoh+u3I23gte+HRz5otGu75nzEuFN7o+A4BqLICrh9RFDz1hsMPp+SLD1Pk8hA
7AFZRufjc/0X31jrCii/ehz1WR0xGngXFG8421ZhuMEfmWaXFQ6KgxTR1kCGlPMaAZk4aPPE9lCH
n/NJWXfeiQourRyzqaCacsKQo7VVkCt6s2hW18hY9j0dy4Y1ES1HwqlrGoYfjDsJs7Q5XbaFyIA9
WGRxKfI4tudx11PCRQjW+mamR0FAojNhk/vrsQJb2GoY7VRXneNzV3dAaGOLYCR+Wh9fIWpLITiK
Ou+dBWJgWZeadjGgHZbLT4W5z8fdVyYb7/EcCGDc4fw99IM7meFx3olgnjkEjBab/g5R5Rk3lY3c
PWdJQc22/T2NTbTNfHpXrIPkuuq7JOsQllkwzC+yFEg+qt/dHRuaNEZAIRFWEMGrEe40DUXUXFV6
8FbtTapbgoC0be3qPRG9iqV7viNirCqt8U60oxvZhJGiREzbZFDqETPrGQsZw3KCNBm30tz2//A7
qX8iXXi7KrZJ0zT9AhHB0WqR0bdjNuFnCAatT2y+ZQY6x/L7btP2tYo5a1h4Dc92FRYkchT1MDNq
OYV4+4pxXE/QopiRNPKlq9TFScyPdMXc2faf9wjKDVlqDRM1Qw3ztn42OX0PxkA3GQFbMOyLAC9b
luRhHulv22Y2bEuosahPWQXDr2k+oxy7Vj95+KsVlCQzt1ZllQubkbe+PW1GOiio/yvwwOa7O68m
a5Y5y6aRwjeBXIz83wXpy9AW1cYaj0ul1U2nvxP7jF11irfIb8qwgydiC6iQg/KGnrVSx44inMIi
9gES9HdTv7ARcRWSgy7MfnCYM8BMFKZcwrMN43Zof9uYbls/Y9BhMCMWZU6AXH9IiWfou1HarqXH
tPZwH1FJTvnlT8T2R8xx96gPnmLv+SnUlXED0/RgskbHT6NTGqdp6dqkf2ZCr7F1ipFzDfAgdneg
4/oOuZHaHdAn3BS9zSTbxNSJeE2MM7S4KGjScDfWSot5uED4qjGp+a7vSd8gwOBQkVN2oi5LDl+C
dHUKEt2dL9Z4prDbFpHkWvX2MTeIKgMNDT1jTCSIeYGOTGNVRMZwUdWJE8GbWa3jwqF5Ee6h1aVq
91/8SFYQsjjKFB6/AbzjDKWnQs6pFibwhxGAPwrXXU5uLVdS3bcrqrCUrxAgga0GywiRzbBMUXyF
3XRxx+Z1/KN9lPrYYU4qyPDv4IsrgEBuXP1552hMHGL4ul3ZEMmFpix6JYHZOFIsgXWIJKkm4Oec
J8zmNHLPQ/6rtkcZxQWVu7FwuZ+rMN3K1/HS9qXVoWMErkmQGDb3arZ4D6CBghntj5ZKAP3OnUDg
T89hl5CAPSo/VGCooSHsQgemzRVRZBXgx1oSgjsGDxtM9GQDXFN4sdEHuZID37Npnc96vp2E/MQa
Qu0l7f37xQ2LMqbiFjvDgQwQbBeLwBgtLEPVpDJux6W2xsCEUTlcox/1sYpD6Wn5hs0MifUAuzBZ
aD1SzWpRU5KVTAQ16DkhLCkWL0/rsCwTPLiR+Bfhe74Y64EZSc0bf8ANfkIubUmq80ob/HyfnBtD
maaxeKml5lmlY5sFA+/KcEO2MRDLRB9QabsXM6lepiro0xqiibngAJSzhS4Y/zHnema3pXQF9rxT
7mCnMTneG0Y0aEGSsiwK+ssFBfm3KrpllY9GtNqcK+uqb6lmIwTIwfB4Pe0wYif0ZmBaGKXxLNHh
IICyEv06c/jbkvfFz77grZvoJ6QjlOBxz/a3bB/N2C+NQJXivs73um68J0OpBxF/vAUXFlZF0740
KVI1hWaLz4tKjBZWOFMnttXGzC/8CXq9f01N0KmmIOnQgHjlS4NPiq6La7+coC1T/fV0eU8/Eshv
ezc01OhiJq0bHeVx5X8DELjDJFhVhHGaxEeKzlc2k97O3sBK8Gzl/ULZdoEC9G1eCM7cmqeMhOYW
zI4yut0xKGzOrLv95YiwtBnziEN7UbtA7EVA66PqShA0p6Z/zMjfXJa+bFI9HhxMtTqVdDVJiWBv
v1Ydak6irQh9/re57BHmOxw0hYX15urQTJTsW3vO/RhXPAxBbq+3DxcaHZY209BOYpJDV7HecPU1
7r6aOtQVEz1D2H5yyMqea8i7guBFc+a4wgHXBBzED0J3fm3qWK02QaNLomWYYl1C58nVp8XaQNMr
6ZecgwzrWRvcJ1RdQvPXs8CrInlHchpmczIroiD3C2DGWBpYInaCAQGmEa1r0XAIJIkTkWdcO0L4
EAFhHjiLTj4jm0jy9FSy0Km3daJ9ujQNGI2Cmiu8ry+n5MADx8sPmt6HE+B6bUwiuI+TqdBE1az+
RsLphDCWdXkWq7fBnR6V0SPpfyrqQBZtzEGa0E6holFfa788ro0S48FDR9Evr/6/y/MzNX9JCEny
9t71Zmd3UWXmDaXOC82bffrnlb5AjUK25895+TK3NYnJALrc2ANPoSRI71zD0DAwZa/Fxs3v8JD2
2nILTYEpCCRdAHCWbPtWDoxGgYg8/sK7iJrzUFUdGRPrYKTg0r4NdqJVVt7iUuzTYQnc3BzvP+o5
FBgFT1DyRJu6UZ2leJsWqHhDXeW548i0SadR6HsYCqqXbYI30x+eu7LDXTO5pM56dMsghNfbINsh
bgVbTa99jAjszNMwVm0ggVf023gqdE3/vHvuPAbRcW4QYd0PM0aYKGe1cUXl5NVRfvTnKlCUqKzM
ESF1aWtoEtEREt9byxmh927VF4vBJMWaMYUAhcgvZKjwyQuRaxxBsTbXMprspYzaJv17HIZ3+p3+
ZTp8JJZJTknVjTDFupik7Irz4WXvKY+mo95nhGp7kKfExLdJiEVUkCqJ/ZXjJGW8mlZ6pUvuuU1n
eQc+hTCstLCdXBovOBtY27i7uh6MvYgGZVKR2XWVA+1L5uwTxU5sEYYMXs97ZXg6JMuRFbnFSNYB
bdIVr9DYZscrI8DYoVJukRYLYz+GLgXhNUJw7drooJTGBW3w9LAMWb9n6+wftwKrcqFGexTdoVNJ
RLWGD5ei7H1h9QB0giPeQpkn5sIwaDQJdbEfWeZM7RSdqm9cDhoBy1NU8Oxk4Hyca6R9Isf4bTR1
Dn8unoPqXfSal5/Ag0YX9LVEsWbYsu0cU0KMedFGxvJPxLFlX1cO8/ngpiP5cvmdeZEnTJC1zXfz
M/8YF8KHmW6/0gZ7AiJnZSpNtsA6+cspmBtoFKSBOJ+dqMXz4A8JTn0KLEAOPQv+2CJmUr8hy5/+
O3+TEMv3RGGuWaQENk4W/oUd1GKx1aQAuFrvLl/krm3UEtkj91lhEzIuKuXoYK2oKPY4MKleuxVD
4Mdtg1oI792WAkrf1eOZF5khE8VZue09OgLsUmpQk6ycEicVXXUnnlzlM5pGyUul2vHiekK9ZkZp
kgZZSrOQLje82PfheN1sCpiwFlKiYK15o9XJ1LLetay0Z2QdvMTp795bqAibcMGnoQ/tkjzjHqjL
vX8iSFPy3h+At8Bp2MMrJSdy0Y9XyywhPCzjewpcgsJc61h7yQ4z9vwpicNp7QoqCjMoKV8s/vFG
+ZbmimRTGKnMuM8sln3QGe/RDxj8IJTooEHjhR8fGTnWSteJ18QKkwQrem3N41c9mhaCsrr5u9C5
VBGowHfycSU37/thSaDzkb4jEjOGHX8ojwewtYz6iVtYjKRv0UFy9tjmJZ9+F5voGt9KQE7i7Njl
lBrFGXz1xDc7HlT0rB5NalIfud3Nl9pjEhm29MTJhEhfZd/D0BnSTkirdPO4AHHB/QYcCzVO/aja
y5fOIDqBjwqVnjozz2kSbQuCVFr1j/t27sIsDPAGYlE7ygu5UaUslR2dPAo7gFEaGyl4rcBQZLhx
EgAyFUl5GJ1fDX670NBW/5iwE+o1V5r6uMVHq23gYEU1YWn2AhEmm/ByDDC9vx8j4J9IO4lGGLbF
jhynJfAwLGxVY00sori32fGSQmphwxj25WLQcJBGuuXLzwghscQisi5EP/Y6+l6aImswCbriCF1f
G7uprNy4os58uHLxk8XnchuA1/ShyvRJnakwkZ57DxHu4MNRKiYrjVw937tD+S7gHyAT3PHdqrS5
tql47JHs5IFOb+mshvQJ65gInFMGTt9kNLDbpPHa4JsHMuEFI3WzzL3B/w0FjHlaVhTCVm0iNZwZ
2ic5YbzwMLJ/g3M0PTnSWgyHZbkfZT/JfWQYfmgR+it4rgHwoB9w/dRuvvsJQB0rENl38CSUr6Ee
w+V8OOo8ZWFI2yGg5/e9j/Svuu5hDyD08MVaNhpxHdc3Z75QvjddKcew7cJPRXispv2iVW+zisdg
Gl2hgx37HKjT0xbJMBx+ZBvKCZERDjb+90sAtyIjOQN12gVGHBarLr+kDF2BHNWBcUZVvaNEnIBn
oUGmi/Krkr05twpdDwaTX0OYLw4KgmJ0t/fGcFFxLJNUcMJGg2LachRhqry7xXyKLOLsvMqZ1bfb
UNmbYIGYcy9LK9Un53hemA+5rXuNoqMT7L5K1lvMGuAF6Dw+mTaAqoVoRsAr8vbZXmE82YqVnptX
MzHIBq+G1q/Vz8IjQUhF/Q6nlIh0g25PWpBDkd5NZVByqQIYd2JTXjhVQ8Ny4X1ZVyUFyj6GEUYL
+UKdnLlX2+SfDkShmdrgGXsobNc1Z04ayySYCwKDdjwqYxuolF12Qo33enpu9ILp1htFlL8sDKTM
Dh3edVPDsfixWNGwi8qzouiZWWXL1d3Lhwf7Q9SrL/AJrnHamJ9dbOKu3OvPcgxAoIf28Ty9FE+/
2utgAP9/YPkLnFgKskwTeFfKHtFKnzU0W55gQ4ctO27AAeAJWY9IDAme+ezhpqBtH9sgaSVqd8h9
niQ6LwTojTPS8I4zcFlNZHUo9/MFrxljwiA2idfom7xiGdfEQ08fcMDlkuoz9WwKuwrK/vwUrXrn
Y0fpFNXqDx8QBUuIn0mvTEB/3FcEu7faLpbZuSHEh+ThqB0S55ZxIvbIGtfR6fWj6iDMc+Jq6xV0
cKr1KQ97MbBCYtz2z61FMQs6JOSTI9I2/01X8tJWr4FT+rze39uTHaVXOSX/rC8jBf8FAS7lEerH
66YHaj/KcpeUUnruOrN5BNjKLxxN/8i+Nj85xCp67wj7ilr0whzOh74yLW2FeX3sKAbbQ7AxmU+7
wPlXHmoIfEdPG65FDNHQLvAhYr/dXzkG34Kr9JZtPgTOXS1zdLv0pxtdRlTYNi6mrHp2AToZ7/sY
2mPUZZSNFO1pOZiTaEjc6NPwgUJZ5TzfkWH9hPJ8I5FeQWKD9DMxUfF2umvfi24hNMPKeQ4DIj8o
sIDmwO4ERcqEymWInNlDkvuxnx4+E6Q/7dJpwVLveaPXvTl1UxAoxNKjc2dT0DjnRjogD4Cir9dp
EFJddY9ycQLagRlg7hvwqYsO3V4JJlnySFSVVCWI/T1B0+OhoYOfodIC2hOyU3KtVvH3kMMzY/nc
1K9npO3FzeLMrHPGg4OuCldBZvpKFtNaBQF1tT07KZ+be0fb2hSfba1yybjjTo1W3Vs9P6kXVRuN
VlbvLx8Z+pY4w8LNa9ZhwkpVeZyuKwcM54wVsbQjgRDR2saldCNINMWgp38Qe6l5e2zDTDPm9Pv/
cgrQOm9LA2qmYZ1HiF0Ad6EP4RURiSrj0l6rYsvA+H6o8S8m+pwThfhFkx13gB2AiDHlik6GmIeW
XqDR7aCtsdPOASwqJTielKm2oRj9WJoWAOdcxi75YVFDujDRSOTHBOA5QZ4K2X9nJKMKG9Z1XB21
KbsPFkt6tEGZ2NzjIj9nQ8JYGF9DO6fum3wPZw8JMmCWBJimwsppCFByI3l+kDpegBgsCZY2muCp
8Da0b9FZWJlQw4NEvESt2ViK3+Y/py9ZrR2UPGhOxHb7W4ZuPi0UitYf1waqOBx+VnCGx68KjSFp
jQnvBQmjkhvUz58G1Oa/xfVlpqIV0781tcRbu82VhvMKqJ2FA9QY1BmY8Mn4ur3/k6YaQhTswS62
b/N8tt5KU6jZucHSNFKfe0Vxpzb0Frg5bwHRqExtVTwUnAXuz/DYKp5/bWYr0jRS3z0aLK5T8aUX
7NoWpaJHcwYummS0GJpOrTXTq7RiSS5j1RW91PgRravs52s+8XKl3q1jmKqN46t6a589afH0r/8X
np+3/kMC46y7aOvKhOpQfe9PqcwcC8xvPpyCMsSqxf75FIqIzDWxEtVpTalEVAQdxwqUdrgYgV5d
4qpZg4ZuZO+fFHWgvoScf6NfRi/QW99jZZsNjxFST4Vm7J3mElcUCLiihilKWf2UaDGHKV02h6x8
S9KFOhLY0M1Cni2f7EkRsRD8kf0gcefk1MLw/Fq9dtZ6XM+70RVyspz/sWCHf3f8SBk2WoDZJMhj
rcWynyuHYUVa+QzKAvee9Bsb9edfH0Quec55R+IlYg6z4EQG+NgpoWkqhtbjReNGMG+QNPBpv6Ji
LJ8vZaqcyrkKIMk22f8Ti+qzsgSNj5oM7idD2SRu4JRVIdudpqIWh/bivCtuKgBeD5xumuwaf9p9
YyGnkoQu8Y2rK9muZS+mdFG0uFmiaMo5QsB7bUA8l3NoqIAzYR2azFlJrZLicJH4b5E4KFN7Pc2D
GZte6ODb8See40/Zfip/fE9upSghHj6rZEQZXVOjDz7oqaP4j+jPtBhHaZPgtxoiIL6CBogGTYyU
46A2VmlRrUiIPrr3MQCy/I2E+N26Ut+in/LRoNhVExA+q/qH9dpyv0XWq8iTebpAZtaPNqw+CEmL
SPrDv1xDcmYsh7nFuhoYluFzrXicXCvFH01khmFakv4DANm+R8MrYfBkJdFAu+NsWcWX3KDLriM7
Pr7ocVtmjOebxR02ypkER9usWxai8bIBDQ9zmCBK9L/iMNxVVYMx5hii3QD40tVWlKLMABSVCJPi
61KTT1JT8geAn9hbtkif58FvU/0+3nweY48IZ4iyrrgXYnFSO1FBCQi6hOIFFQp7wlVC7cJml4E7
Jrpbf06clrEygHzzZp67jKsLRJkExhb20Cf70HKT/RSpO1KN8uA7iPSaRDX+pmScfwUaXIN1snWq
rCEzLfyhFzC0sFcafx0/Wwp7yKKQXdxetIT8bUc8eeYtdspr9kHy1YhetZ308cVLKjh7SEZnt5Kq
AsyAKmkihQBcM8npuGA9L1fWQwEAYSqBJK9FZ0jZCXaJKBBLrTrBcqJbXKm7RnMMT/8GEFIzZw1c
ckYQ1h7GaekQ7B0iz11RUSvNQFmZ+FrBMdW2SCAc/970rhn27rGFREj9ntV3cxf4SThrKmdtXqzD
Ks+qmoNkXklUe4A5EEJ8YfhEFG4gKfrjiFnoryblEEzcvzPwpPp81ICuCqRHTIsaeTP1rsAAcFHx
wWauLgzp5+N0K2RTCOjk1DJ5iaBtcInLcjt7iv9mx1KB3AZg2RsJX4CbqTHsNR4842pLGmYDOtD0
nRSJpwnjv971qaSFSa+gHoNkbVZiJmHsrRnd/5waS66QejzSb/bm6wc5swTLbMZX65E2Iw4fkuEa
m75+UZ3O+KY7EHDNIBwWpSqow4vVThQtG+OlXS83Y2bkIe24cuKwTOXCRrwzvDFWHRWo/FvyXuKR
rwylIEo11HrOUR01dL6yTFVbf7dLRa49TtrETeWameP6Mx8nnWdCPuxw/+ZWOikSBnCC5s0g23cu
j0pNaufRnKBN3nZLqjD0BUNUfLsE6LOw9ixPm+dIBlni6cZOaqE08H9kYFBQaxBx3oj7QGYc3iOz
JuZkFJRoRAawN9Itom5jznO2Eg9eYbq5H+hQMlRJP/XSdzxhZZEV+BEGQ/SCgtRNYyqcss1+VVWN
r29VBF7RVHG4tCV5odZO4JJPXW+hygoL6tG0kL+PeSqUN+sDPokCk9kHj8gF3El8nS6/s8VJc1tb
aqXLpkk4hr0IdmUjlV2caKt5ZEQIet2H9TnM7KYhHfrq/0wraU6TU/cleAqFpht0UvS7ZDuUMUym
oW5FmapYR8qoiBEXrcOkI8hNSgZG74edGTTm1P43hWtVD55WsFJHCbc2uJwI3gD5gbHAXv64ckBI
ZYG7lW9YyXTgpkDBKf1zK2il0bF1M2xYjxEXmmQpE9MZdrysLDxZQOLyuEvkw8MwBGFikcZ3gt1z
IMGlUDfK97MVP9LpNRRb6h48FLyZsJ3PebzURrRvKGuuRFZ+USlt66tYtkabTzyXM/7sOVlAkRSF
l2aS3aMM3B27fW9GzjT7/2FnUn/RSh5Vb7O4FBM/fIvNifF102SttL0Q20TFvhk0cz3foF1l0kSO
6nt9O+wbu3bbazexwHijAbex8z+4fkAvSkkuLaqk8Ln7Yn8rNrYGPuR7rRDHYyA5DuHI7BmvDB+D
XtuaM711H5KnnBLV1YVO8+Zm5kXzZuFPqbMXCFrsnbo8ah76lG/GdllHQ8Xb4jG9mniu0GaEYlR5
yCwk3PFXpYG2DOfDzcVbxnvVFCWVwgRNg9K6RCuWrlXpe4Vxa+KsQ8aJAL67I9Fr4Tqdsk5+hNDm
UHuKl8MHEBd9VQjdyOPitKvw7l75z84VLby0ueEEVe2bn3puTvuH98RGQ7C8jnwgcWKU/6VYx2GE
8MdCCh9QMwEu/Q3hspM8exHFfUZdfqyXnORcJ4aQS+QckA4QvN+K/W4wRRNzqmOJmm4C0K43ucfF
fdJy1JgQEwS26dvpgz3p5dPRJyvnBMRlYWri2DkJRgDfZhKWlyH3bno7GkiqPxPaXdxL4EOxPLIl
s3roHaJR8ZaTXS+DGDq0KkBqf1In/VTu4SxZNnH4s5DCc8n5lzVQ7hvzhSiuoEY8DlX57U5z9fJk
QC3LH7FftVcJzul13eWY6iORr729pbZJd7cbpbFgOr5cKToCX1RT6v3ZA04du3O5peKBGF++OHTR
EJeCteJtQ9RJd3aOIo7A6SKzaOkCRu2Lh7IGMNUDQ/OCUAI9NxXMjf3bCAHqlOjJK+N90bKk52wU
tFEzzK6OsnyN7RuFrv9LxwIEkC18UA3Nfk+15TtOkgLUDRL2hI7lzTGDU09wbO2GfCGwVJju4oRi
ZSDt0ELLNhMAWwg7f2ilnH+sgRl0PREPNy4vmqjA7HNK3uW97dCzIqv4nKKmmhCQ1xUQn1pXAd6f
srQn9kZw9P8jmBLvbgLN5z582HqJ0Iez7bfi4EHmC0nzvbMPTAh7kI2qA/EOj99tKwWOZJBTG34Y
zjT06z/X0GFIEx5lQEKZwA5/EpRwezhpA8e16hSMQbBZ77wfowYG6d6WB+G4y/HcBGw/CB5Esppi
+xK/kMhbfxtB9dy8Xe6kkqhVuILkcF0Em2Xo9aftWEoLjd2SRTpu6E6wDjDby6xvWBqGRieOYImj
J5+sSAHSavTrq566WbKhjZfITzZGvK7kshlYbF+9tVjsL42lyPqN9PGD+0toWLR67WxUDc7Jjr4Y
K41Wm7Bo8NSyIYP2qBlyzYsBQSQHBDrcx7u8x/bx/NxA1yO+6dTj9vXpz1YcrIKQy0n+AnXo8WZg
DUk89fqzCbgIs8hPTuzW4l8oGh9rlB2MNSnG/mtpj7xf5sdzragKUTEU2vViJ5LstiDcUFYWgncg
1Yj9cqTHvj8nYn/4sHfSB9DGW9Q+2Ki4Q5oeVaWMVnGPC3egiyLgyrLKFrjrS/GmwrPW4SJkDjfa
HOwOkTX7L1jrTfNaQSKly02ciEtl1br034UcbxTdschKYxp3kQvrtAFXJpA7CQ039ZA0lrYc5wGW
nqA39pTJ7ODqEV0SCgGUdRPpeTrxiZe/cuG1xriAsliVAAvCgAu+9wmnyW3PYXmLjEEaOKvnhEjC
XB8yxYSY1LmmO2e0wLiv0ap04eN6YMPsl0wcZW7EBiB1o5Oq62y/052a0c4kNHRE4XCMRIxqyaUg
+drNAFkJ5xCEciE9QvSqdWr7JQg4ExkuW7UuYQq5gEXwY2d3UiZquyoGs54H41QHZfkzJiMi486U
LSnuNdkkvyUsTdI3fprnTTHab9vSqiw3/7N4UoZ5lKJPnx+XJtuwCGi49e7pwkS2RHm/84VipcVO
vynEydlwNe+c1pbrUIUM5K79M6C+LVc0WgZ0Kz+3IH2jZrFKz/VY2kciJZDgvBapTkkZuSYqKHlH
xUv1vrI5PYAeyZ3og/6YPGFufcPcsuMh5wHf5uIA3dLJWfR8Xvwe79/6uUtNUcRLXkaZbHLD59HR
4kP/HDK6HqpXYFI5e9NXNRmns/x5shtm3PyK/BHVg8iiq/mi1VqM1WwJOgyEUYAv4L1Le4RJqRwL
34h05DFZWDgyD/6PwkHlhbCafXoHAPXS8EyKITcz9yrBOM8B7JTEsd5SpOsqzn9YsEfEkO0kk7zG
wPfSPuU1PYrlO1Kab5KttYDkWszkSGyD5okdi0WKrTN/yDeJQcQ/3zjblU3Tsq0F69MLx4arg7eM
6SSYOsbybtvXZLnNjJme6lrzoeSTGDRYe5VfSklUaXAkV8gf/etbe9o7s/b1ag4Bi1fWqJyQp9we
BrDS3ccpN1/JgjVa1o8Mo1INx2KL4uwWgLEQVks+glWvAj242FkUQkYhRTBQ/Cm8HQM6Wb9JGsXz
hpXx1MtTA4FoJzewkTRatIuu10Wmhxv6GVVfDKR26Mi1DA561dGXI26L5k+WvVxZlFpr+8Z4ClVg
9Q/87bapY9zUJ0tsvZzcbLuMAbMWNJCx5V3YyDMXNAUdPnBqXK5c5oJuJSh0u/3yHDD/MJ6F+uAz
lcyt0zSyYBLsWCI6JK7srND66DprDfcC20dwAYdUq3DfrFE5wDj94H2Dq5TOfWoIh2gs+a0oRdnC
tOfvvPiMr3GYE8EDS1sB5khIeFkXTC9mdNURe+T4tpJG28VD4PqYg9zQNfZAx61P3DbZM2qkCM9B
Ee+9ZBKhTHZbzAQyHVnm9v4MwJj9IYKz2eryq7GUSi+qRp6sSjOiL2BkeFizqUnYseQfEfnt/LhQ
qLw7jt90oSzxoNxZ52KRadXZczp30IbvTBlvCb/ML4DUASClxo3R3sq/amEpCa/5w4F48FTSE85r
wYnBqTsf/jnFm3KPtNvN76qGFw6j7i4PhOHd0fZvzR8zCFXbEm6Ms0q3iN6dbD9aGYwlZs6qlEIy
ij2IJVAvMuiGLI46Np78fqCiy3uIC7NBaH8Nu1t7hHgIT/xF3T4msUWvoZwSsPYYO1WMFxhoJv65
8pvF+klSGEQFTTqeA3/vI7psuOgNPKvMzm2VYwbo400m7aJyAB5t5f9KAq0ds+ZGNTQbwlPfWpl6
dS/v35ilMMBPEfoLNIezdDlCfLMdAbaDJxnvclyx1LFWsFjVMC7nsixh7mW/a47cZPkQSsd0gbjQ
jS5ay4+wiPVQRIGAVQQujRQpjL84uGI6uuMwK+cr1lsl2pC+4GDNTkIW0W6Tg28sfOEgUr8C9nCn
lWNdDwoVcbtjiqsyGmxnOnoBWQ5nX2Z/5FGhpCD1WQnyLul5iQfoE+bm91JuQZhC1VrmF5YSfxVQ
aQ6LPmmOraLnJzj0Wd2TxbOIkm73fQOBN2XLzkGiBQiM5L+IWw5JvqLD/vzBM26nHz7pjJprE//c
GFy6MbKqXwJWqrUWbe1QPOrrjRxPIsK6mfIaEPDGyoleNP8D+9rWdC6/JR3tIAw1qklQRmwBNmxU
c0L3g3t0x02TnjdibvZQJbBZK6YIPECQ9JVdCHK1zxrZic1kKPFQ/hvrQcaeJy6Vb31B4XHN7zis
H1OFkl8wiCA6SfILSABWLW2QitdLUtoJ+kFbyeS5FCNaxmdFkdxx9uV0y0cTs1L2+jXJM/myQCTA
Zg7rVEeI+xZ/OQr0yeUX3ukR9OdqLQl3Dn/swB62Y/EpXFAEUgdLZs2lxsLxZghnDKPulw+TT0qk
IrbtNxZu9tWM8vINOfEC37thhzFGzeG+UVnAfa7FCX8fa9OVtpVNYwkBrxG1VXxPXs4b1jT0M3Q0
wR4QlLHkm1GWOQi6I/YK1x7aW7IoMwsodJcS7am8y6/cILA5YwGHz12kgLVQPcFRE0l0ACvHIWev
WWYtuTiz+WQJuwC/7USZ/iIg25AGh0S1oKqN5OKcE2Ipfpj0BdYtiEOwNW5Gw2Un7MY7pTkAwaTu
Ty77nxjTE3KavXlZ8gfIAuEog08IiRdBf7/1HqQfx5dIKCDNdCD3sT3skJk1v/o4Xmlig+Nu/f40
+TpSG43LfjcSMxs+O55t82BKVwT94H7p0KSAdT8TSIJCOEOgj9EXgvqqmI6tKpWjFCYHSiQFcob9
UGQERXDOXDPfIJDTlIK2xPzHMhs4+AwkL/7PryfH9iW+CGhi3ZAexXBOBMTBi7iN0hQw7PfuWynh
8UggBqtjat/KNEfW4pwO+g8JCLIoaMmop5QcGkVrAzjIgetkJZQfD0qIOT4G4IJTL6AapLx6OYnn
ymz6vjwyuoWmJTpu1H9b9hnyNuu4xNmAYgw59h3uaFHf/qB96uf8rMkHariA7xbBRQQnOAgXqX6K
OieLcOxQi1D1KgFSDAGXo+B3QxskmpQr1D/9AhJhCLIInBWHMLeEY4aLXci04jGPzZuADqdQE38i
pQ8DgYtmmTVJwzLYuYb+tLrNZP/6uo73MhxKXCmJ11eaFJAhwxQSc2Q/NW+PN/n1Pa+VAc9cFDD5
mhB6d9cF8M7U2RYHs2/BoJz9bHoX/Riv8HVpEW/tHg7r8zQR9KAwTHMge0rm4b97v3nhNjl/qTI6
sxSHP7OSZgBq4Eth9RloVJ9iUNcpYV+0u1kmx+w8NcG0OBgPRGbHXJYMY4/BEEMnYThj0wP6H/8s
ybZkqfTklJ1sWNC1QUQBztcw7DLj09S49lxvKjLjTgj+WYoOhVLgS/vjTKy3o8z8LDwnDdrAOzfW
w/WdvqEpGjZYNdM2RKCAhInZfGN37IrsTN0pxcEtQbYj6ucEogt3KDIdLgGxP8OVXq6oukNFKwxT
/S0WkJRDFRNO80Xn5GwAcIMrAa1K/r+O/1zJhfP4RAvHsAsfBm41FOoRmfMrcikMt3X3iDXdMgic
z/bAwYTPLXSJTN0aYEGuQy4h75wtAKaGV+Gzk1MRsntc1l+/RqewNfekryfiQ94twPzT8B7RPXgx
YkO9JZRHW/OW/EB68N+3ivp8Wv35S8/P2qL4Img24/wAZc3iIX9CicofK+UE3sEdPvrKhs+nnloH
9yk4R3Qc1jZ2jA64/dcNcsOXBc1VN+n9Ch7+WwRdbx6vIsXWULco9ipBbb/HNu97Gbaox+HVQqrk
twtwQ45tsMjko124IsLF0K3F4KybZZOS3Jjv2DFdLpFOK//U5dTpU6oTo72uvzSkmlxvWvgoBezy
vKeEUuRlIyk7wrTn8DBYDS+PyPJ0pl8A2lYW55nyOc5y9HbJgIclLc0AmC4PZ3apQRdK8N3G4D7K
CB0OOfoJxJasH0fbJEUmnHTTfkLS+QP4XaqZzeo3AcIk/dRfOxf2Ly6FAyDbJn9gciXYx4WIso4l
PvuOkApM3cD5upDXVtYh3qrbOcPq2/QT7ExAzq4qklhaK0Cww34Wtpb2KeGQeVj2rj5MW6ybcPZO
z4rd6Fgne/gMu6mAcwuc2bd8K1NDZyvOPsBnnLbSMH3cVtkmf9ahXpQ3neOUr6yz9b3RoPXQnnoa
MOYRUDAX1wIZVXZBZ9Bkzub5agKyNHFX7H8zghiAGTWDxXKEfd2j+crcRlIrYPThJ0oP6YzkR7vs
d7GHrSiGqNwKlMMPcMirxX4ydUZSmPhKNJw0GX3tEI/hClz+Z8x3waYLbbzYnfxS2IKi1T1UIw5f
Bxz738qEp1NPDc/JmnQofDAELMKMNSaVlvj28M44H7Muaj3TKF0fe/hk9ozEC/dw0C39qHBvoWyl
uW7iu/XM49qKUG13HDcY55BQp05+4HLPuK2P8Jc2qTxDLZXZPngJtdSuI4K5skxp90ESZbGGLCpj
yeYSz6Gt5l76/vO9/l8LndVHln6OvVLnrIkyjAXUibHv5cbm2dGt7zrbOPZskafnxm4seOq+wqwI
ytO8+fYbDQhCGdeinx120QvqZ+PbXfVyJB9ly8BfL1Eu4Qy6IIiOuwPjqMyXK0kfrHpkcUFryqNo
TIDDgV1Q3SCl3ken+OzuVID2hmV9Dy+4d0QRaqsITSeVbLF3yeFz38PuTOX+FI0aAGds/A9Nhzo6
WLrEjigaO5031LOY++kLdEnAkBjnmDAO8SkrXzLB0rwnXbH7VBjPdn7ZeBYxF+souOpI03BzuH5r
sv6FhWTureVJkIk6GKtYoWAARp2M86krI3EMzqeY1YXq5dU1/EPj+j9eaiUik3OGJgfKwiYRlgzu
qyFLYULV/qwv9YVCe6BE2jC6iZbayabTqa7zR1IQHIbGe+dhXAoWXes+7F0+X1p9UNdk7kDbbpIn
Yxq74vDJU0JBsN8onnfz2pNqBRMAScRHwxJP5zLaxE/38aB/SYnzmQWdvZmnqLU3TD3Lsvnq6FOa
PgTu7Gjj9t3baud0fwicTvfFwENx+VdwKoAoQ5mwd2Zv41hc+/JX/VPbJSXOTwsuongbeRBRSQ2q
mqUPuv5GvX0SEKb1VLkrx6cvwygz0xvigRm41y+BI+x5cqXa0H+hiu6keqPC21KakY7V0H3Vgxok
375m1/N6QRtCzXwpzDnsgoyp+YFF2StFBG8h4Y4BvQIqAKHurCbnMXIVHtzh3MVimRztz888HIbf
9+6lHA7oIQRAdMAuxa9bRpCRg+NBpWygI79gd+xvu/ynsa8nWmI3cHmRzCIbv3TsmAf2i4XbsyZs
C107sbm0J23QrCHJTF92XOBo0i/hAXWCJM+a1/jm0lfvFn1XWr49iBqXHozVdxtzJHFDMfuBTago
6Jx1mdN9RRTq0LDXqgK+WPXb1pEDbdSRXEvuaTEmmeYVrxLCcxJFPQrRZSOdIx4OFgWSBwasGkAN
Q195UC/splg/z9/xrOtBdQ+K2eJ6AWl2WWotQIPeBJTxzhl/TbfhkhrGGr78cppk0QCTEwviM45/
mvG4A3qiduhWUzm301dNUShgNjGGTXYWNm5i3oxLbixAr5h+1R+PA5KGAC/B/AVnnj00g2Be4tRl
5hdGvR0vRl+HDUWCam9uTg9H2oWw5/57NlRxL3TEAUa11KcLDFWdy5H5cEUAVfts233IcUliZe6Q
fckggqzXlrQIdozSOlUVAu5hg546LBVVeb96igV9+AwX1MYR/V4jkjk9UKFKNAX4jvlsk5dxl2Sa
UdsDyr9O0ld/DYBxTBYM3KoGqipaTPFDc8ea09aKKop2hhMdwTANyVBqyCeOY7j3M+gijTtsYD+8
fDPIKc1RCEnWbGHn5PDr/q2thpQ2PkjFDW6KC78n/DMPz0S2J0nI/rx8l+/GF8eia4MGV4MBqKaf
IMxiofhicPKfGepFT0Bi63Vzz2pzOkNPVfMoQpK2SH7Ic5y8eVibk6K2XOMGlcZZMsK91N60eo/n
as30oVnDYJbTWoVFwxgD2vmEi7OqiQW0FqsT/jn6WspZbcyb3+AFE6Ozm1WxVvjDNo6XBtIhVzpS
n3m6xourBr+scOFrfLe0+lE1dR3AOgEGMRY5sdHjF/JP4ykrkxeszSmM/9hIIfieMhptIeCfbvMP
Ol9Kny71CoxjNRVxSAnw/oZJjNc0Z19H18lloohICL58m2heLMI2cB/LSAlCbFCwjbtU2sswcDru
Bn7rAK/yA8S8oUuLTES1GlUDHnjCs1HQIgE7esw6av5iQf4qK3iN+lP6gA4P9HGIL6pxG2Zqxskj
r8NROQYydDiyKZ5lt8zJ/taUWpQmQzl70QIc3X7Qs3Qc/CTKwKIuSAWB6Xhgxsy5fVJz0v8SpEPM
eVft+Wp5HGEOJJbGV4E6t8mE/U3XXOBz1qR8FcLQ1OxWps67LWxvp56IUhTUt/auq3gIqVzQ8z4L
n0gZpa1oFyvRcpvZPGpXy6gr4gdj2hMcfdDU0fdJUfIhg2ZuVcrn5FJ6LPiKvVK8/d8z6cUuD65s
voq5ZGGloTm/BuirFi6LS9RdbZpz/AI4aRZzRAll0F8qMopwQDYLpbzJpsmeE6hhMZgyaWEcb+AR
dlOka9JuWVYunZ7x31raI+/E8SsoD+O/MV9bWq/OThny5oeUH4ykkLKkrb215bWp9u8FN9npLGrl
jPtOG26B4V1cVAJiGlKkiuL2wQyQvBDmR/BwwEYTT2P3BvIYeMK7Ad0uXQNaJs8hL5i4Gf+wYTdc
NbRF9V6KrhV9lOH37SkYXBmWWebQxI8hRLcY1AWGBJQzZmfHzMMSQ74NSbEfA0/g/clgHdW0Woz+
HHGXbEvHnaNv16kp7iOnw/KAmM6TGvFHYp0KyDnIQudNDbbdCw2ljKVloPJPt3J4vaepNwVkXL5x
K7DilsthCGmCNNtGm4o3Lq/OUsIAoYRz8Ek5La/uHHEaVaiFb+IkrHbSMNwW/KWXli/T2aEmbXfs
IyndgL9d7tnl0yDa0bJ7guTn4oYpP7iiNps72VnerHPji/ECD3iVJUDCNuSFQoOouXhyKznV8wjk
XIStH30rBg+2gUO2Cw2EtUrSC5u93bg8KT0DiGSotO6lmLtdo/M/HVHFYzgk57XyktDBS3bJSqFP
5I+IhcsoSkhUXRH/N1wmCkBCNk/qqqvrrlAxBFdOJAyQP0Ijcd3sdyoIGHilxs5JQ8i0NHNHz718
3d4OQg6c3cGFvdG7xmBlsmDBtIAe9I3KnusbjQxzxolUkWGZKpDgdH8qJPliLCB8ecG+9WP/B2SR
Q7VrAG03YK1FAM+KwpUU2T4KW9osMx+0bzUiQ7Qo5aavDasVMObXhL3JKMrR7rsaHzu/0zqyiXh/
QwWXPwtikf4098qaWQCrI0vv0XMwZ4miTwi6KianHljWca7Y6wtUAbqhdTsyaY3reYZgZ6N8lVB2
Q6dRTl7CGxWt4VJ3JunoPEuPjZIW6urNwnxtBCPiUh02c7u4SozE5TMPvvo8PyeM+r12CqAVVziw
mDq5mmtZI4x+gmLZ5Dtk8vEe26TVGOH+b9AdbnSYi6LaAWnOog8ckhFkLtWuR+FkPrR0W2ETSbeY
wyKIejNY+12Se3bhLDo1j8TaUWTtiwbTdaMKYwGrqwdrQI04Y7NfN5jgc8csr5KKvF5XH+tcwZTC
xRxxl1mgSlWQChnezuR3Zs9P+892Ml+hk9JWS+WoSg8WvjwdIwz7UrBOfLtKey44dwhErVMhrG/e
+G3Od0Q8G+LyrVUc97h9ePJwsyfWi7QOXlGQ/6R7Bb2sWOhmgAVnvKponLE4PrG3OPxmF5zs+gaX
EPWxa5z4uDdjwRK3PwHSMty77SXJH/hEJwyZjuC04BNc+rKHhHGLDqp9tdCWhv30K7oJ3hhXIbru
euhrFDEDOQJKCMOtJjrvZPOVdgkXf3F7iJtWG2PzXfBMr0ScqGmCqSpOOmyP9bUSxv0V3jKLozpg
zVm8dhv+qryjiqZ6oYi9fmtcF4RdBM5QS5NQEmRBdkvvH4mrJS1g5j5UifrrpW1FWs+Kk0uleSlS
GG/AUy9Z6X1pd/sC4MUqtJjxUze+bzM9l0WB1LkqiIE/5GEBv9wBeLQDqApKIfqGDhcHhYf9V0W/
1O3cHHinVnrwgGq3nseyG0vm3inEvo8Yj8jK7lLXJdJNwH1hNbM3/j8b1peBQW237c2LN7bUggAu
qInlef49KYQCVRf6SkO+QA/t10bGd8SB4CP/m2s1ZuBQciDAwrlusaLPu1n9fq/TGlppZvUBw2LQ
KsKuENaVNAhcT5+w/a8tPrBIj5RDAmG4dZowbQQqRRcmNB7obQRLGMTPcMCBNONeVbrzGrApVbHJ
lTE4/lnG/tyu1LhS5AEL/wT7gg7ZL52E+Vhsgu6/vYMQ19npFFsBRC5sXvif5mFsv2cWdSNBjwyB
FDrDHFUfb5c0rYwp609iarb9sOkcRsvQ5ClIk/UnY7oX1xmWs7x26cmPFf4bRtLMIvgqCKSuwQks
zB81sdEFkECzKUclsah5U9zn19JqR5IO2QhWoqs+7uhq+oAW6tvgKZcG2AwJkZ3sXUoIdcv65auy
TV5O64Eq29XWu4Q20D0R4ezSnoL1JoMphhxlb5NzuQ+Mw5JYabeI1NvKQELzfaHx2yOj3UyNLVKj
ZU+oDNrOb1csWPDzM12Q0Qkr9uqAWb9RmL3eHVv9+dqRky7JNAxPZUnM0ZcYoxiHD81mQ3FS37vi
kfeGAJ7+husZYlQNZVyMhrly4hpLVVtHoM7ZJ+wh+N0Sf71by/7bxnGHI9d/xJaWICPao0Vl9/OV
AcbHqgAafLlOoZpQC7hEMDpsD8tnD6EZ0ourV/6rwu0NPTU4MzBtj/uRhJdYlWjHDFt5R/m/my2R
uqS/rBHsmEujUgJycnrVF4n0LholrEs2bSrtVH4T766fdCkGiYsr6hl/2yOwyQUIIPqTW7JuuIbz
ZaaocXpUpU7TmaG7Ft22hGZ1SX+ziGG5+d4njOJU75dtGdTL/55LL8isvCQdc5RwhbGQJlaPlNHQ
9U3H7tJRC8Enzllxn1F+f5YStXjES5fbB2ArdDF0BOW7gLh+fiF1rAR5tK7wixq0LyKeUcPJiQRR
6AD+9hySkakl19vBji7QWj0vakUrxz7Fe/NvuxWqhVulHOCJpiP4OlZbQqnNWNX7Nh8creEIwXMJ
OuZ4tyc8/YmspoGB2JI9PEVe0yYUQVN6Tk/qhDTD0tZD3scK7GFaMMp73wuKj5z4R7OEjVJIHD5L
Mq+uLuJA6o+o51T9C2T5UfrcBbI5Oar1NWLlReJSm7JvnEqD+UJZ+xmLnGSRWxLbzfyGw8Dqx4PS
vvnogzQ4a5r+GOE+ujmH1N2LTxfTbAMobvemezJyxSmUN/aAKFXN+NbTj6N8aAGdAk9/8dYpJBlI
MDg39lS0FHOIUJU4f7nDojqKa0b7bHvbz+YZxlFSoCNNt8GUYZB5lsV80z2iND8hMY99qu6bzsJI
iSgNL+I53xDokog+/Uqr66PlFPbV5RIycdFHjMSn9Ek6GEfxx9XZXLnalU8h6v/mkl3BETNXb0Le
4VhVAnOQLYQ5QifddfXY6izIkDcjBSkKd5l8QASrKrBjZFqtOM01PMb9vKS7GVpv0ILlsFjYtMBM
noYXXD9T3IRSw/eVlgojYX6AZJEo14AJehnFLrqHH+5TQcQQe3iSJXeGejPv2gPsq0cDZoPpD0Qq
3vbwMI0xpq2Dij/2ZiUwFJDu8valQm/7iyLEjaqkD1NTwHHe3XubJgYRHtVHQeAyGf9k29OVFXmB
9mxtzfxMy8zWjbKUTZQAr7B4L7L94nxV6aeGfqyB9THlrKTHcZUXNFlxZHc9GMIhgd42Oev+Ev8x
gK74md32tBZgZQ5/SzpN6j+yU/TS8Ecv0C0QqvFUG8EOm1EOp6HXtFPsLlFMR/YLwuDAx+gOe7r7
tyotFnrGwjCAOgq3d6/GDaTNaNANGMCKVyUrItvspH8rWlhkFrcb/K4jR5OlvG8b1U/Jgw2DBQez
XSJZZJIBW4wOUBKbXRgrLC8E6j9zBCF8aZ0jy7hWlF8IqlKWtw8ymgkYjFtYhe9mWIkd5zZc7xsg
ylByGS5fKItGbWVDVLirUmelG45GYHuQIac9nICG0LOsKZsamc2cX/r0ARuYYfFDZqIZB9KzpQg7
8HRXEHetGzuYULbX1wIBVr1R7ZCGYJ+tAk5Yib2epNjlGJtOSX7pcBR9GSAjlhtZ+YaJ8hALkO1K
+g5Kj886RHVdQMez3kWUjpkfqcjf9YiNQcVB35yc3uzQGfQqNOHolAl3yYp68h2004lKugDE/ZU0
/2p2a7gXGAx1Rg9qpOiI6vZZ1lJHox6gjq55hNZtzrAVqoQ2oee0azkEma6bKiEdx78YmPdAAWdR
JkgLPMcVA9O1KqyNcpZ1T1Ck6RfNaC+AZ1FIgD48d5YSRKHqPiNFi6z1Hi7CdPgepDl9AjUK2YCy
xZfFPFTt+RPuOSzPbBkAvMhvbJrgr9Qg/QIJdbTjB22Gwf5cy4o61zXak/lNNYO0v4hUcKFnXn+4
ewuu4g/NUGbnW4v0B+Ny4VTRnkaLHmPVv5AWY96PCQ6mZxmjftW2fmcoapqJRm0iseBda7PVfOLL
+rnv0/eh2pLH+Zu9HEEwwItbU5K7ZWlDWf3Y24z5eywzhz6uH1O3ZrlBK+qW8T+i/xS3uIZEmDiz
2NQIwdsOCFOeR9gnA/jwzXCRKKx/9MLvp/hJyKGrk8aQ1RvL13DL3tVqJEtwl11bhBfg23SG9o+T
ajlb4Ho7sBoQ0LYGVsGJv8qtW6gllPaeD6Le+kKtshGiDRv8vBD6HYfwQ7lOLg085lHi1znlXfRS
34MTH6bO+0uv+JX/i1T5ZICEvqA1NXOF0Fd4wAIQzGC6mkh+ooB+1nH6GXt3vmP4RcKWIYfbnipf
LPSXP+dRLEiuQ0EBQ1OO17MXn5x0tN+Eoyta76UwDwlBpmSksCDQiuniLRgLOuCxF1kEThwidx/P
5kpTdyTA0wkJW+NUXDtetuvUHPZBqYe389sX51MydfW0EYytO7QBr2tm0x552RtE4sjPF4lCbhu4
AX3vkUSpDQpdopzHHS2Pu3S/rtsrNed9BWFggYRL6mFpTI8l7NhoPWFghyNQKQLhs4noIkHbhlIm
/5OnDjYhcuqdrZ3UxLx5kAYzOxu+jps+eSTfMtMQtKuxyf9NN5mu3NzP3NOzkRGWnpNk7BPRhtYl
cJxF2hKthxTrXD7OdCBgPDuk6NDVZmxqcYER+EzJW3zhgc6FyWRV3wCIg0KSpj4EGehosFe8iVJb
CeZW+FLSnJuML2lrMPbalKLWS717PNyG4xFSCevUxYM9eL4PUOZJWG/F1NQTdDSC/skjjXBStkCH
EiPdnr5/QOhQlV8CiEQlNvhLzr71Z0JLAEVx+E6BRvd5ehkU3m70SmckS9FjBk1wPW/IPAZO4/an
zXOrhH98i/yYk7Q07ZgViaOlHwC0IAc9CvzIsjjxuCvbF9F63f6dgV0vKUMMD7Qsh6ARAw1f4l3D
K1yU4Z/maLtJOpQOWbRlBgjoqVD1WN+/qAqd70+kVf9IVPBxUl1RFyoMl/zKWBEqR5JFO1ETjGxg
e80nWu5mD0efR8Ex1we8s3Np6DujLccpYQKW/xcFgzVTOKoPlXyPAN9d0wqXReU8wKZNj6/2Fg0a
jVtb9yye5UqE+E1at3sTo/kIjcmuQDBS6jG8i8Musd7u08wSxKwWySwlC1ZEcP9orgXIfHwFqANG
QjqHF8+xBFUDEwOQH5N0PdH21Aq3Sdbd9s3Y65kkAdnYYDef1e92hPR7ax7C8N3AGjLyMU7dikBe
DT5Cb0qyVdKAmDxWEAY255jqOIGu0lOj2wZy1xx3z9noggc+8NJNIOjqzWletefQ50GJ3da4OjLO
vBxm+Q7qB+tkJW7o/ZvHKzbc9ekgtBujBv/diMRgNcT2LrqGOH7mBPotHdMA07FYuiTzpRnCKrx3
6ccIOzZqWrxsWe9Srsu9z7pFX5aOA4384Y+13WG/7yay34Dzl759O/0uJdgbUnIh2p5YH13JVDFI
+qoYE8ygsczKYF3Y3Tcllt1T3E3gRHJVEyvaz9zhZNRGW0WYCYvqcTIy4v0LcA+oi2mD0sTpsMoF
B49WD77w0YYO/mIK38tUe7Ln/DTZiFcCEsmTRTBtL1EbXwtlHFkL/6I2cNejqdejAs8jPLqqk8pI
N5okKi/MOMX8/Nz6973yFG1zQ3mVqD3rpE+LBD5OoZuVQ49x53uY1oTCkN4+h/foputapmfv2cR6
yL/GdiwR5PIa8d0gydgIQGNtc/mEVQbamUDuVFyKJK/l0RcttI2ruTMAEoc/f+ujc/7AvwMMgxTR
apYd3soMv5yQTuVfTonwEdq6iN9kbkMV9DPMHTPL4k0BL0psy3gtRoBZ01DtDW3edzXcdfzAbBGk
1uzTSFCxEBWfK227Yi0MMMEVF6aQ2hOMuNuh5N6Ktp4PGPTxhPLcSbZpdUkF4LWCm+/C1dzXQeTr
OfH3CLWCrlv/q5xbAvbtHuNjEnTeVZcnASNEsTtLZOlyjihakiC6F6Nb53j+DTlbuM5Zfh1wwYBD
38nc68TOINzuG0XjbeBlIz/QufS0IINEzS771nsu05kUDX6uD5nMpGe6EnBGzDNMotnXbdfX7n6R
w6yTauiQxFSHduFAUAhnyRGuLLq1X3ZHswDIjpSTLa+sfgcQIfwxIN0C7ml6Htjg86UzBrhAHSSS
MUPwnv6XjQ6KyD+PWpL6y0DCQIFIJghBFodpzjO68sOyMCXejoOZChZWN6N3V3N8Zz2OLSzPHD6u
zMAzqt0jar4XWowle1kI9pMpJbFz6xSLj8XxXtz+kyXz7cYOMiE2o6jMPJ3HmtPhbVNB+gupDb+a
dmejsYZd7kTdvF6+ZAnERTlmQ7/aJRhNuHI0YDl6zFD6jgOe9Gnk7Q5lwJRkxCbbADChyVy/ShrJ
L1dGD5tKxmHwVEOR1mlshi3Ekn49ezv2xksQhwznC7ccxm1WfVM5qKrbMkc2bCD9UT1KasOUOPIp
LkwyKvYld6E7hofNzNwVdebMb2YnPCEXOGOYIl9BVM5cg5kgQHII+5gk6m9553Ssqf3/rupzS2QQ
4dDB1F59eucJmPzwOiAvHt6IMZU7IF9UBTQ1ld9ITkdUR28hlbWzIPNC/ptXDApLr6ZeQr4UzEFU
DcGG5EwBhwMQHoOFN+dUjFwW2qUbbH/T6cZANNWCwpqn1BtD4DSh3ZyolP5ZloRNvFvI9RVMiyVY
mESycqDbnJ6WJpGo+PMREhW8JQe3vxIFdpmNerKURs+oyLr5qn7BfJFEgUYeS7vM4VHJHfrpvd3m
WmspyZf1EwDuLpKQ14NYPsGpNR7Ms0SDxuPDDI6GjrPP1GLEvAi45cbVizfaaUoE8NciivfOFuXK
qCT3oMtnET+FYlTGiYh/1SvGUQ53V3WSaisvvE4F5g4vR+jjv4A1jNT6wwVdTMUTy5f/VrMwmFfG
gKt8UQV1JARn0u0uM9t02nWZdwnP3PC80uckzEM7iseezTJAzTUkRdmGpkYaeoOCsbXEluWe1+rN
xZCHbfAtscSxOAYOjtRlIOXgQrYfjVuJtb6M7Aikvp0A23jgFiwJLdFmXLx0PJY+BR+OSJhHispX
+mZw8RDEzdhxBneBYYZ1hg1+U583ZbFjvBzZuMtmqmEJJfwSfGMiQ1WRVkYFiBnxw1M300ls03Pn
Qc6mu+Gfs18iZl7Mjv1nCUSQcbtcL2/PYFmHyvj6Dy0lzBBQnyUFkBBPjAunt3zCwsYapqvQnqPh
isU9ONaCiSdjRALNAuE08M1nyQ4hZDS4UpfneLuHDqdrdXIrw/3VEFTTqY9jaZPObQBEKYARMzsr
Majm+G0R+cRcZAoVEqx58wgqIiZZRDOxQ7kOo4CAOAAKl3rdA1SMdVkUOpy5D8rMFtl2Go75cYU+
IpqjaD4MviWmZdysxxiVA9pCvqvjkCB6of2jRX09zKfDpxyLThLgDsbbtgkf2BM8RjTN/cFFSY3N
kgOoj13tzw0UqJz8bulktbHYJ/McYBNxkVt8qebyTINKrPqpzvqnveI6QWiHrapgh8geY4EHqapI
nm1O1/haqlMYc645w5LmaX47IgwncdYR7lnMhy0UiyAJK9WojFOq6smQ9CdEbxZQ0pAVtKUk65ln
NAeF8St23pJ0YH2yOWSciJ8vTd8EZcjUY7C6W1w6MgTXCXHFRJ28SvkZwX5ZStyA55K66/jCvdzp
hOtCNWH7reRPSDzGQd1p8rskZaDn9kW3zr7mWIGelT7KUre4ZCGpxgOs4uweuo7h0Xhwctpfmoh1
eSgrGZR4lmx24S/IFHFNXOooRqbewMzuhwRT4ZC2DNDwQReGn8wcQMTmhlvpy+EYbSlHuR6dNIbr
y32DuQCATG02Ef7tMqp6wQVO1zLmkcvDLLPzlIfu1KwTGMurs2y8UeKXmWINWUbMqFEQhwFvSsZ5
k7l03JesYaFcpnnIoOJ/hrBgrxLet2URPJJpaQUTySt7ReIcAOX8VhRat7b1NMGbffglQxF83Rzt
FEHx6JWlwyCBLdReGb2MWBEyXZYTv4N+vFPqJXJ8eSlkUXa8apFVQznmO6/+J6ubT/Nov6VdbIBQ
xxpG0eYVH46jKU7JpaB/Vo6J6jsbwTqM+ll0+0jKjWaxHmpXbNUfjxXXB9Kbrq7KjMDShVHp/zSU
sAjShpX6QdHjTjvjfyouf6kBv0wRztbNtId8dUI+3HCUKOUR7SZ5lwlEsKh8bVJzoc8gPNIv4jyR
RZk+xs+ZZPOkpkJJQhloecl8ow49Kf77HdX/EDnsocUNPpYC624vYYURf9oFkpOOKOO9WlprOgBm
l40Zyr5IcjPaGsKVt/2vaU3X7ggucMOqvbTghkAHQZYNSl3DrLxhk+AI+o6b+hihYFeQ+v4yDnoG
W7xvFtSMJ620WmzFPvOxEl41IgnHH1hqcMdkibTAGn6/VArAr3T+B5zUabIjrxXxY2rOWJ5LS+gF
UtRN8/GoZSbSJCbFcAhcOaJzdHvF6Kc8uq8Dz5f1vRNpRYHkKUHN6nEVs7D1cwly0Yj7beiUPXRJ
H6H2mcGFXx6pwAAAKJ8yo+tXC8uWzqHY3DFC1CLsdyDfKb4Hd3z5CW/HCkDJfwWqPzOnzfsopjhz
VL4WSfkmxL/lF1AM6kqmy4NFNpeRg9lZLyhuoct8lgF8O8nLaINy9BqGCZOTfd73gVfFSJ3tBz9W
XgSHkaClRvXmJ3tAsXOVgYyD8Uq2mHcXXKdpqDg/O6Snt2tyWa8VcRdk4cV8+URS0o1PDv6mjkM0
hVyg9R98WLemtyrARxDi7ECY7iWA6lDHtiCvSFfIm649+YcpgxFrkPtx/8FCCIyrd/5Q00wr5Pov
3/i+uq+gDz6Q08YK7PpN1YVW+W/RAxp0XlNVc1p0FwUvAwh9+I6a1Ld1y4Eq5wU1alIPh7skXewn
3MQ4KfPZBgEP+OBwGTzkfSv2eeiNLGi1UbgcSSaRUwyE7+gGf5B3Rs5dSokczI481LtH7KmvX5CN
cKORapOLbI1qErxGIxEJ1QHo+BqZz6rtZ2gXTZZ8H2N/Mus5ptliFejTkfFnAizT+oM++nhAz/+b
kK84OCnBSFTH4Otghml8e/wRDnSno9YgVuLSkhRVzWzmOwqkMw7Hr2py2fgqVbK0P1SfglnC3nic
2qbH8qhzPn6V/ZF/LjFBkpFinBau7wKJGIL6IwgBGaI6iYMVlHLwAVIAIOZwOmoIOurbTCWa+2d0
bzed+aoN6iQwtbUCrjr0Oy5DcIyrObAiTRnedbnkVFLQBKwREit2IdSFZm8odvMMYQ6Sparfyi60
hNkC3Fjr8SnVgTT4BzxpHSMEbBIgzmXhTRffJbeOqs1IvnEYSWlWyoh1Tri6XeV5oOEBv9MmClgt
hr9s/tvOmNnwu+4eVYUEZTL5cQFsD68tRd2biwUUHmM4hu3P5VBXn0A2FbkufnfkPm+DihqlIt0s
/GnTBRulYhToj4JtDnsXob88hhJ2kTPYIhbTYi38+UaAIVI6Qs8TomEfeKKXkjruMiuSLzT+1WRT
Ct7xAIO4Qs+yKI0GPtnVCb34rnIsLs3yff/FT+HlGD1im6XkV47oCSOyum2T/v/29+68rZ7+dQGc
532nQzyE0VmALTvvc3NPJdUIlYCqg+iZdM4OQ30yBYGzuyqssy4blkhS6Lnj+z9dwlm4/gYIUSQb
uVVU+y1OP6qWRTbFxVM/vk6Vyy4UDG4oaYTpWPjH0dGyyNJdMHjY/mgMV/j1tSd6dWikAF6XvpoJ
JWaCH94tehYhHCYwqfjVQ7eXlGU5gT/w9BL6Ic+MuMWoCDfGKx37liGOV6NsS+RJgXc61arun9Kh
m/SWeCXSiTe9Q8SO+02CyoDBfDpojOMW+MZKZaOM5jLxl9NCn9g9mks1UO+goRTa1rtJAmkG6KZG
TSvjm5cGg01Z73UQWVarOV+udqgxqqOhfK8u2sNY07Hs7PXqmxPMz9bkVXEGu8KX3gFPG0DYKHBF
qdSftemlj+PzMc2KyMu3RDOtw6wVvXHeV74hsZsShWTJLozejjTF1eZX72chLLfDcotmDx70VltO
XHD/EPAvtqlZ1ZQxOGXFXB0wPe3+RxdNu656TtJPd69n96Ihe/fom/fsVnGxsAO2Je6QXbihKRgM
iqCcujhYB5rcE/HggE5u3Xjhz7ZyR7ZUs/gs6TLIwe72R7cS9sCW5LOb/nx04jhnekqa1ILGhoFN
blgN6J7XDU/pFqVedbD66/GXZ4/viZpqiy9TqP1IAYLSWOPpzBhpbRUYN8e+HUn2UTOE0yMI843g
Q+JpYdd3MrZa+3Puq3JFcA+qrROqmYq+7D8ODbkCw5XfGoLIhd2lyeypkiwBJg7pMFJKFC5vhOIP
0npCVN2yD6fd2z0xrKBt5nvMVByceVHt5GOadU7xKmaSryS7q2TLh5Y0sDnIpDH9QSoNCAiTzJb/
ywr/bfdD20UQmhUuaDXiXp5pc544CQmuvh0rTtNvff1CY9cKi+FoeUceUilHfBWMM9TYFNM5J6CM
92l3saupNUtpJRPN7UZRa2Mtd/OZhPzO3RsPj46S+16uY8x9xSVgrtnYkccyOZg/a9a7J4oEEb12
vaNB+O6gYE9+9GOjTnNmAyeHOwTUyW0fxY9Lty+MZhgbiIe+QG3AFgtvbe24jazTFMJGVfqy3km8
qvXfeyShLnt5SrXW3aiopYiyrj0Q+Q06uMn0hH/xGQ5jXbrAyD/69zu7CYlXKJpk11i0Dry/m4sb
v+wbwURXFqEIIi+VXMtjwevB0zr3Va3diwxDhFXNdbsrojAjKz9xP3W7rqN+vgpwdN4kh9cMXb06
joFQMFpnL2ykyz8cumZgKupuSy5NhRl2HrBkKCeMknRd9ipZcKbcUdxM5q2nI7c7Dr4L1aZznT/H
VC9Q89KCv2eEdkjEXH1gPtlTaWV3CJB3mz8KGdS8RDJsARjDqLLklaB5rMw5PCKL1z7q/l36Po5e
+e4bQ5ITJ6NpsJs82TrVgEneY2+JeQ+NgRdlzrkjGdqW9q3oBwjP40JSyWg8wXhMpWT4CQ0T6Z10
VMtlNbfcV0lehrhhORJEsrxKxfzRgVw57ARsdU+gqp3PlU9ZVzARdAMVdbNQpgu0IlVVNSpzL9VY
iX+aFWgAyMtQmUqK0lCEcQhTQceZIP185lxM/k5zRmZt1Xh4Mp+c8bl5OT8umpzPArI9ercPLJpA
QkG+u4ww3tQbMCeDddaHmwkQbGDnPMYu0bYhzkMyzsJffRzeIYW1Ieg/73lGsy1DRd/sZ7IwdsxS
sgTUtnqoNY39b8VASS2gln6urPdg8ZpewjZkiMipys6ttMWEqfW2Ar1diO9tNJYAAR2Bb6w/3ekK
mEsgpnzvzCc3ZnZCyY0KLf1vmUVN8bP8o2X7HprLZQ3tAa0wRYQZZDFB6GYES1wEFsBxnXeWDd3G
aYzpnBYK2q/IqPGahjq1cgkQi5Ag93+DZxoK76Nn4RReee62XUFu6aowvgyWS82VxrP1NnIwVhJX
b9Lrd1ecgpa3uq9swKKv1e11vUFwALaopAMTeDlsPmDKzQ9WBeBZKc7NrzcU7m1WlztovUK+bGMx
Fba4o0/EUUF66b1Qf3UKQgI2pnyGFp8QI1vbc+me8DrmRQhp5pbfOXnXD3JzXrSbWkKByqVfavGZ
DwV7VXXkcOGHP+NTqJmuUCopcSBzciu6T4eLwCSuvxSik42OV7CfHreD5axzZk/TBTZ9uGcQzzc6
1ncTnsswNZ0B+XFOzGZbxhMog7jUfJ5v4TOAls/3LPcrlWIqXysOsqsyq5dKXvhw7ZfH/sDu6yf1
1GUE1DHLXPu4OOg5/FjS+YqfIPlq+rKmlnJ+O8NGc/apLkZ/W425uXHNw7dJYtmQHFwg6ohbhJK7
Hp3zYkxKKhmVsXBnH7NzlNPj9izCD7guF6CdJR2FKwZLuyDtEv4S1o2ilE98OGolK9O9TX77W7Ub
lAtNeuLspSphvlk3na6YaltGeGg/4EJVtkFGgeOjsj/QpHXyMgfDiYKu1jByYyg17A529NGjLtq5
XXm9BFjlKbY896oDIF7t3kCut8dWVY9pqIvDB4ZTT+/J3heFza0OgYHs2oJfMoM+sTrD2Ci2LOxV
2wl7tD0KKr/rxIvEG3sEYKTa41L08Ej1BLeu4miFhC9TGJoo+LGJ3TVjBm65FFRshdeuesKVinvR
OoMwXaLAEuF7vmX9FlWLl4Jyl/S/sWakSKeTRDyjBOR9tcUbP8DEviB13/sMjPviickI+dGM+HC5
O+WMQOlTGapJGXE0VE7YstsYfGx9S0Bt13HKLdOtMIZiP3DrjnVia+b5qeRf79Dn+IIIfNBgXl7m
s7+sKXRHC7A4jMHySbmFszqoYB3UHlH/GTkv/6d9dNe0hFSp9j+S6GoJUgkt/MXbPwG9CTR9nDyR
uJ5GLicb6lggud5u26RswDk3vr5a0rKGPBIflGILV3+dYAs3gag2Vb3BhZhhCSGR6Q7wdKQiY6D/
NXWIsCpOX/OHSfF5M8hPuQIvd21DhPjanJpKvSFTLBwhrssBviq1Rrv/rdkpY3l4dn0mmHYsqQje
rxPcONs5+p3KR7BnJIGnwehVHK1+L/HoWPYgoabjjRNplM232r/2VDG3jKLo2p32iETly/XV0WOc
Vqm+w3eWCnK8JICVHbYO54BRe3C+i7rt+0pydrHgvo2o5NRkmfO5lo3CW1Drlgyv+vKeWQ1NcSjQ
NyxVEWGMQ7fI7eZGQeGPqQO5BMvJykPIiB1k2Drq6ToiHrOEMLwieXjLvZE//WTI+K8ZdLk7+brs
Tn5lDTYHzavglyzj8Lrj2QjiqpPupFaXekH8Dd5sERfveVhD0J+ZK1qY9P2gsS8vD5qn8zVKVTpD
ILtKjgPARikYTSDVvsMn3b06Y87gTX1bh5Qhfe16xrMEvoM3AH0OUUFqwsy7rhfwlTxCC4I9WA/l
ozbn87qresdoYqP/OO72IPHLs5TWabpxBhZBLL+OPMJD9O3pxEsi4BSrKtnAa2zwMObc08/Ai7hU
VQkQ+hVUgANwLMuBb5kWwJsfrjD7oxfqMyzy/5w5ANhBHZ0kwjcrzUJ8cg1TLNx/Gjn/jrCfwh9N
slyup94XciY1yyqkRRFgpuhp9pMtaDk/P8FyG+vJIXeAl85qcrU9u2vSW2vygBmnja03S8KNH7QB
7W+9RjJduXOhRVAzQap5ttEfe45HwSWNKmIJ9IgADS4T4mo6ZWLRJHGUPBUr8wz45/zT46hyQSWt
bmwRUlXRgSeYTUhJ6m+G66BeMbxseXTKSDgKMluitANxE+26g5XxazGPhjX+YDauD1iuYM5uq8Ht
oY5vW2DsK/ke/uocv33j1wSVDgQfz5Og2CY55hmacuczoOzRAKixXPnh51u1oWlQjXW9PdbxKcsP
YewQljPW0Nd6NphwNTmCKGy+fC5eMlcN2IJIEErmc9QSJJE45fORAH2c/6PxEZ7DLOjf0MFsEXq7
77f43kut/emnUzlNVICNbHJExR/COU2MAf8PR8NrzaBnWOaIsRFHrDcBYWHT0zjbEcoG09qaQIpM
/R3BzmVY5jENGmrhliZM78hhKrrg0wihNSnYU+mr7gfuPl6MoXWbKIwcajNK0Mn4kZiM4FLYDzQZ
myXJBubM15AKCE+T00cnaMDs9WDkoCqyICl5lxnveyPHvxach1T2uDtiyzJZxBe0ZCF3+/u9HcT1
s3aYqBH0yd0VEjV+ZJ1j7MJYbLXhkJPhvx3uznKDjWrxKgzvhbGwgWfNOYJFmXevIEwzZh84ATQl
qIBjGUhIuu7ccs1I9eUsnDCA26JzgObU6ORz1kQYMbN7GDddlZpKwJpeWgEK78zbLRkm359G787H
65b1iz827O5vZDtLkrfwq1/N4nQNsNfYnLULr8Lwjik++KaSgSmax2EudS6raWfbWPy2wmVOZ4no
hxbrgvGQrr9ggRcquumnOVjqAyLyc5KCqkilAMNd2fsegzDz3VckwLCaN0eTEeZMxcn+b2U3wmDD
mOn3BTavGejwPoZ83QFjXE39/u0fX7jAV1Utz5kAd7V6+sFp4fzKmCxAUWyeGPQH8QzoJ5rI8IGa
DgwQf+nPD+LoZR9lbDC8JPnJpOgbUxXzgJA3Kp0erk+4NJH+viQHPD27kisA7g+vCKUbgwVyvMTi
xb2fVk4Vq7HDcPGJBXCow4Ay4ajNsGEl4Bccu/+e9iD+JfyWFEsn4MYpqlmxU3dav7GIJs4o2n2G
FNSOS8SrfqB1YxbE5v2zl5tqMsivcXj5l6yJDm+kWsKxgpVKDqgVTx2wV7+RnWt40aX/GaUHADYb
O+1n9uBRnpUk1L7LzV2in0MOi66ywRCzvOtMBZinRrTov/5glV72xImz0VTN1C9EjzIhuKT2zLTe
wRDeT+gnKFXsgTptSFckATmReytWz303ljK84y5a4lQN5xEXWK45/RRnX+BhAqsSuop1BCNGL7+D
X9AVX2ls5jkImhQwogpmbmwtHjzejUFSi8npvXS0J93LpjSwZVV3rLPZrxB8RxpbBSxtw8KzoFzv
T+rQhibYLCGAfKRounPn0/XUNvOu3AvhAmben3u6RsWkLfRGvoDbkHdVna+vY5huhRry3x0QV6Wk
u5+x1LzNuo0BiCTNbx+LOyJql1A693OYMnRznIXbklAwZUXBM6Vj7O0SCBJyqC8mvHWgLfTzQwdw
MpyFC8mhqgCy8nw9UmeiKCFFCbz9+HuqAvg2qybukV0qiCHZnAVlov9ChvtH+gkzedpw5KjraSy0
14lGi9+ljWmKGDYvCiJp2XDJSEwnyERcG4xR6xMigRj0pciWNCAuOLCI4cby7gEKoBurzgTdkWyX
U2J7WZgg7ACNICUqbjyhydKK0qlpSwgknMzw9gsNYK7zqurfQNVaD5aIqhSGAn/+8La3iPd+pB27
ULvVJDDLSgQgqJaYTN3I3mxLIUcx5Tq8seUvpNivcgPnBXxkYXhLqTyotLb6d7tNgihcVf5qzhIW
yl4YJ/l/z4R2FXmwZQu5rI63RaOFUfZbbwgKnxsRi7dzAJGjhvwF5vyyvpVD63CgnIaRoWuXqvEe
D/n8nwlOrk1scxQBIInGPwQd4UujVX0px/twfEWD86J15Csefo578SW/F4mjvySWjhCTY2lFspGn
punADNrDumUYuXzyI3QVLhF1e7btw4tXImU3ONj4TlQB/kpqZN2R9BZMm3hrd7IfwR+ncJHsyAQC
EwNfzojYP/aJuSkA7hHrcbpfRyyLy02g859qJQA9JfoonP1C3WkAhcaWG5aUVgxcd6g0JysCa+7Z
GS1jBhxao9jIYSIKkUsnvyB3jQ47gGwKuLgkDYgWiXRDIEnaoRv0FlwnfcbuPUQi39nb5yIeHPT3
u0tjlXWWcMnL3tbz+fp/N82YkgUr7vjex0nZxj/tifnjKE8cwHx/eTSbF8Zt3Ds5PYbDIMn24tzh
Sc89Kk0UOl8TEOFykfNlKoRxjVJq+I94Lb1maI9d9OkRHYQ33yvvTgARffQf9sSnPqNJ+b1TpGYZ
5Jfmruke+k7X/XjEu9O+cBjxugFqYa9wx5OmhVdJdkjDw6muw3ZY18hDPznUlp8FH2Ik9ln2BAYY
qLHXY/LBQoF8NNFyOD5GJh5s6n0HwL/AeQaMk3De2pZxZhz9qiPDaUyme9x1tWr72Z+ChsYhaDgy
CDXTCY8xOURpsva3SFWtO1i5TbAPjjzgpKYTd/BdXnR01TQxpiwxTDMAtBNNUeWCFIuEexUMMZof
07DgLxUDDj0FrECIfwsgciADrwNOpNA7xYhQ+i58pykl0AkbENVXA+mlqETFAd9zO3wIdQWNxVjW
oJ5/EVWREuZ7zvLtVC5CHLVxR40Eiy5lhLtaLmmZjA7T8qCIDdOXflLKFx26RyVuQSk/1KTdBMzl
DckUkWSbI2HXYjeffVlqnFSTpUyYpIW0yzzTtMjFt5zLUgcJpqF4XYMhJd7Wo5Y2ppgd/SRiNImP
8XGZVymT89JKdHaqj207nGImbUGXDvI+T9JHqTvRH4gsxG+N6hJU63KOEAon8av+8l4mUyy6ZIib
LRlFfWaxno7S/Oc24RGLbDF87YyZvYI75F4Tco/Yw0L+VkqyryexlOS4yeJBrjvhu4/dTSSXLATp
hMrs7f2ICFCOQfNTa7h+YZhUi3xPf5fD8EdOJMsx7/ar/C6Ne+QRvqRxQ0QwzOILX0vr2pqpWAkb
6y0lqCi+o9nYqLbOs71YO3wKRFzp5SXNiJ8WlHPJ2Jzsy7hiqC7nAWlKsA7Udiqx0xveUJC5dwrR
zYeZQVPBe+Ggh8h3lGebAoE6mZeOY3VYvKl3x8W0E2KFtNE1BsssItG0E98q4IDw7XAX1cPgxWgm
5keuQiWE/DP87dNuyoteUYuZSNHMBfNzVzVr+EMgZ+VCsb5oLoAEeJzB3IvvYT2fEEB+WW0QHvL7
mV1vAUN4aDbr0+k4OnRT3LcExYr06rMfbvAs8YwbIO+vEL6WNGTswRL4p63UTaHsVBkFUwK3X/uQ
1osf+o8ylBWJBPz3K2xJIeWs2VJZg1XlBzHipHCm04hDAPPKQ8tQMP9VsyZrSurEKsQfZf+5SAnU
DbBJ4gReCFhllBD5Ka/husAaU0zF4nt9Nq/mIlodg6fKk9KmmeeSd0oHEwQxdFLzTaUMmM1S9s/K
/ws1zBYc+SsFhJsq7c0iVAP+d2BACwrhHLCSRi9KVb4bAzh4cKqsXw8LEekHYrsuLKyw4ldcvK1+
0UHzCRQKkyz9Qx2vJKEoj7X6c/xufjdjJX2HL17jqhjrwEvMqW06pBn6kDjivAXAVfNmaB2rEZbT
5QCKvqf2KzpVz6uhWniwu/tncPHysCbP3Dt7MmLMwz8wTmUp983Mh4VBKEcXJ0V4d0oowhDsV7+0
bQgtk/ybQvw909RSY00pseAyLTQN3ojKvMwoRiy/07JHUEBdJPdAc3LmIukVPBWKauMLZM9WOEEF
fZ7O19+YsUXora/bALsZkF4gvu2YYS29Pdn7A/XWNY3/m0xOnA5pLjT0bGiEILbN0G7fZNcBzgdE
D17Uf8ZRieKImZnyx2FCAKoY9B9pMGwYX6PKCAXanHceh9HI8/v25WqOaop0pqhb0EgT0HrEvS0n
yF4Sim9YmwTW7U+VC9mzmK9IIY8rjWNsYQK5iT5UO45KRINBPcmx0eZKOVL3fhVoHf5DI65u7H5q
GymFh/BEvaay71T+yHYPwkFS2UFASgW1y9jE/nrTf14gSHCwTVlbkEzbIoXr6/QN7ObR3q51yD+P
O14QWMkebUSt7jgrlndyvto7dsNrK4Hx8U8GBti1Eb3I6YngSiN2mObFKKXnLMrfIuXmO+br7736
CBF1+rXef12Fkz6P4oy7cS37ncWYYCro48x6MFcoSamGc4fCPtYsz6pyugLEqD6ixbN+52l1702S
dO9o2kfXfUJfV7HbP7I3gV9TarKv60tse4YIjXeduTpyxUrHFPve2cw6bpBCUWLK+RfgXkuFKWc7
UAZscbc9/Ebb3y23jqHtRhuBg0lySwdmQi7t+kENAjac0fDSb6BmM+HAarDEyFdf/w2VyMtcnBcE
2TX4CSPDp+DAOuTNgAkeURAHcSBypPbK6usnSA7wfUw8VnttIifzFWzGTzOO+rjsBAxR3LA0DHYe
aSbND2LcJn2YeYo8g2yJShL+xUFn6Pyh2RuR4m3vai8fz4MmmtoUZG5Y3iKhDoUturCAwh4B3EJw
2XMn94UeWPZFVPRMrJHXmOPZ5OPn59dASReXc+1DTm6CTrUvwhAtWDy+l95VoNnJOFbuat9WfGb8
fhZG10+iWSywqEsFMY85brS6gIf+z2XaVDyPGQKzCdlNotOjRdlouMdUhbMJxpgQAREany1WVjKi
wATdjIN9VMFdxcGrLOyFLD1mt3A+xW4O7AIlFK/+pFq26BqylPlRR+z9v9XMa4pI5irXL237aiqf
CKjYOXmu+Ii4avDftREwD/smsY2OqRIvvmsmYH/SmJGS8Zmd+XSG72H5D/7XWnFvtgEphfb5sKh+
WDJTWLmLr2Qkgl/sqx1TvxrT2dFW1yzLwefNQNIWhQtYxHjaFaXxFyyx6Oiwz/QRLpTOn7WibVbF
0FQaHgrWU5pB1qMFzwIxmL8XvNl562rIDjQZmxSH5CUDugLa1oouLdtm6oyHs8UUmkP8Oz3jyfFz
kQFw9BMu6KRYNHPFD3isl69H44po0bV8fiC1rkRLOscgD8T8dxzO/yCeOF6jffzRNU3sfcS3WQmO
RgyHDdqqOdtF+MdMk7IbdixSqoczjhWg6zF7jB9CGOL5iO2xfMpF/GgnFAwKBvNBSXDlL2c6DDOQ
tH6HZ9hGO7/xC75vpGZR7qrcUQfL4594NnqsmpCQLKa4k9c8Bu02LmlTf2kCf1wp/9S9SIIxyC6B
XUeffE+Gf4HSniDLZW6SpM48JM6kKTcjB+TjkkF/Mu0FCdoSd6kivO3cQd/S/4/QkmXqvv75/4fv
tWdqDcLWVggxytSKXwOm1gWdgFC4LEj84viydtra2VC82VBAOV6p7qsx6GzdkPk3CEsT9DPvEbCU
Neuh1EFovO63dhGrAYZPmLfztbYEu5ac4EISV+xPARi9pHFl7j1IJw9n8SGvSsaA7wX5Smja/SYz
u7+bRX6Kaw7bGI0X5QYdm0lnYZRUNoljuK7eys/NEccX33mpqdeUglozPSnmcw8TSM0toie3HPMJ
qzjFSlsW92wAEz3sTiPoKI+CuQqatWzBsSRTerqYNOPoe7zGgPxtG7p9Cy6M+yeyrNA/12mhMHd4
kE86rhaH/w6ZxnMHLbw7NKfaXQw0ZeEH6S7qfTqwk0XuzKYWdkJjey+Mwjt2NSzljm1ObERdbaww
IPpSf8ByFy8vFdE4FAuegtWCwibUQxJ4NduHXW4vM7IEmyib045JOq/paTD694stMjA2k3NfUBNw
kmnkA8XjswXqJDwg7TCmiq0eYrDNFRYbtKeUHhBpVlmeLo/WTsPSoHV1VKwuG68oZbdLROZttspl
qzoy4OuCKVU6qWsCS20ZIGqd4Lhov+1/gIfC6wU2I82exbmUCdz/4U5B73PJ6XIMUZBtIzG01wsJ
poVoUKajL0c+Ywgz055bpQb8dcjWTioSoFwFxKMz0a2x8J9U1AYrlHZoJrwbMuW+xrqgEdt7ivLo
jf/DdvrrwLN0hpn3AMRA6t2xy24+8eX7gg0EXj/CK5xMrXSzGVAbhhpfanEycNsiAVcD3NAdWaFr
WfBCcD9hc5oRd9cHEy8YKDpDlOWjoTOmDbl61ivfeLQZ6uEex/EYGfnuBbNo/RV68balxxNMxyog
p58RumlyZfY3+GVJwEqvqvR+JtEuDW5sPQFzuSxqJwuWqq/iIXRJcpTTSaEI+SNpkUC0hFHTLKEF
Vz0D3oObEMtPLYIJizgz5A/U8lvwpUMCNbX8wJQsBPsDh7U81MpsDWvjgmNqAT4UU5ayIeGfGIJU
8/yMyGypitMwUUlJfg+pT5SPPQ0Q88A7z2qVgeXIxDsMn8f37ZFP1PtD36KpYMSVyFO7UvanmPNW
ucZB2aGGzjFkcBtuDJQDjKZPheKJUmjD7uuewbo9TulN4172q6TK3TGgKEjMeub81d38jD3uRmCx
PH29mnHrfrlMJXkT3MWh+SA/73/dOdLka8cUiuR8BKXlewue8iuMqtkv9xy83Cfq5OQEgX9e0uYD
JBkSkPx8BNxmn5I5hzQmCyDuIDsPCFOaImj4jTDysYsk9tzrZ/m7YkFEGJWIEMen14lOK+59K8Bj
f9IcrZ9doYMKgPAm4L1rsLZw9Q/YvlTstU0usywUnq+eG3BVqDL3E0dqI88Bl7kx/Pol9rIi9YGk
U079PrXZ+l8ZTJlS3NNq1uZd4sJdCzbCmizoPC5MchaTMe2nfMF3rVaSYbU2ci74oHRRx60iRFUa
1Lkek+tEU/p6MFLKIwQVHQt7cRtG7LiyCXBmxEJiU2nSIgHG78jd0wkijzfRWSnzPbsdHDgXYzJE
H6gfcbbjCqrJWUI6GQGc9P3I/kL/HDiUP9BqrvFyYwGGBQ+DNlzlUlpwJJgeFu2/nV2QM3CovnKg
HTn/Oircse5XMKuui7zuzvvDz43cMoRj+n/salt6mhJSu4uwYXBF/Gh4bNIn4EKmN17qqNxeO8LS
m5ihdyeUHsuOj0GGXlQklwXHlov+rJQZLDUGpFiBy3qfT1K8tF7bH6vC6Cojjl+KaSXW8s0hwHMF
Drz8AO3JciSUkovaEY+2ZXJsmiG85vG0jtMwGfNetDyr1auQq7uFsGs16VbmimChKnt6h51Xv050
an/hcfZxXL87UGqAaFHo4hhKKnZpMME0WBxeheYiJK2+qXDcEZSEkXu2mANEbjEwQGIGZOYi5DTN
m0lAaPCH3dboAZcPS3WkQ066uNmNnC9GX0KhBmoRhIHzSq6QjjGWBfzisXtwWaAxAjqyyceWUgGv
keq6y3ZdsXEHArERrNA++wIWzVcvFesz16JAg+J788uBL+atEoPJ+oDCEHWxLGhFjXqggF9ur3oX
2WTXqz7pZCgznVoNANvcIfVJI4RlFMDW5/7yakUQ6/ZDEqV6yFB8+A0lv7gV51dXDpYDjA9xMg0Q
0EvKVBirfEBfIMB/LAYX7ggLl2kRaLNIKyBy/AlYPEzJe8BHHydGZFMz7hXqU+aIlup74cZ0Burj
logHErTYzTDSqS0FctAsKkaDEqzw4P5qWD6fbgoK7dND+Vg0bRgpHs3KYGINw8ZPeF67kLAB2d73
6iCuATl9hcg2M5YnmX3AeH3ehbEA+R9nLzOI2bRXDg9jdzqaHLdFIIRPtZpHtgykahYPxp5tuXGo
Cl99GQlAWkiT/c2LfdWqfJC+bkfCS+s1djnr00pAkIHUSsA3j+jldFU96v9z39cqSzeWL1CW/Xnv
hcdWpbbEdL44nabBUAwdFb47D5/wrqPch7UO7vXJ+Fs60TgkH0gzKLuH29vm0VSuKOj0zTyJMilv
CIvs/S1uVlbS23NhcJrJQy7VKAEDYZY4yslkLZkV0K473SzVtek7JbWfXs26vIXGVtOZoeTDakRi
S0Brz4Tezw+kibXdFsl45Vgh25ZpdR0oXjHtBRzz1wv7i+ZIbVPaSLNrOBQ4WBi9havAOz/gHo5I
5piZiyn52glmREGHnevtmAGcBTAJwlgiee+jLL2JUTwLpXofAdMjiE3wDpC08MlD36IZprNRSvt+
/oAyHSbiAUbFKwTZY4XmzE7FkXwSJ1xITBFzOW6I32KYBJPUb9Y6tEYQ/ExsaWOvckfAgV+ZZkrR
7lShWDQ8d3oDS9lYi1lBsvlXUpxPNXyZbcztxUXnrD6RIJiKrFmCRI2+FG/1L9nli62XKs3R0yh0
/F73343aOtFchBjCW4xel1bZ9RC2UNev85zL+GnLrnCtlwGle6feTgWzoeQ/uBslqwQRwRPQF0/v
ofzP01rj37/Qk0GDnE0Gck2+rHi/zPllU5fK3THgw5o/ngZp1XKlUHwWWx0Xrfs/1TewYEAvA1DW
jYehlWbMipufhOa9J+RAzCtKvxOFwdIxcEEH70pE3B8ScOExo3kGZWVleq3z9GWEC0GXmbUAQsip
RLtOHkf1Egok/m32V/OeK5sh7cFU1wQFBEsJG4n+KAQY4j/QXiSvgaY7dEJLx9huayruZ3/IN+p2
GPQU0blUw8voZg2zTyHO8EQBLXpJCBpJEH8yIBIjuMRs2sxScx0Ed9MPg0CPHaelxfMp0aSwb6Mq
s7WP4NCN9hS04NRBemIEYWCbsrqePyI8vqlanZqqAIxqamUMTIN8waU3LPZleoHafk8a8TJcM5uN
Zi7VtgyZirgZLr/+7JdnfflZgBHUs/ZwBGrXTl3jc6g9N+Lhpgu1PX90QO55BEAUrfuqYiVNmCzZ
ZqSy4Bs1vq3V2GIy5CAG5EEl7dE2t7WttvkYViWLYSAJRxHYs1lmhOihoiT5gyzO4XaZsqcOPQpb
mC+l/9d6AdwCJa8o+zO/e9q1sqvKatJ6GMjf6+RF3rS/EJAgH1QG+X7atVF6XCYryMsvkXVeemmV
3R3XkxeRc6IobpSwrxOkuzxGSdyO0b34SmzWF6LByCp/eeiyh3OnmUCxsEnzRFtg1ahizi4cRm3I
bLnMFPkIK/tbaaLRRFfxsPoPpD0IEmbhMBO/oOlHYvukqCBMB/AJNoeSh1lQSNAwtF9lVKTjs0iH
sPVAC7qg3fE4LuLuP9x0iie2IwAMWksMEV9OBap6Ej2CNR01BCLFLQuIYdNiuern3/vof8GT1D4m
7yWuODlD7PLz41YotvSCDNKDoAODpoF5nHD8JhMnAaL8lCBqR+hzxQXRsned/uezMmLlycMa0fMU
53SMpDLUedsZ+F40i62ariBAhx21NWSH16PoY4v19VjczGhbfpK/ouzxtfZmcsy0DO8nxBVn2RJY
hm51wkE+HqkPpYy/ZLFYJZ8BUCnH3hao8lwBDaRTAVOxZSW+FrcHOIDBL8SbcpfZMRa16yjp+cW8
ZXLlKT0Jc5Ld/Y2ngQKnrwP9D3SXkTv69JBTzpbQkOsTOk71dH+Ptb3Y3uzgLRZKD9mMCSrHAxB6
iYz9Fa3T49RupMIIfTJbxlP1lE7vZRvjgq/CWAw2t0XSyzYD/10RJNIna5O6SAN4Pn59rqW6IfZQ
CbxvVaaG6FumFh7TrXGFpDjtaM2tBmb+CJUVanl8LUTuQgtzxn3LxpM6qtyrRDCOlWSNeq8dXXPW
ZTvx/z0Hrfawt50CMJNQfkV0zGZqQkyk56EBvCpSfjm9igWR1N1PNlIoMNyPtOvHO2zEWzRik3VO
s0YtM8k76mFuZQUaOsd1E2Jt2kXtjYlFoxRH3bkzNTSmw1pLQlMLfN9gChr9yNgvINrTWwSwMEiE
IjgxAFB/eG1meGHcGjBWvkkGMFHSkd46iiybwNzfjY9D5S3/PjNZ1DahwknuVI9C2mEes14YVYy5
8Q/9sKJPChKPwGQGIq5XoIupidUZwhJrMr1aLT2MfCen85yRDDDFUetolUqANNo8U7PnoKh68H6a
1KuEHYQHfiQatVsDomYrmFGT3+mQFNSjoss6aDlnf2yHVPRCcLlSMxnTK7otdzcam83t+undS7Kt
Q9s5pb+F7z1Z2//i/Uv7KlhyvuzVveWeyJCToNIIcMsIbMK1nDs/RHkE9DuTLUdKK+bVbFfn7+EG
3x5sQjeel6DmNpENmmCrsAr+wjelK3glQnbzaOvD6cExzh3pTPfMobpLi3QN4kmzIJjS8IX90Suz
7nzd0XS3QyKLa1NKEy3THTkhXasHeH66JksI7MsposdRc93yi6hFH3ni1qT0q7MbZvgog7h69kiN
O0+5eF8v3x7HgOVkotIDwwfW8OkfpitT/1wK+JRaWeOZIUy8eDK2t1nIyqDvHvYOPd3SuD1+Tf1u
XjO/p783S5oWQ08hq+nPejZS5zpVOPHG3Q7wr7fTm07PyVaSiiVxU6YdP6bfRfFcJwb3/B/Ol0Qe
xi2xNVG4w6Ktf7OYROTPbHNMbWp+oP8qhxDlzvuOp5mR4nDTOGoz2QHsqPguEKcKTqyhSgcPRDD/
VKQdGQRsWm/4Ds5c04kxsPRbf8qbc9oeQ5kLeaHBn5fSGHPdVLQNTt0a/YGiw5dKJ9howx9+cXDE
k1aPSuho7vhJlPgBUHaH73udSVi3RJSvLYTAaWaaSIrk9+eCEOVdZ1+Qvsarm+JpMyR9KQvUpGZz
WPUu1odciBOebCAkqiJc5RXVWEZiOe0M74P7sWS/xPmKuHUo/lMCkmQfFy1iD+voiNe3xxnlvfcB
Ln+xZnhPrfbpPD08apUP2vBtcRzZNqjqU6UrNFGLyClPLykVXx6tyga00696GAX5V6GI5oq1f9pQ
bHVIHL1JndNw3K9HozFpbHFgMjqCcjyHwclrX8LKmBxBYuH5OXagAP7L4YPMcnDhlRBA3SZfkk1e
iWi1V5YKYW8SNHK80uz9N3UK+Nl07b2+pShNdFap58ozOUbp+0MSL6LLCtMqbUEEzuIdHf6Y0bvk
9NynG1Ue1w6vNS4sx/fbkLFElrtiMh92Y/BzqEa0P98mREs8doOz3JEnYVbK57zuHvdmusbP24RM
d89l5ua5ZUENgmeKDRTu82wdfvupD3/ym1FcshUeekxQhJr5P5DxWJe2aVUPcVXzO/cBvjZX5wWV
6EwQTQKHzrzlgFJLJ7AaN6Ba3hqLCS5ZmU8RW06nrV94PG7Em9eDmrdIVfdb/11B6JcPMgdtLVqc
GcnA+rMhZkTvhnMo2R29J5ResTlubQieLAzVe9IC4YY4UduheurzBjyB74UkXOgrxNaIX2yTUpSc
Q+B97DGiBwpGqm1m8DdWTxjJ0ccpXrjVi6PNpngGpzASWSfXfmhQPAoTZGTw8R9DIIjQDWrSH5O5
J90zB80HSToGZ3NxqanU6XMyUR04HasZ6tW0IqTxCErWMqUp64bwe0tun77eksFScqJYIsprT5NM
CzUa3lrcQe0p1X4uBqs3MwzPMV47blAEtSeHAOj4HkXvVSOjIDAu9Xqac3PZURiflhPMmY9Q+sGw
NDN6m5yJt4EKH8E2xQMwAiw+rszxC1xPr9a8afW4etvwZU2Jy54ZoDH2Qf5kmk1ql9jkw0Cp8e/O
NnByNCACIh2df2A1HtE/mVo6/oB1fJPaAZnoXnrHin3/SgL6rPGM1V2QRiTBlj5E/0mCMPGrAzxR
rXAuhdHd42akkH7XHz0t77gfLfNY/wpgFprJM54Ee2Nae842EP52J0IuZcUT3ugX2IXZjUpmq0qX
u23332dYFcqmnEgRrCszB+a5CVFFQyfk9hCovwwkbMYHyrP5r7z1H/Z3shHEBuOVVKurfyR5B85h
6NkMlGhyS6aeRYc5hLx77pfU37XDEHF4XxIojrxrMnnZUecwDebW7k5RwJBDhyHvxXzb+a8Dz/jR
7xhf0Ej4dT71idv7GVR01W/CkvG6o1VvH3JO7uvON+aPRLBVkAT4+Jyc8XsucUpFKoQ59UO4Qsdv
dxNh14PrxPoOdLmt5+kITrA0jXmdkOTNrCUR2eBKdQ3XWU4DUNRRV2m2jqfoqnHPGwxZTHu3A7tj
MSwL6d9Ng8Cz8h2SA/C3G0O34AIsZEq/x5X2w422CcUJE7AwivfC8aCv7NKoVW0wGFY7ukVNlLnZ
fGJ23ecEBvcvf6t8wyWpDkledaS+Bl74M79jU4xAVXvFPRjNr3G5GYK+QzEWraFXy+ew8Mpk+nOC
jHvQezzFHWoZyAIcFvovrDmnLxsLg8QvuqzotZriOULWVSfA+9Nlq2iPlEdTTYYAkGRMDwvP6tQ/
nL6HFW4qruG5s901kniWxoqdilTuQuqUl+iTnmr1UjGHvykGob3/yFe6BOy6agCjsseL91tC4RrI
1gdt2JnM3Nw1E3sUuDVHf/q2AoFCG98/qmfTMsCpmN8/8QOXX4tfBlObL4KxsrklFzkzbLu68r2x
ejfqhC5XR/E3erdz2W601neVj8Nrw8Y2PDZQ/JDxN8kNck2tVYodp4BHFce3/j+pcZwEvrsOud0/
pcfcZpeacvavPIJp7l8EvWqGgW6vfsy76yPzjzd8eImNjdhKT2daCE8FgEDRO/q72p2HQ8oNXleG
1fwv77jWu+tjLiqtEfVv1ahUMZRvgiWcLujbIDivlhrEuEWPf4t8KaCcwCmK0XBZC9tbT4u7xfnm
FL0E/n48RyhcBKLuCY/5oPTljVXE/lV983tqI6Mz+9UG5quva6tRCMiyuCaPMn9mNsRM37foYSaa
XEHzDyZA4UXQFpLiwxCe/3JnmVTpBkjZ48+D6cki73tbCNeyt7HvoazrpeN1Awj4yHyIKKM3k/Ql
6Z3/kP/kBySfUCRQ6EEN4une62fMtvG6STR0yTpiTLw/wZ+H1A/qXPy7CAjOqrN4jiMl9yMko/dM
bMp67dZwujmCY5Ol/IHzDaU5/uSpxF0B/ItsNAUyjKagpmJBgtpc+PP+8riRDT0+k3w+mXks7kWQ
zpxgbQ0PxMb8zcbZ4pK1BeIrvsTM6UqQ9nXILfyh2XtgEMQQRlaZZXBBzbTAyjqxtdRaDGfWQyIM
WZNk5roHnZUDoCblzeBn8nK9SGvqGQOehc4CAy12BbbfmIbdnuGiUBjvHpN2O8gZ8uALqnCAY938
yvx57HBD1fcADUwInA6gn1Tk3QYgUOnxf/jOafqnAFcmm24XXoAjeKnKD0+b1GPu83y9oi4pwzN5
440uGIq2rkq0e60ABI9GI7tcCyIdg8UrO6YPBGh+lFMaF3ny6tZOe5fgruXg1DBO89ZTuBtOcBfh
PxVoFVogzcbYPMIlcBiBn++vdzChoAIb8SSy1vIU+A3s2GuuUimrsA7ZQhabkP8LB6IuLpwb/aZP
W0rI85EDm9HNd6XsfUedHMYery/pb6Tjv+DYXIWb2YsEWd8Inabd9G/IkDsMZCd3wsPf0+IcxJze
Ly9a01o3TCCNXk6xqoKP5TrpcX7u+LR9XUfmyw6Tth2FkcTG4UUppC3HbgdX6QWnDrzn55zKr5KL
ihZG3VNIQmdpHToZEJuVsa0nEgLKrBioAyeGYKqhls96rsjfPlNZF1VdBdOggoLtiwq4eoKNufP5
VYLHEecZncX9Dh9uYGK0IxA0QPtFhu7fPcZ3XG70yYOYuUwgPWUhIpe7wls+dEhJ49JtpkeqvyOo
x84NucVI+0wCHrHS54ubUQmZ9BKDcu0DcHmA1YVvzsjFd0yD+AOi8LHuVsWqqaaImNZ3SHo4YzgF
vi40NjP9fWfX22KGmi6WJpfKa0xsW18RKkhwlwoPHzuRQm7423TEyYLUP9Lmb9Sua2hmfAsIr0hE
GY6trlZcPbXTYzKdLd7ULCvjcKpN307leamdsVHuoCWHVPWdbN42QYAP78eZ0hIIMLhwjVgbufka
h8y7IGb22Czp0WNhNeGlYcwmjK8aErItj+TkNyGdK3rxzsZij0FmhZ12PjMvP2JlTvhDpRz7xzy9
TTYzncw4/dOXd4DJ8U1T80syr3y8Ix/qnc/1+unTjhi5HfH/oakMSAPMuKm3PkATTZ5nqmjUL7KP
/vaV6n9zv4sMAC9H18zs1u7eptKIb+W2yZJ38mFAhBDXegWDWUWAq48ZAiGOvTP/J9EewfOcxy6R
0CpZceOh7dyT4FWogY7zikdfquETuae6ZB3RQckMCe0hPcKfvW5IbdxqtyfmBnmInrSi4oiTKG4R
PCs8LajlGPZAaK7IHEBkLmYfP8YudVOsF570W3ZL4l5v4/+4xMMNvmcwswKykzrFffXlG1pSini/
bhlZWyRfq/sad+h00Exp8CWfON0uYi/wJ/Gw4GcmmJ6SmbO9whCccxmUNBm4sY1nZeXiXxsper1r
6RxJ5f5bBLNVs7oMZP/2tP3jkU+aNNkZsd8HSD6U0Giuhy5MztbSg28426waM4R3XMu2sYwKabBF
i6LmevtxwEdGXEJWX3plQQs+OnCU7S0gynuTz4H5V5yqJYdyLt0vDEBEhn2LoXLJ4HESTh7lk3Q8
anP3B69E7NOX4GQ7z6NRDhZwdx7ZlXP7lnezoMWZNcYNPGtCueb7Vn1TTywzCjbGCy+OGxUcefwV
5M8+KGlGy+gWXhv6NJA5EAG5fW+Cc79GHcUMrOEBXy26QRF9SUi9qshbz8Qv0FrmOLl4APD9mR1Y
CoE8Wz4wprwTLVuSw0guZxcdA3Jw5Hb8nIyqr3Cpkrty9MYixgW9MISPIztmoMTKAoMxY/LnzZbS
S0EstZTeMECF2xfZaz69utOaDoOMCUzStE06a52BfZ2JDe3PDLioAgtvhVaV36L0U1MJfJc166lU
TpmcK2m3F2MwmJNb3le+kTDyUUOQU7rU+DG0k1fO8N046aGGvuznWXWLeDvi4AZ7l5lzG2yD46vZ
kaYe8efHvVkYWq4+Ch94MW5RYg5ynj79n6mxOIcg+0WMMSzPZmXjN7P+ozK1MeCWvgFUJMtxLYEL
xdX4nEzVpTMC5/6FF3dEjWdEfiW2U0N1AdkdLKJ0qbbSaa531gwgeddfgzFhXSCOi4s04Wn7MReC
jLJsOn2HKKaJMGYjLijgZ+Ahs5J77bU9N+SD8r/nvTDhg/0oqwhDargf7Ok0Y9CJ0HFjQjE7dLVG
un9DlvA70Etgnsfp9NGhMrRI+L4dal2s5ZCETYGmkJrCslYRp/d/mr0Zp9p0oqohRK5kqltd+lZB
asH6ehXo09lzuxjvm6GL3WVF5JK9oMtrbFPzpdy17+tCWFHhNw8xBjtR6GAMOIPNfpcnQh+sj0ki
xF68HP2dhljhYoNcfUdONkrwEIeur0bAjKMtiCH78Hwnx+2qGlAlwIFW61JAgxsas3JJrQHDJTm6
lKJ7bSKdQ8YwJn8nARvmeqfzVlLC6aKBx5FT1hSd1/R3XIwvZBzGQIpeiTGo0nE2TQEGqHzFbdnP
ppXOsSbYdXj8e5KizjT2bLesZzhcHhnzJLV7f0Ojwg9SXA9SlDqfiJckNC4s3QaIP8osR/L6JvPN
cUaMrEll+FQ5wS4ZcZrM7Guhe4JR4XG6auRRUsGvXYYSlnyCgT5tNpbZEoo4Ro+DHEyHmMKE0MJn
AcdR9xrePG/MrDQamQs0wqiiqC7w72rW/AR8xKgpDaV7VmdT6CPApi2ZcVl12IHP+XTW5sMCCQ3u
P7e9llvpIl0Uni0OW5nAuZltL15oUY5dfbX3tEwDyd3A0RYWIuJ1IHTVD8IAvxg9BpdHxh4xqbc/
/u6WqPW9aSU8ey7PGxsQ5V3srUtqefT4UFq9HKl5nvn5QzpESY7K5cNJQMHrHMwSyk5IiybafPWZ
F0AJzSvCzTkf9H9tdfh5GDiLzLey0zwWICeYEfCJc0x7QDPfpyd4rAwOQCf9uKtQwGHF3vBse/Zi
YuiWgxSTKqavKmzAQvqj0WC5Wy4YjrdIYxQZ1jHduvXQItuV3iQQB+G9rhUhYg68YgWxpeyWRwAr
re+R0j3qLV4tCB3Q6M8NucvHHIrkWiegb7s8w0WDn1MK5Ucqk32FZx2l0BHyRXxS1iftAOcqoS/b
P/eCun65msONHE5bEKSu/frUckoq1Yg9tsjMEcwfs3milcAlClONhTLln7PHkzopdMAVBHkJIONU
v/u6uvm5GkFZV/D3obf3/4cyPpqEAZ28/HA9nbvr0uto/ulOjWlPWzOYUz9sKeAJTIBUE6tavnzf
broPTaZhLxVY2pT9L9m2ZpqEzCV8NCw8BOepyKtUjDQpNkc09D6T/NYeRPaguGAd1V4bCRtTfOpU
ajF+0BnMESoqlV5uj7nlcJw2jdklWIVvm6ndy9Dwgu3zbYpuUgySvHh/Gzy6p8GEivAArhOTTNhP
ShIdwvOtf+cODRjSDOX+v7gLdz5sbh1TlYMcOvbgZ7Jd0Y+rDucIibDw+JTFhgG6AWvqzJmugy+m
oxuTY6Q41suFTeCvZcF96FEpB/kuIal7C1n9Q9kjZ8auDMjPcD7TC7kdmZlLhVMkGn0Yokl8hXtS
vewOyQwjXyH9P/Y/DBY/lQ729RMPh5zXKkmWMyJxokeCqU75P1Kj/FVKMUW6+r3fsymy+earEaxV
+hRUYu+QODQ4mgM6gIHQbB6iHsO/WZoJHPbAhM0Sy76B+g1cAa3ifBC8GkqmC9pdQprMXw9w7C+I
l4ag0HC7BUpfqjtdhgZoRDGVBgZ+IDqfpA2lvQ10wHGSMGyutabtfxw42O39xpjA3s0KR3hFNzJx
eIGr94rsN762aF7BUKm+4Ldjjx8grevs0goCPRMP01O+BtjEh1SENIy2SJFgSj+RQnyBtDW6g/Tc
CMDZ/cUJ8mU1zYBS+Q47tIzaGokG7CAC7N/QpEpaNXwlhE7ZdlbMulMd8m2Lg7pX4Yycg/5O0TEd
dQfw/NMGpYO8NF8WmfyGDFwAIJRNrbtaJo8UonmzIl+D6qpnTJsqfZ5HRFKRmKaaPiE/mwvMBf3y
hU3imp3fa1KDjhdwvIB8LKIO+hsilwfoCBfprmI0ddNMqB+GROucQAtnbpo8e1M1KYxJhZhKQzDN
uDLQ4DVcdY8jJkU/xBI3Uaup35/MDPYWpKwiQsuh4XE7eV42FKqS8CFYOPjC0nmBEbOsoA2l3xNU
UXoKcKw/puRw1rj0AXjT74ebtnwcDBiI6ExxE9ciwDAoGxiU9sOcvdDsbC/qlLXua1tag1tXKZHf
/1tXECRXtkOI1E0uQqpPjNdjRVMZr/rTt2Zxb75YQj5b9q6ygkOzhiB4wJVj1YyKadpij3liZmZb
4XawZWCZd/WHXhZ2nQvcVbxcqzEYYoacCW1ZORNPfgymPPOjpN+N6iGK7R+yI7XLcotmq6fpuh3a
z0ahY6NLZvtQUHRLHErk7k+rdjxfANfXVmD04vcNcKOmlzo1LPik9sL4bAyEDgXuDGkp/9zOQMxJ
rEEKM9oXVPQU/DRgwUbBrB4O1uSFLQJaFLRLqMHZLI1Aae1mlNGCMIq6uFDnoFJevmW8Zi5rvP15
e1AuKUDG4ENDJGh6z4FN+ZVxBhPNhDdHsdIirffo6Pw+qfiizHIHYG8gEfY1L6rKMw/t40+SO5vs
gtiOnb26BckXViWbajDpCgh/CRUH6Swt684PWf3yd5Ptr7UY4ovhtFndZlp+ms4nFPVXfq6EpMkV
szQ6FhquNHdQQ/tbJDbwi7dIp5URYF+pT8t8hVqHwOke0oXeg4r/qHYCjUhfyrMemmuajMPXQ4sT
QqNg0vx+zIci9Z2n9UGqC7XgtX7N4Z+i3E4e3tRISeOfOTBf0RN8EBuySm2bH1xhY3bVuIRjkvtP
nmszZD42I8+mkeuZ1V6t5/nymCTp/7soPrJ7bgX9RyF5hjqG3N8I1tp0sRUBpkr2WR8TBLIOwlp9
IcHP4xCwt/VwpnJaJCBaulVTgBhNFO/3eSGiLz3AcgtS2XOHWEz/n2/Hcfi+TzhygVPjkawX1zFR
5j9Wi1+ewGeGY4qT2tPUh12hL/cT8D6rs1zdmu8LI8++xwhjgGciiujj5xTnwQJpioc5e4ROnCTV
WmIKIPb3w4iYH/qmwvbVfCoFfQ7Xz9eQDSSBZJqMjL0wo4Xdrah2I5pEdPTRs9TrNW+4ueFkiExU
tcRqRww0EqQfNW8X3VjFv2G2AzBz11a4cg9ghjfj9/TOCdOQLv8AaT+/gucbczjj14pQ8T6OwbuS
kNp03ZVwMZBvHmnFdhQN75XdJPCuydUT7pIeiR1ys40Teemw/qXxWlqIPJqDly35A6+OM9p5AW+K
p8WuBoJH0/GnoFAbpNcQl8WWC/IYUAunbzJQ1/zxK2YXpuMZqXOg7sHNYRCoCLL9MaDQtsX+VfYQ
gCclnmoLagE2zs8Qesn0cynN0ABbf8AQPuJXpA2QuZ3mY8VwySZO4gE/9NczAMy+2TwdJtJzfvDr
lBquOShnmfduLnaJ8rZsWmnfUpiNHp8u4Ll4bKODxaIFI2PMsywLIxWXpNfCOW1U1F8OKfZ6HtiS
cRv5dnevtf7VZ6wZUOTOkyDQJTNOY0ryoHpUget45P3R1mSpzO8/VtHQxv5kJX3FAvx3XVjUoHJf
8TbN5jrzRjf5XFDK9kIP9cnNiWtb+Ncl157jAPXPLwXlvLV2b+MSII1rPPE9VYjqjFk2yaG3oCAf
qXeFv2uWc1UlMmZDZb1+e5idyTgoR1vwzT1r1+iLcqLMjpx0VMqxwBHDQisFhNrPbaZNekc91oae
wdZLg5PQUsFZ8Whf8r7MZKJvDXzgbK9Q3F9SPEo92Uxb6RB9mvjulAmYHgmEzJWfhAS328zIiqS7
3jj+J1PgTtW9kFhuZ9h8t6UHBWpIAsDwt8rBTeHtUZj95+m1JiioTWsj5GFHQNhARxeWdgUtYULk
l4zvyn3JsYnG0AHQpyEWzgxvTSVm/jAklKyEreR/4H7YiUbnAgKiu9FZQsFZiAEogXJPzlr4lX9J
lgpx98F4qvvdYa7py4ljsvXbN7U5j9yfA2uT0FXQOp93x08gULeh+s19tFcK1RQM2Qxym1HxlNDx
ZD1xKqGMpYu9zOBvIB0fUm6UaSj9A9xc8uH5BlKMLvRTHAF/NLaMagkzURRX0pugJ49zId302jBY
pgqVYihHCxKL+mp7zO0nZpPKPsoAYTP33JQuNXmty/439sHHnKC4avD5vOo8bf32zfOBdjWQ6+FO
45picK3bTHynQ2H2CjOhfA26MlHSA3qtFU2CP97nBecVLOXKD04Z7s6VavOuFs8gb+uXd/0oBc6L
ojXYuby1kTZIpzV+niPHjuFmqACtHGjxYgSNTH2jP+or8tHlIQec0EIn0ehKko6ZamFvKRKN39sG
l31IW231ip3UZzCyGNidQ9JRapBtPzRYiDnlmRSE44e1so1thVTRLiFHD7vrQd7HbIx9/VcvDa5j
kNid+nB9tn8gDePxI2ai4a9voQ87Dwc+wE4Dz8yvYacDuCK2ltDillBH7ig4z6LVPyRri8+EIEPQ
g/EkPKPm6CZESuedeMZq1TQkBYlKTKegbTxw8DAC7vL/3+O7rjZF05segANkmOCOEOjU1PIPoUkG
//u7uOfFJ7+75Tbrylxa8Mkw43gcv+WVIOqbNZQvKdHB7IMlM3eEY6VTObm5MqoPuGpM+9HvfM2t
yZ60dx+ONWs+YbilvzRo69st88RaVmTezGlFJriuLk/y8F61K3U5puqkUvUM0qNuUSKgWTnWhMRt
NeBXWV8ih6dw9Nxnqttrfs8rD4xTfYFCAqXYTNT3o4aZlH37JW9PuYnM83Cn+W8NEaSk4gadNlJE
mzarcuxV0TojOG9i7FfMpOdu/txIoyW94hq0plFsUbDPQC5ZtBFIyDdCfd2WV5Bs4AJ8dLB5mu4G
6n5WV6hSz3JJ6xgQqk/lbhR/jw717n0zkZA2aQYLaqGD1fu799DTMGkwcsG77TpghodXnTSOgOyY
WECB+XhtCJGegvqhNY5pcmC0aM5bFKhlv7RGWbSCiUyfBZiUENl1SEH0McRuYTnoAFbGXi0wRUEG
6lUzdcO+ghf6xThoJ/r5Phw4vcRL3ZSy2gBnLjxQ/bndj69ZlyrGbNdUETMsLCvJOh+e9LwYq/OZ
o9tX/0LAoUPcXOAd4x0xavYDNf8VGlL4LOqfPLo+hcLP10p+Qfn54rbhcMeGMylb/k6VfVYNdZcV
I90fotoIOQokvzFYj4vgtfQdn3S/wk8sBsi8DIs1gPEJEtwYIVyIq7ZH3KQjXTYRNB66nY/uAmgD
Q9fCC3Rl9AGY6yQeTe9WYRjEJ31Ae5YMaIG7Ldd1Be3MLc2eHIlOsto6kBSN/WUOW+xigmB/Khsy
uiGoKcYHoMRAEylJF4AozYSOteWN3hHYwd8AC+V3r2ElPcqak6BB5byUKkKufH+G8d3WEuzJJ+v9
T7TQSufSiW+AeSQVXQNmdEX3E1K/4g2DNLWDeRVEWP9cTcZZedNy8Gx/sMfOjhGRZjNl+cENWs0R
GKMMkULNjHlGd3XtnCsWF4FNn7cxdSsCeaXVBYoQdhEPgkLDznRL4HEg33Relx8gOYmrN+NEMHj4
HqUhd3wXqrw7Rlu4wlBTNcTecaTguezF6nTVvJYPs1H/vSPrH5VaciJSnIXUH+KTOk4ttwj2kLN9
wyPoSEz7hs4HSumo2bLoT1StnBvjBmsvOL/aOd1dxNvP9NaWGOUoteJLwxxkTCD7SrhR1ZJE/YjL
MqdoPBszoB3AL6bbRaql2nvrJyA+qlkdJQaJT+tNdF3uLmVI2Nnc0zOQboYdfL2zzDKjA/ECxMKK
nJm4Q3QJ0yfx5y0rHuLy0V4kSvtm/HDcIPEZswFE0IBPqmWWSIieuBn7G3QICYQASkMYrPHsRChi
g/ozu2Zk19pnQyIWjJqbsbBclTrj8iMXM1Aagqv4/GVDX6PfTVoCPWQWW/bJlM5Oq6aTmI9iepVy
BnLJdegBm9AzhjDfYklDnC8jTlRyNaf191lpjt27m0LxSqZIU9YZaR8mkCUQmwrVF5Vph42W3jr5
WvBsXJH6NdEKanoWYnobb9kRZd3U3YuuMoVpXCSzPdhGwaipdx89f/kt96GdAa62fOA5snkmJGmz
4bbDDbe/biJxAwM7L7vvU0LiMSEvs69fo8rqvmqhEX5Xg7FIPQGeY/EkWnsnZfAwzMFalW5fsWMK
tESOkn8KL1IW47CREu81pG+XLrQ6VKa6EVjNTiJeMd3MFlqHOuaCajZePi3omQ+w0R4H8KnWKF6w
J47S5f94MPHb9JBWcHoUr+hCt9GAXVO14ElM+Zt3ykEHRaFrdUSN39LdCz75upFLYzqkvdFzbakP
myDIBwuoCKQ1SpggxtEzblOYVRPG9SVlVv74EiBlW3b27EzQhEJzf4TL6+drX1MTU5QO7n5qUksz
v5+biEhenmr2BDACbEJNcQZmtHS2BhgwIF+Q4LcAHPGPfwn3or/MLN1xVy4xBG9jzUNFUPqySfNV
EzU4UfMmo8pYiFKwejj4pgjVZCYrHGTX7+IZvCWbE7p94DDyQQSL+2AWaq0sZAkgmBHiB5CNcrDB
UUoEgfhV5jx4Sa5KhJ3B2m/FJllsWH7lemxqebE2Md7qtCVHGHbdbG6ct9a4dhQOO5oFw8CPdV3h
QyKCOdFwo/0HvIOnCHwBMtISfKwn+xJU6ZR3bfcU9M5ercecg47L3qyJcOSAYvrcXyLFij9FS9WX
bwkHP+inJsraxA1FQQ6VZa1Fq+kMEJ68KWXd7JZ3PQRWYe9GBM3oSy14+Ub96mdQIzmHG3ajzr1A
f9WzIjOQD71o95ufeIQpqYE8mvztLB+4mKTwS1Sx+h0q+PS87RddhbdnJne0PG0v+snP6kpFn5/5
quUGhlgFyMrt+cIZZ6L66AG+ZG4bVeZdtRCnxWCZx8uSTfOtiJ063ZkFFEzwQnKcPxNMUbWYt1FF
N1lIP1N6FeQx5IgnWWnA5NZHzzzXK3tMi9a4QMX40hxXB503HIOcMJrjMJMQwmSRgztjG6oLzBVT
UQnhMu1V3ODY1TEBwo6oU45v9qXCDZgW6RZaB2XyKWTVF6LptniOnobkb2SKN/RUIshLVQ7yKbAv
Yb13g7gj8ceglsYgxgZeU5Y7HO1Y6z5K0i5nluC9ljTv6qVs0me/1+6wPH/21TxVE62B/QYZG9uk
JYWvaQhnSIMUaxTsd+FVpaTCtx6i9aGE72tKGy+liJkkRmLjanyvsQ2GHBDv7+yQXYr6gARuWMua
Rz/x2v3qM86RFeRm2fbXUVGFo4rjJ7YH9hN8PFFBC5+m6QAwH51Ay/+Ci5CnhGlUw9Hbh87nClQ3
Z6DunO/nx6B5duM7TEdKME5nT7/DyNgCEnRieQ43yqoTvh2URU4NkaOVvVT9WsnczxEWP86Kr4Ki
2JZUAlFMxPmve7QlefnAXAYP3JPy0/IqptXKC8MijGVewufqYxz0dBaFUCV0V4jL+IXGPcDwr5+Z
Px4fPucxJO3OXQtfyAHo7/i4xnQl+X+dXiobzucLlONRRVlkklFUXUl8E/6/8PhVs41I9tsSCJM7
aGcikWZbUshg5V76Eb9dXO25UEFtvoVqwQZKKoeBSnwf/eE1vlgj4Cyo4azfw8+vwj2SC0gbv5Pe
ZFrPYKhoQgWHvYVyYaqUNdn3/HHCj2xTSvizRRyfPMJ9yqMKBm8n0nVpBweUHipkcUc3TB5IGs0z
9882vCoLs7jxqHZ4oZeEqEqENybOiUhH1pVa0uy1Zf7kNZGj2heRp7DekKsw+8sFOgevFf/rhSGu
hp73GXlAGhVYg3I12SIHzQeJa75HyAQEelfHXbKuQ8uFyBmc6JEDHu7IFA3KSzGYQfL6CLXWmTGo
P0LfkMBXkeuBHAskEh5mL2MqnxqTp0/NpWVvOoYLUNdiVbDGKtP7eSbzl17okchjC5XC5lEq+xa1
fpc1TG8WW426TAKjqVw8UaHvRVYn3Y4Dj3zct8kYMs4xQXKuudgx9V8lEVULtXgPy4Eg1PUVZAtt
hIDCqPkdohnD2+i7EzFS/pmZ4SvbQ0OlPPJQHJ9Yfg8u5wx6sxf/9ObC/WSz5ZGINoroHPr2NGeu
jC4xxf+k+UEU70/GECyViQAJdif50AVFLWciKIm6XMJPU54Rh4su7sDZnBnF4v78p0vbxHdTtPY7
gjguVAPloewjlS9tBiXcqp7Ht8yfc7VWZ5jQ7U2VvElo7wcnXh2JOPOr30wq25m+o69lUi6Cp7A9
VtqgPY6nJpnmPZcgv4aqr3k/3JrS34YJH771FWGzP1oyb3ipmu3h63NnDVxs966JdhZzn10ln2EL
+tAYtoFxcltvl4QEBCT5xC63e0UzF0GWBGChf3DMTXeqKXKzzgohSwqvedHnNvoJNj8FVTnhV5Zf
SqtOCFzLi44fDtyWu7Glas9zKoY0hdV61rioGNd7N2FkqQlDTrtkyiTpC2WAjcBlIIqnSZC31QC2
8tdTz1SErw81Y43i0CB/FOldTwRHkFbxfeCiZkKA59tiwwU+JAzH3V4U/c/im1KkvTPUQmTEn/O/
yjIE5ktgp/lgLbgp9v1SN8U7iiqe62ebMwrtqE8g4xVNAxc1eABGtulHUi07MPxsr4TeKXzW9P6k
+uKn59QtapiyQpAv2L/Ao0EH8YnRTjN6MohSsje/LJoVZ9+V7pju7vcz8ALXY/euyc/FE7Xd2F8H
h0ZzXUQyAArbcgyul8ehB3wjBaUfwW+abILRJG8+daeHDf0UGQXYw04BUaqGjvUGge8GeWyjZWzU
yoPqMtKPWI3BEpNN7Pj//V5dwdDCqm1dzZ0+D+OrMUfnT67nxFwxXC2uloIcBmB0PvartqLfCoDD
XCQkw3YMjiOV5A2n+8gV4QUJ0EMas11eM3yOLD83tew2oHvzAsBWh/TuH4chg9xNGnsPzGyV5al2
qQypoGAYQQjkFE5keT2d60FjVfajzInqQyhRYZ9v3Rz7lmCybAayq/YTTdpKb4K7Hc+HhHyR1SsV
V01SLyls9/G2aWeL+7vL8Ri53Uk4SrsVxmXFg6sGlhr9/AKpYWKJJBrVx6jCF3PdaJ/6al2dz37I
WT/CaSFABHfGLiLEb02WC/oRB2qOewgMohcx2rCjddLZmH0Tw5Fx9Y7juuYHHfFhefXdTi4DJHRR
nuQBG9pmpiYFB0L8JzIHB8ohIfiRwv0mNyeFLnzKsvfBJzEWav4/xZ0whom4eao3HY3g/LJ2lcC/
8ZyQ1Lm7OaECuod3eDHkDxlGuE3knofI7FGpzdKrc6EYESg9ALGrAzU5limg3lBtrvXHP1QEjqt7
cVX+OwoRejlPuTJyZOF3hHu5awMruo8kbLcSEDZ/m/YTGe9SA1SYQeaZiVCWCMMMZ4aPmvA9Eojm
fj8l5hcQeI5CgkKwpuMVDkUzvnPevzpfhipndZdsEo9XpZUoAMq8F6k+qbPMlhDVTF1fCjKdPiSy
lq4vJX0IXAMEeRn/prOAIV5sPVVSzmk1BFVjDKT+PxImkt5RO3n5W77KAlL2uhSHgyi/Cr8NEtLA
qA4D5ft2CwcKHQZfQS0RVmpKxDGqscjhkWy8K4fPtlJ6hnswmEWPCIYiswyvwOsETPLV3r2Dko07
WwQ3yUR/GvNcLbWpZCt6eaHWd7jNvR1YizqmKRMAAL9bshorvBklP3R6mzj3hOuU3UjmwVyxFRQV
0wmNCxfz9Y3WNcqA1XzdmkupvI6pMADZ52aYt60fAkhlZ1U2lnH8lHuvfCIqwXR6h3jCzjlhag27
t08Frw2HPLr8xl2qdb1/Zm9XNhQuj2xTqJWVx60E/g2P1wcshgVYzY8EKH0jptOaVy8uMLvp7UO7
n+29aW4b8+b2TwZneYWcTJRL1rMrqHs47DpaeidLztmaJHZQrxlkO89YtSCheeyRsAWMOipNQM+0
PSaooLsQSaIgnSkx50JjZ7I/BUuOlJeyI0xbU1Qw5XTOdwbt2QefKRuuluEookfoPEE6dlaMrS1J
Qh6MYmoHuHA+Fqe+FCdJvLkzBxKNspKXuEPgl9s+eIS3gd4Bx0twwad7bENftfQiEb2N255RSywU
oDqcEZPQk3TBYgBLiwYkLZs9hSjiDFUzeSO6tk4sM2j7gbXiQZvzw1DyBSFxAgej0dd/LVoLy9Da
gPAiXzakggg+W12flIk8zM6I8XoCWQslYzaXtdlCSGUYKB6afBFjl1pUv6cr6KBzq1CP+K4BUonc
1epqnigOk7XSPxki7REWIF6+nT55kaZmuU0CMYdoL0Hzaz3ZqNiv1m97naZ1kP8TYhcXEn4VAWXo
Ol4Skfzr2hr1KOtl+PJsWhMxp7zPAnC9m2XdXqf5BNBA4MfUb6JydSiHFhiDh5ZnOhtElQeYK0KG
ESDGBajmraxuJ27vum00VO+ClM2KLmX37MfE5vGrzrwO5OiIxq8Uai2P3/sKJS7j8QVU20vPp/C9
EJOA/xQFOCIn7oMY56DaOI2wV80XbXDBHp70Gv75tkHozQgxQ/fGZKg/K7Rt8K+qhK2AcS6XCOiR
cEYqKWdSrJpAYGD2wbHtNOzIxP3ScJU7YkIMbB19ZqE1Jir2S3jPvpoVPG2pIYaZ5gYnrC284tYO
Ol9Ig2RvDg18WbVTER7/6f6LBuQvfbdQlBDf0W9djWuHzX+rsfk+ianzjblRZPlmjCajDeWymU01
JUIW+hlKdwRVMljAUZuOTNNYOtnQjG4/gkvJrHOOpk/0p5ixJ/6kaENt03klwNz7EVQFjaQk+QzU
FX7kwJgO5gCt7vinmHtyy1KreyUXy10sxCblF0WWXaLyY16RuW2rnhvcyEiaSk5COySRS8CZ9VfZ
j48L4Vaz69XQN3MryPlyDZxcusN/SAq4ns0ZyYiKYuFqNW7OEf/GVJjaW1Z5K44+nPBuk4f+iMYo
qyFE0+W9gLZ6KlJYB3vD2tDd+ch8VRk+CONJcHBXJ68QeAC8jQFUy5Dq0b+kY4FaF9RbhmIT7vuB
XxgrjT9eS1Ui3ZOtX9k5yTI75El35xHeI5cCm85aglsxSf6iTgBueeJydIHSchV6OD1PGgCDn9b+
vLHE96doVlcK6YcZSTJqzUCJ6+1iqIvUqxfj2QPLREc4mji9wMYOj4KGfwH/jvrMfRnKjhz1TfP/
p2J1v4q3PQq8UwOqNXLfPAHa7HAlDyy6n49fhhu9qiqsiehvUbxQ6y+JtP4JaSQkaZNsvJXfbWOP
TZZ9MAahKFhl26WqQz5xzkkIgB9HAGlQIFriw4N7Ky4WK0qC2yoVGXjRPmkQ8ou7Hc0nZo64O0md
zBJ0f6bd3PVK2+4DpnWvn/UXD3sElcWt0rK3zYAsKc679XZprmrS65fNdOh5tNbLmGF5JBRGs9yN
+NX3Rk3/4tSDcHgpDY29R2ZKIkRP40aeR36L9+QtpaYY3FUApFzxRNlykHsUZijzjBNXI1KLmIG3
3NSMYINWHsrdL6Q4KxtPERHyYBjK2p4LEjfUX7V7/9/Pf7Acp7ClVMZV6f1J105++VCRpnzEaecT
EoML8M+gWt2MAQ9/j+IwAZVjfj9vG+r9773oYDXC2YmjI4OxuUNzEXiVLC2SoCiXR6EwyA2MTA2N
vuzkwjGiKnL/BTJLhNiDPB6PxJBrdCtGSb1OtCq3WrYRhZlJx4Xdo/JhLJi/2Pt6lid7rSsEafxV
BQw3ziJo9PbdHU7I3psIsdhTPbea8Cz32N2Kb8ebiM2qBcvSA8mtsMSKiSuP9NWkiod+BGt19oFl
5IbmLWleOUX7/134xzTVw3nYXGhghwsdQdV9fzryl5xGKUboJSB4VHmPpHuB4kVjtqzlRk7Dioiu
lxyxS/3Qr1FVUJnu7ATwbCkf9l6kSMWZ0i7bNsOIxD8kXbJua952SUq3acms9Wd1VgeXTzVYe2F1
izi+1sekWcCGlQKC3imVXCOMga9O2pzUD3NRWAjGVCXJSAFXr9J5o7dZo0WefuPVQMB1214QPw+1
urd3VxB58VNn2UnRzGkDg/kLL3DfoPM1fIWQivXgJeB0k1JOeMsa2B88fm/Prt7uaEBAhGlsN2UY
mJUDicKjd9TY541qOQCqXbGGvMEx1fgK/WRVa8BsTe/0eQUSEHtGl8cCWtek3WVwQSkbZcl5wAFx
5kQhzp1uTlynIYx6+yFt6ZZKsykNa/fjxLzbkxo15Kd/MRcZtmFRw9j9GPJ+/MVhoea23IeaS8sq
R/Kz2LWwdV/BIk35Zzulu3w5at7A7wbxDGPUgjeCZMl5/93VWhVqAdUmqKGBzm9EuELoQJ0rvt0t
0/BQ1KnldzLokuaIDLrKH2ij0jBfGQAlaMk3WBpCIwMlWJg4HB+d+S4VuUQoypqmDmsYuWTJibyR
N846/JXDz0p/uLFPAIA5u8d0K/ZsrPT5aZob9UNMiT1y6w1bbLqYW9/4seWPPQz84dZeOU4DARZJ
8RWccdI+RMqzeuDcVKxlawSzqm+uA39w6FY+yTbFYUHqOLlYs0uVD2j1mgfosfjSZmQyHE+1skuT
djR7BzQCJG6BoG9DAUxhE4Tli0vzRaGXsmX0FBrTiderMyjZPEXKc9PMLbawMzd9IiIEHtrk56O5
Y+pw4U8qwnXNzlnOKUVNtUot3vws4TKnqjox6Dt9Z+Z/2A3WRNb6qD2ys4Mf4MBZuDwZm76TExBC
E3b9odUxVnPyxLXXAeY4MWGjeDQuhE7+kINRLYS0orhpBMLrGA7dNDmOnjyscJ0OK3Quc/w3QoEh
++E30adi0rSGDpjzPwiidqG1odked1OPbNkmdi0chilm617aFvIwNflhDF81ZBtge1pVYj0HxxRW
da6hg6frkXYPaKB5BKKxqZW3WsjWPEumorOQvjuKKDrn0qCdRa67MdJLVC652TzKhXDAxAN8mLbA
nmvFpHVAizmdpokXYA04A+fupqUbU48aOex9qWZvs1vGqIwNU0NmGCjBS8B6+rlRb21CaUxuKfaY
UxNfOKKMkSqGgI5zcSZOONJDmrG1F3VPqmqp56AjW2w5viTqk3LrxktJ70SCDQ2j4yBvkk9pe9mt
nrKB9S9XW2G76WJ6d9mHCxpxyCWZAijStUAJ99N6l4iI8gvId/cS2x24uIEYRYKbd5FcoU4saCc+
xFY5J3a4b3gThX2CjXpYo+wFFWXbT8HeNfcmWT26exrR9nq7oIXunzozq1XP0C5/S7pwZPcsob6j
sb+LTsQGJPm73syOkaoJgyaFJxToLsf5VcAAy0ivYqIfu6QyI6DVl+H+97eb4QQSQ9aUxiyGTxnG
/0w2PaM5aRWG8Njar7sXFdBcS5Izncnv1P09McGCPT60oMQIRVkUomJpoQfhxNOHhFnMIExlNLHy
RZXA/xOeDdfC1po4hmtb8PvawWHz4njneQhh4VpbpE4g11FxME7X4xTWhpe0Fjcph9QRDeBw2WZ9
pa8iF1UA6HeuG5W4NMgQjiR0XVBC+t0b8++S/cooz7ekDELqxDrqmIiXZrhLK2NTHCW8KoLMe1DU
bfWkkZx4DkxcwF9QAUbOWWQ3NXSU5soqnc0PmGNCr/sAYR/G1qHK66d+KB7sCMxJB7J2584qoRXN
a7ikPI8OFne5axH6IohoEfilgUXxjw7SYmf2YuAcpxBE39ygm4ehdhyZxm9SimimatP/jQDpqdvY
V674nEShQW6iZqA/j23lRKHX10/pTSwbBRp6bUUL1MFbgufJ2YCOmsrZJrXVweMaiF6aS14e/GFU
CApcu81FtwRWAq1ITM+GPnH3Vt9tljpCKssxaEAuzTtpsF1XZn6B7yjpKVMgdtpQAqcJbROIolYE
u+PllT7+GaTA/gWzcfzqYawG9ZgyHOzhq0KAX27HhHN2rnMhPPyCHZMF3QiPUPrD5/v2DO1c6gTN
LQbsQDxWKr3Z62l6dt0kMAs7X8dxn9tDoax2jF7cR/G7m2TRdmg6bTu6Wg4+GWdAX8g+dgdxfIDJ
PtyaZ2O+LFjv69HT3HFJFEIVCNzfEIjm7iRz6LJFr3TL1GALeRAEeTGf+w74sIsfW8lQ9vQGTai3
gzDD56X0j6CuUmv5vkJKzx6FbGKcF1a1sFiOD5iPYdBy2ME8kre8ppMZUGIW0wjVxKzkLKi97zgm
mAfhu18Ts297wNswVkS8p0i0BhCGIPgebchWbV0sU1GCSDhc1kUXvbHCbAFJ/VNAKKkrIURuS37R
hzXQ5SR8tXjBYGeUlafDyj+awMxFyqAQsPfpZTdEsdJuhnLE7q37oeY4S0NbXtIqngHdXgybHHqp
1V0OoblUTmy2BMr/AzxM+KQiB3en5O8S/oTzOWy/zXFGnlFuJM4QmVRJoKA/8iTYuWQB2vPqSpdn
eCLfphDimRIW/MhXz6/lIeuDWicUNh59rdurkPPXZQlMcqmOsFYCAo2UrU0efZbGXK0A/O+RKb5s
FDsNCzv/zT7/qOs/HwPXfy6P6tE456BdjgHz/rG309aGndNDOmsC05LpylnzxpqO6FYk9pWH8sSM
xuUpTOodf6nVta/CP03Mv+4A0AfQuqr3zsVK+91YgpdIbNGJ/t6EBZMQ36al9cAK2Ie84sdIsiOh
angxEVj+NKLgd9vZTlu/IYXAn/ptPGDs2R+/ZIsFYLiri8q2uAoJcW+0tD3ffCxV+dxM0DzZD2Xk
NXPg9p9vCfNNSYPMZxdG1EQVc+W2LXteFE4gCEYwv94y0BfYhRV/y72V+NLZv/5WnibfprGyTxk2
zZ/M+d7KXTB+Ontm6sJrlWaU7JatzqAt7vxCD5gTtAzTMKAAv7AdWKC5bkzt9v+xVs89vjct8jWu
tSe/OHH6ilsd0qD9Jzv8VinDa9kgboDus24B0p+nUuwLRHKW2Ehx2pda7+r7pe1f6v1W2fBPGnOf
QU7OyvoVTaSEdGIgIKdpAbkgnr6TC2GHWm0AFd7uYradbMtVolt7Tc9gUkxCO00w5BGFKWO6x1xL
I7NRVlz5tmP8vNY7JUL92LpojE6NrpW6bM+f3XnUsftrkXqVoXVex839/RYVEJW7pdmn/vBSXxYb
s0TzAPReb++skbXHosVHc0O32C55b9kjGzHqNB9TnauLyenoCV0mRj+I89X8JZ1R7p7rj4Hm6Dp5
ijQPf3zKV1IIRrb8taJZ10I3miBT5M6l/z43AP4q7r18r8r/vRSMD44ahyAuEXYfgM4thyB9iMrI
WT7YzaKR5kkI9kzU7JkHgmtRlph/hCuSKGNk79UQQePCy+PBMLFBOSSErd+9RVWcWlvHkNOp7oXP
Lca8H+6WMzah4lhC93go1imuqIvrQqWiqayc68S8QMoSfWADoo9icWx9Z2105ApxADeZfqEH6fBM
USmJFvD7Itjz1ssK0RpVmqCtieC6f1TgseozvmE7Rnh7v96N1fxui1DIM+DbR6rhGS11zzHTojVB
aHq9ZSp9jzB1ul7+XpH56LHaN0++c6wagXTZZJmjOSmOOk4IyV5Hhv+CgQlp00+7ywsK2M6ynUUp
MFaiR/uMYtPxUrPzQt/QolKh3bl9H46rjjzF7JHX2ZxHiSO+Jv2jXnFXM4AI7F+B5p5u0ixwOd6V
ObJ3JvpKiWcBQ0FyS1soAu4BjED3Usb9V4FY0cZCYYq6X2kmFhVvJRZ+q/LG97UGcHhf+DA5zRZv
jiMU9KwFSBcsMnixZfm9H/VMTb7xwl5DOQnLOZjYvGu6vwzEPuw26ayryRfJnBhLwJ46C7qk+Y3m
KHN0dZzSMfcQl12P+ME7hhv2P8YA54XhxS+rn24SqaqzbQxbDtfpMqDeHCetoG3OrmH3QEs7itcu
QUuTtF1xf+KP4DV0NBCE2wnXGzRFntPR2RKNmq7AWWSrbj8d1Ioi3bptdyzmLPjV4I6jhUitNBCJ
Du+kLNYyhAAH8/rQtwSW9tM774LDngSE2iCqzESfOrwOqCwxjIGVko8L61XdMd2t1KMw2bIv5Yt4
8/4NYqGUUpsQbvxM5oQezTS6XCSx6J2pjEczSu5YzmaKe25eNPtl9Se3KsKK0to3JbmSGDd++9YI
CfoO/iU4hPjytkBVvB/fLzDwCV/jEOCX9kPNmXA3wVrZSWMtWvgzCx3E6NDvcGSSwxtQGcaiZlvP
GLI2d83gwCQJbHlBO4x3sWMoM/CYDMH0pVL3kLA4BbNP9ZQukpMWmn2NNb8oAnO6OcJD0Un/gopn
oca9lpiv1BDPexunHa1fKRCPZMRG6xtbZmjfOzmJLwbynJTn6jYiRT5iO1+HpyKQ2NmqHWahWNrE
dLW08mEJHQToGJ/dD+pgXkTiKDNhtBG8UsUDW1XpoQfxbIeWzFl0CZbz6nBj5V7PcJwLdZiHIOjz
58Vt/6N9qfp1smM/lf2pbSHwRE8ha7NdQ3nHZrbZ7qnvhnZfdj/Hjga70qShFFi1abrJ3bNz734t
RwcmSz/cRpiSmJIEhwvXO2Hs+2ZzG95fymQLBx5xKJVNVwKV/Rw6rW14rDSYxLK54DspqMly1vJy
Lrnqo24uRdezqz200M3v45cFYvfyIBeigFLnytu1w9OTnU0y0nOBRjR6HS5cBWMokDhB2hJ+61Xi
8/5cxNJ038luWHQvonoAu2qzhSl0xvRQ0ZYOe+mjPpOaAxP0adjv9tTu2L+Xd4DWtGe0otcG67KT
a+30vRQ2U+WHXEW/Gi3R3mvLs1ZKsbHgsGTeeklYaxjKTd3CEUUPJL6i+mfcnApbEKsHXhoUEpHF
uiPPxo8jVKm8V5P8BmWDA8+YRcMh9OYJ4pGQnNU5KlSh9i4hoZPiWPGHCNJIDVUfXzYiz6Zb/DZ6
Xv8CPw8x+F+kzdlFPpsQP+33vgnzkr/gjphPdJD6zL+0NYPuxLEW0ArYK98KeHDY7Ycnf37XT3TR
mPnb0AUvra+3beDl0TxSuS0sZRcpxBLxe4rqAVBe0Sxx0QwB+l3yki0V4e+GLaH7rwzIzBFqVT19
Pk71p+POisRkONMecRsoAr+q3n01sm9m+mZL4p5ieNVbbJYLGseQKh6BFp/N9JWDPPTlyjfpJM0A
ihH+uaE5/GfADPoma6FvhmwTfPeisP0PTNVpblRghi5YTvkIH7kW4s9PncB3+R6paQy873cwi1GS
RroqBldzuGDWt3dxwbXwKUB/mIYsoiGUWo1/Kd8L38CfMc2baDissVjssfscJNnl+MA78ieTB4MG
K2Nj1hiAIe14uw9F/KVxj3tLvJx9Qv77JUrIbSbCghlYfMWNAlYCup0yQgvkcKcWuI64S8vxH7vp
jmdaIC0KD+ppjaV6zkoYJZFNgJcloFjccjOwWYHaR7lAqqqA4eiTFc9v1lLqkW1D9X5tV59u8yEL
w2gsEYy/dBZ/kFXHkJ4Gt9T8sxnaaSl/4njYeojW8LCFXV8u+55bmr/JxrfA5nfxnDM0r1FOoZUt
153WZsdR0dRlEuF97LD4njS04ut/4a8bHuT2CGuRuSoQF9f+5nnwh2vU03vBoWAN15PrrO+eqPD3
oZ0EaK/I6PYxyq8oFwt6+i3Fu6LaDliG+jLellp3+mtSUa8bePtG32YZwTaixjIsHGUArcl8e/SC
Jq57Dyi8cZNpPfBafdrQymMdgiZhFzrkF9BYD1ZAOuySemT/ybVXnDw9HMUZrJJd1XnZB35oGicM
cO69XGmkISAwzhpnKls4WeAq4Pyd9f7est3n/vf7kYD/eJ38j0hM1ep+OatY5uguA+zcPO8/lei6
t8Lbw9bDFEPdZB59tmRc3lr8WQbgtEUpgVuf51vdROzpVMh4ApgSl1DRujew4PgrXP7e68hVogEi
BiDq9QnEKQVL/1z7LhFVo+bDnj8WGwc4NGOdqLAnFP0dsupGWRxnELcYSbeJW8smWIWiQqeFbYno
rS+NWM+ULVzWzm60J2GcO2+E5USUivrpjfZfU+QYRv9cHhnq9tuWnbfR8B8R6TBCwMtBf3nfoyst
GuxXsPXXNQ3llXJyXbpg4N0CCmgoWml+raorEyKcEt2Ipdd/6uOB29nBT08wYxLjTsqDjX1aMlB7
Ie4ZKjhLruKjigpo/CrJq1ovYG8+NZCIbOucFI4HSMGxJlcz3SJI3zVsT/RGZONJe0cluTUsR5Pj
a4nJSgw+yqIwWXPxpDlxnAxXwdbBcPVComlTl8UHxDwdEq7cf0U5FqXAx3HYk7bAJGk+2sQPsFG/
fNv60CwXETuFl6HlRPqBLuVYAnJZqHuRQtcIzsqDVh7YL21C78YUdL1S+XGWDEBkWDMJVW5+ygVo
WAsEKW+d6tJB5IPCotYjt1jC+R4atL2/sfUcspALtLy2S/sJDsho2uEbywHHC8vQkuo9BGRr+eer
PsEvGCKnFO9QpycLCcvnFOVuvKzchGKYxyAKTty6HZ7HX/sP+wwaMpO3uzDXpRt0eSE7QyvlZzlr
DzK/I7HDmHjOE3KwOHqs7ePaqwIR4cyD/saY3PEqe+Owh1RqpFLdXdu/7m4tWrIGjXy4WAOsHise
XHQUfUUXu+HIHZM/oEJRr3rJdM/TR4spa2QS5JaJEtGM5ZTjhpSxC4vEOcTTZTJai4al1861K4Fc
dhxAJrRKok73igwA9R6Ju1WO7id7NTvIeLfycJuMZq4fYaKUDLbO5kjLKbisHnovwkABxOYCn26P
qNG+v6IzoDG5lggOVtAhi08wvvYx8yIlXh8Xrxbvk9VxBFe8R0sVxc+7NiECrW8NxK/4k/M0RC+z
i62oYCkLKY2H95sw1KIkCTZpRefZJ2lMec/8jBkBqgVPp1hWjiaof1582KnW4RKQ4aK+s5yd1VKD
/igyZ2joKUeQ2yy7i3mpnlF+Z6NCxxeqVRIL4fyup1LvexUun61BrcaSLOHvSw0T4M8WuvCW0C4Q
iE1COv5/spvBSjOmR0z1IIGU5u2KsWPUIOay+jfz++Gu3jB9evUj8Yo8zP/byinoe6v4uGg6y2C6
qVbip8htiVZENKXVSoSGqKaSjUbtjuIw/vtKeQc4rTGyUhHY9khGYuFpxvT6jT8DpONiPvVUWwjh
dsFHfmhT32A1yn/Yu9e+g9ekDmNihMAMBvFI1tY7wYJljsKx4UBAvuB3+HEOPHuiZr08d/d8TWSh
oWKLLyrqnEhV6LEsvOy+e7TTPWVu96NJ5glva9/VGmCogvRCjETWILkNz0vzXd8PJqXvkH8oOVwH
hWPdPUiE28Kd5Il4EfKQrDm1ImpeJgIMwKi+qGiH8NVewB80bll5IS357KvlM6uKmWvVknGg81Rf
tSAkuhTiU0WJeQpUbF7pi+jpP/ImBcBDXeBduKCzKhkZDNW+4h+VGblKafaDFjOpgC1BsV6//xXV
RfjjKDTnwmyQOWVBUybrDLymdlttKLsBcBNVPrXYuyuWNqDqVgvr1O+NgxZLNWYriKbk9fqIOi6Q
13Uq3JWwXJj9GhBGDoEMr9j1ftzSv5TPvfjxexT5bq0Igt+LzQZfUNmtnGAadGT0pACR+Xn9J90N
tNO5jrojDHZot/eq65xataLEiJcEeIIFOK4Ivrom6zwlxR7Ci0RfIjhtvw4BMZi1yTuMu/66GzRs
xik6GwQe7g2is+TKTXzmDinS+kk/inDJ3nZ2y3K3cj/A04Wl1s6RU5+ZovuwGK9SdQvhVz1FF/ds
ZlaOps+XS728s5BXmCvL19TrFtKd1NvfYvDyekjrEUJnoIrhaZsluV0+RtTHxNGk0+X68mi4tJpG
i1BZ+DlSIZxYUa2M4C1AzM6ap0KSsGLdquVcmjZ5qAWUXWQemIxcMTg+zc9/kWR5QHdS64QgJulh
S0r2CF1/TQHZlUUyO1K1CutZFUhadLwtr9QqCo70m+VyvH27J/SqnXtPUn9cBbDyd5xifo23C/Vz
hkXgQ8Dzz5STxOevz+29ZGyUykNHUxIQHMicUfokTIPJE6b2uLvF8DRgUnQYdorh2O/2ARqzRXX2
x0Aw4NmaXNGXoVZwGkV9UC2UpGQ66k/7sWgr/y+akc/1Ov0y5Lktgn4XetnHT+1X9tlU2ZpjVwwl
fJLEVObTCQXOln8Foe1eI9j77lvlN9QZC0bnJBygmxyMRxYTX74Nnme+ozDZhk758DABPtJrvcVP
QmTIb9BXMOFbrPDFmbRjN5pryYvndm2yhyZ2JOhuItMlG0yim/lKCEYAWAKwe/qFgojqJl/r71s2
6cihlg5qiO79dYFk4OZBnWif4GzR/GfHq7ftXU4VOSke1+vYO5xYGIMeo4Z43I7FVNSb6UXVAcoA
PHq1639wDbrhaZYttiOTx6WRNUK2sqDO1tmnCkBCpl/3YKjqlFCQXcCvHjudjXB48oiPdEjXa4Cr
Ns4sMZh7Q88KptzZ0PBttY++eyXgeORYeTPa2IeimtesuyAQoCGlcyaempbXusNigkakm1+W8+jd
EANgyKwH8yoB/ONKS0j0Re/01SuI9Jqup5VRSsnkX4sRklvg8sJWqFb8Q4A4ggrZklaDZsENqqBZ
UYn6zeIjFV4snigmf2ijztvSQQ4Hh2X916beV2VMc2tgep4LH++egiBNN1qzLt23BWcuI7F4S4Md
EjVi4yMXNqnpNhWyMUGu7a6jvC7hEAhLblXpnhQkoCyjWB3TAfAvlv8NhC0a6sX6VKT6ustoKPRv
hkTqL5pkRoUaHS1APg7R+7Owz30rCC1cEMwN/OLxKuQjBUqdGJb4GXietJcAzIwO4rHlJAVMHGDt
aBi0PRI5V9QZWwQUuXqPJ/441UNW3aNT3fZVlJpRTjfsTU0kgzhEI9zqR4lET7Dplq2Vl940ic2Z
m8BYB6P5CzJZ+zsjLFyE8qAzncMVCIplSEHOP7O7b263JMQ0qZ1rNY4MhM4izKSjsRDFdoG3RnnE
oj/T31sYpakEPUCnQg/m0Ewy50JWX3RQMhshmc2X0BAMNQsCHBLpJwph51NoHYBm15AMNgcoBDpZ
9yTUh23nsmziawfImK2J5WhpCXezGg/+hrM+gvMsAewFHyrDuWjjNaMRyH9Xh5ZbRgD50dSxqIKB
q3MhJeW8z7aQP3lvI46fkGlmQypbU0+dArAlu3BnnNDVEO+LxshXbGCTd6hJhSxBanhAMHVNdF+U
Cu6PreSeVrMuiRWVCE1kgH9HDNaL3bFK/QumabQ+k2LIsfptbFf8ZqmGj9rXAmCVogyQjRTtx3uH
MdLdqjBypxrqWxCF+ru0wTCoMF5L6yT+W8d+Ffj55hYhQEjolgS6imfdW04dvRylMFpSlpA3Zn1b
qjR1CEDo6dIRuUzNBnHo9mBmABFz9eyh04qGdX1NxwVxIPeuf1wS/E56ynsYb+952kK2FYjvWfG9
FLSXbV6ouC7DLZgjALPx/9XyaosqnaTBxlXsO2T0Nmg7JEbGG+5kcCisRM+vZb2AmHHWoX9ls34N
zE84DehvrH8qHY6sTS+6NFKr1C+YmH7M8oRdThE41ptxq26Sd5Qgk72fogu8RMM/hvcRFJNrIAfP
jLFlVFa+Ic8zpl3wM2Xzr0QMLG/GJazqdwudzuycLPT6Xwqxehm1mUimAKeg7yP+li2YpP5Mv5HY
JlZwWaVN/fsN6bKWTUuqb7Lw6iPmtMMQGe6SPGa3tCoya/tVDjYECutLJo3zEEMGLOWqeIJBLaN9
I/HzUqqcTMUsrguF4uTIf0HLFE9JciWTC3vJQQKsAob4kLgXBd50ixy/CB7Z1vbsQKZDssplgtQL
zR2ziG6nnjDs6fTZo4Aprl+OfCjBRwn3jXFs9VgDTX2qMBbMS/9J6SfAlJOtE6oJsXBNBLQAgzVk
wJVGC/d82TR1wZ2KBsY3w1sfM/O6yhdGlgrQyBPq1TCpnvAjLyNGBmFVOplHjWlr9jNKiCUfkURg
OfM3YXPJJRUUBwKNySeKInoe791psinsjLLTUpNtkaADxQQACPXZzPqRCHKuxWzBhTR4zLv6ucp8
SVbB9fL8PGrOItxLU8vNivcd+6KHgVQwgFOameBK6SAJTbut+RjRPpQkLzUtzT9MvyyunDcCt9Vn
swOMm1uotvLaJhE0piSDW/KTpICj8RcUGE0Fg26DcoVsELu5fQ0TWWIzKOCYkpjtqwS12JyPrIN+
bGuWUT4GWwc3ss4MuDZZKp3ust0PlsW5ygdbqRzWCiQJMmzxlMwADx/BozPdUAT+BeTsftn4UtrS
+g4GPh80cGHttUSLmxgAAaDd4TzQuh2L3z8PuwK2b0fhUW3/7YaPNTSAHYpf75lh/cfapX42Fsi/
vWNFR8ok9xeDwZioxzUQgN5hGRQM6oyS5elg7gAak0w4NV0TEzt7N21BERTTL1C9cYvmRScS7Jvr
NdKba4qfvnIRI0kJ79azPZ7n6hme+611bMRBU+MpmUcA5iRzxKnKrK/pm/q36Lo/LHFFpNxMwcOA
MIzsGaOaKJ/hDUBJbeougua4iboZ5ckXbK9Ph0wtFXrONs5V7SaR1leN3pkLWUsZ+/u8+8PYPdXn
mxSXb6Bxi9VNCv8kbhL6iVd6fjwtLqt11LK2MuDkS6Nl4PxCZWeOgBE28ZWBDKLcySgbJKa9vDDt
e5q84hwvf55aJU087qCKUecvTeDf7B1dc5ve9JoKdtNL16086G9L058VkapyXLoMJvzw/BJkLuxz
Wt7nShnvT2orijnmzQDflSmJEiqnCDcwXTdPpE7cF2Ier6iPSCDyNQev+r6HmoGDrhKEM8B9Sk23
F5XfS9xKevdn1sJ8uwutbIy8K9asmrb132ag08uJNYXwgobLo8Uro3OFXsPyJ4QzzRk1JEB5vN+V
E1trlsCzdDtagQdWMYRoyubXjB1Q+1WHwGESi56jEunTIgr9lPQOimY+um+RcIKZsk8bCB/0SXE8
dvDLXtE+/4vvoAZSsrgfiQMJNQCo4HRLM5UoAnR+jsaKBNIjFDYJ17pCaXgoMNnEOwqk9kb7fgiP
M3owG4415Zs1mxM8+lPcu+4kw8kOiDWTO3M45lPqTbjTwIrtmn6fXtO3z0cQwu+/2xdAyQS2Ni8y
qfjyOESI5GhF/XZClsUAIMh6RAZJ6Zf9DUa3g4FFBYPdFt0UvLRkYikTyUdSSLN0uykZ9ZVeJeYa
UNgubSz7guqcR2jciI7/2mpnVxZD5WhLxosb6VyfVd2XdWBnndB57b5W7859LjFCSH/hFeoAgOo1
wgDC2dCSc+PULLRKKwkFBB0aPl86iC071TKEOEt4jSCyd66D2dRsX/XjpU1gY8Kzm45B1zY6Zrvg
9y5mVmnOfjTvPHqwYskDKmFz4LhsS6KLFtcIrFvU45TiFGWldI0to0JxW/OwdHfmNaYwkTtiDnlQ
Ag4ey+oCt3mTTTgWF4mDS+c83bZACoMRV4y7MwxQrvesWQAW4Zof7UzgA9HC8HNr48QZHjcCFQB6
ZpobjwL8eMctxrYA1QMBa4egaHSq8Dvnv6WY3nLJLEmS/rRz+dRwnNnMwA1bKQ20OsM89Ow7jfpF
gv39fJHDTLU+KfEp7QZTPWtS73C95zqT2a2tah1aoEqzAqyHNVDnry1S+ZC0EpFToGAdlYsGDc9Y
awLw+JPPqTlU8yGAeK4hCet0ALnEahvP2Ce4mwhjG6Ndd2azoWeFIPdh0o5rsDewa68fw6JOSQxL
TUrShfm1JWQ8P0I3tRPAhP1AtNNgj6Vz9oABjEaR9nsvbCOGYePVRQEyhRr0/Zct9RqJoTgskIMq
XLPOl/P8lQu3ADt1NiBZyOty/27Yn0IR0L1pbwQjL1P4oczqTGn1M2Wp8D3YOukVwVd1oBNZvghp
pW7BvSNaBwOR7F0+FRRSjCsMjbUwPz59qWbpws6j/HRVpZakFp0GFiN2ucCuE/ttlKmafHevF8DG
gOaGX5LbEQuQLqPiAayINfrUiPo5VeOBgZjyYPwFhdi/xspZkgaQE38KLErVZGMOZUMoEXjESg3b
6IgxEu7/+ikmSCasZ2QYa5kdMSaMH15SaGGws2LxLMpCk+Z2ijHVoaC6hrQYsGcODOLlKDieR0PE
2unstkwM3p3zoX4icq9J+Et1QzVKR0ckxgj1x6eibMVIN2vd3XbbRQtZi4lYQTH0iwtqVVKVf89n
pqTz8aVK2nbQbfZhZXVcm4ewCZjLDzcegfr7tut1Vr2+6sDtLTc4z6w3wqEWG48n64EtjbF9mQYO
jQUakmsz6LHlshf54wMrjHzOxAbP1HTd9JHlVvrIS6t24RanFEXvPA0xbstqKuE6V1jUywwAagck
ljABBejExxWOmKVkmFKV/sTtDPKHY7WDEMQlai4mlM+ZoXuAIsfpAQKWKxschMK4e72JtOxqIsW3
EAkxAHLCDuG9UnNw5WkAXVPcg0oK8YvzDhuAH8CCSlRRZ4ZXaT8yt3/BYLrUYL56f8GHUWp2hCPL
nehBr3D50z9b3FERLh+XDsyUxizQAZa4KhE98+l9bJbRnVw1SP4ymrvixT3FavdVjkyNbTxTuRp6
u4Ui8gikC2Mzg9WMlsWFMXPU1ppK0BcqAHuqFnEb+ViLLJmYohfpv+wAq3g6iQAxjaxd7AXbUxeO
WJ4NuHTdKhFoeIV59g8eD4BFHH5TpYEQonkSFh4oquIeg4jiIS7bcHTpzXSncR7xGQlIjVvISV83
PpW5bu7CxzF9sxVVxt3kNvPo4N4jwLdvdaXrKK56LXbEddEdaDFBi+Zl/RsBWEWaqF8Jgxx2KwF3
d1xK807UWsiN6dkxthGXC7kK8tpmsNITdueoa0dGA43tgKKgUKkABFHRpFUpg8awKAhGi4ZjWqUK
Qr6wkTh2eMDjBDjLzosQXskrnnFCocHt+m3f/9BJhkaNiM64ySwUEe34cLv+pwtS5qTMBg4FCFFv
bZ9fjrCutW7RM5a/RxT2uPGIIf72slrFchZsbFp6HaMzSvlRYQtAYUjwyZAm23pinObccIXNIpki
jXRX94YNJvLw63l3zkB0uOBAqw6Ke+UUBpedEv9gtuomr+0chf81P9pL4JGHgfwOxFeAZLscASaC
ZRouAGiamWTloVzO3JX3Q8OVD2FyOEIAow98J7XvrMUg922s5DJ2xkfZe1rJ0sB/yI46/bg2QEGp
IDQ3J6y0rs03Z4PxQRkzJHVPKYm1drFEVbks8A53f+KHNM8khz3DmHfsOlU6pH3o5tOeemyrehJ5
rJtrYeUTMhEIwJZTlgAf5iDzT2fGBEwyRmCYtlC1U01WJbGKYZT07LSm3rxsGrn3pPet3cuOk56e
CB3x2xCkDrc9HKJuUBwxVsNM8bBdEhzgQZaiAbxF+maJCxgEj3qMm4gVxf2ztZeWit6kbODFz4xP
Ih0E2VL/05SYarJEE8UVv8gZWLob60mqA1Ivezt8PrzpTaV0Xdj6O4pvUoIPP4tWjXeddrcKM+hQ
mR6U1+EEqBFP+uzcnXOXqYXJCR53Pt3KHAizL6wv4Q3jheB5scBkdOvf3izSVOTCT/hP2rkwiPYb
F7UKHkBd6pppbJ7qz30sll2B7FRB9FEMZ7heeAam+iO8P1PkhcMS3b7JCvKg5RnP9tllRO98N734
4rFziEtQWRdevIE1XQR1JDtYJ/WWbmKIDmF5+2svY0XIM6hHbnkXiuBMBrsp5+C8+pQzibDdjxT5
ADlOmtdX81oSGIgNmxFZVdGaLaWoulJPR6Q71nOgPSehxoKaQ1yhRW3/qSvVaIoUOsIseH4vKNMZ
KF3ZiLtUgtj0QW/BaZjfixrmagEqJmMDSc5P8YrQbQkz/b2UrZbh2EZOm3lmv0RO452WHRfHDaAG
WME8nqt2rFN+eZZsfmTVx7zr5gWIKDfRukF1YFfKxb2efIL4IwnTCqA9TspQt9PF0wKLdo+S8jGD
igDSpSOr97EUD5EuJ2G6fJxfyqYOkCTBB3U/9fB0Xu+1ARf5GvPCpp4P5oTl0YcY3eiWmSWMYjME
wcX442TBHNRNU1uaFJB7AqNcxKFZAhVLRasAxea0fgtbStlLqmeTDQc7M9J3n9gVTQf6SrypfkRQ
CVfqFFs6WqrJa9anf1ZW0GJTaEOv/2S+66LMmSHfuSnsA6HqaAoiZWo0EjNnR7I9Quc5d/qQchc1
kG2VkIJVosIzoFHTzSuGWX+N2WAqzF8CYuA681KsFa6CgTfTBbPPUFdUTjiczh/dqlH2Le8LB03k
GK3sfpY5ZagI1viWKZDMztihsCVgDcBNx7CMhoa+zqd+UKaeJDmfi9ge+BxQMiw0TNlG3YgY40D8
NjrRV0PhZqFXlI909PnBawGLajfw50yEWMuZTI9dTonYYQ1cggyGEbtQ/4ohzgadcQw0x/Ss1z+C
OK8iE6/PZGy80P1UnYApMLGbrF/hivoiFJcooNaGTzy+sToQhplxaEt5ED3hBuJgZ/MEoQMV6yJR
r6W4lrhFARDJvrmhmYS3PviF5W7I0+iCZHZ1yrlmNFhxezqgjWtnh6tRl4JjwxmgYy9Y4uyzwkFd
9kZIJkK18rPCeuX2/vA3eB9IlP9UIBpUovIktCExtAITC2t9UjGj9fO20VcyRkCXsP5Sy37FFU+r
ayuqTCFztiQVPfrPFKhLBUizn8otpDqQEIrm0iL9mzhrqjxyrorr+ohUEjuqaFf8WNoM85hH6ZIR
8pSjtkuZjMtak4Bp4Oy6YXfonZN6sk4ql8o4c0ix/vSMYHt6H6ckKkDXtFRiaUHtg3ILvPvGy4Fk
Venoy77UUK1VoJB8z0Vutd5kMscqk9KFfZ8A+upfdpW1jbZLX8VSyT02z/HNG5APxeZIvYW+53Kl
d9+y6RnzbSVSJgydUJo7eLv6zB53SMNXwJkGa22EjyMz6AoR/OBAFCLlciARyXf1s0bhjKADQeWa
nnZOb+5Me4aIHzNToRltpyHTtG0h19wnM7fDNthv2vKsxokQhlDxISrovzqjuRk3k4GJsuKmbZCt
M4u0zQYMjYEmPmKvDR1Yr+hfGOD/AsclufyMHe2B0XXTlaJY0VrZ0lLO4PqocPR8rNa/xHZnMFYf
jetGQDubtzvwTWolHrh1WP1IV9EFhiSNEWLCE9MJWaKp2PdlB9kMUFpgWckZdPEHklZ0uwMvYHaD
8LsYm1/S1339HEfC0IiVB7CXlN4m6nlWCzd2WW95tIxWhedg10+d4K4eOBABYh6eTvsg2BYEfmgy
81780l0CUsubaRInHEjQGCS+TWHQjdPST1RA0MC6xYa4qn3DB5JFeHw6CtcAQ6z283BQUxeNmX9Q
L2xq1V/mIIB+ECCBPtl1TRRljNwM/f8u0LDEe/N79xgL8Kw1jItWw6l5y1Ra8x4dTfZVNdU1VtPF
p08CD0rp9sHGE0J2mUF6lZw0HFplRhlJ8c1oHeDIfigR64Dn5QNli7ScDJAvMcYjgd0fY15jzMHW
ikdkqJ8ga6UKUiCw/ylRA/StDCFA3qzdpOF9nBkpMTg225vwRrHiHzi2fm4DHwhfdIYLAI+gYkZX
hLxyzNlpXQWEvqKF6jbG6GUu8hkb+S3lCq6qcgN4KQc4lNwhINVoyCM2cZzz8UuV5XuDSiowxIrR
oc9ld50wkFZFLSJMXZl1b4u0CWSPt34kXhB/CO2k1Y8h4Ff1fvVN0wWx0IcbjvkYttOd7Brm8hE2
zLGtSHaFpRVzKW10pl2cIMETNxP3Bb5HRCnsbOFsTVVb7g2//SK9yKSwahpuWI7yCw7FnpRdvDuz
uEGtmmyPAHDcWdvlGNG0alHqoNeLhlP2OAmroq4HJFSbxTBFNImS3d7QQ3e4CCVVpACljskQVIZH
vuj1ex0KCPTkp2V28IVsfTkXU6bIMlsGhjIe/rXHMt+pv2lQtA1QNNYytFoKavDBPb0peoV8o0J2
t980QtgqTi/MsfOW8/1+gWTJ0cC00/zl9/T0e9m2/sxRI/Pa0EENDk4SuQSmJwHAga9Vsl3s3lfN
VTdgdKdJH76fJNCrl4hRrxGschl8+zNTPvLaBTlCYo9LUhlMtK/a4Ek6WNGtw0SAdJGH+AkYvrJe
ERGuml5aDeVq7UybayM/qgrG9/bzxVRED0j9n9cJVDaQPbbn3nfQKseANpk/BI+E3WjAGdjAoyaa
DJ/eerGsP3YPLe1KA9GHGJEh9eDa/llf0B92lOGsv5iE9zAacK5pDp3bHU8mWeMx3gZo5YTurAxr
WI/64Oqw9obvrxQoOpmuKj+WF16stQ/wNDJA8Xk/P0w4gxfF4/6G77w9OyYVN/GEbLSpZe0NI4j+
Ul523CfGW8DC8DcaYi8Wh17yWf62oiHHJ+vl8zRDnYgz/JDCqAEsVxceiy7LkbM66vG6HJboAsUO
IDMoQyANPdQAbSfOPjh+DYQYDk79L0mXHeOldAsGqgHS6IXyXKOdji2W+JSbwytZCC1++KWFi56o
4VqUCCgIxEU0qXpLXX3ZLjEhQd0WaClpdLjojkAsKYuwzbc8JJIDgGaPKbNTA3/Q8TSqfRAdM7xR
4Tp3WB2X8dTWHidYnAsSdhA4QHzJkMU0Votny+dgUYtpOfGmjISbz9Vd7SW8xfBKYxU1xCR8xb7E
SDkAlaPpft5DFwd1Dr6SBuOOHoyJc0QmsQ3q8zPMchdhvirQe/I/ONLmiTVmJzulOcCUovR6LxVa
onwu/umQdj1iSN09euaatnZfzfghGSKCwiZXMrQayrNDN1CdoOwNDUdlKAKcH9DqofWMH449BmmI
43c2tAxDhvcsZu2nXk8uUZO0Z9iEREsxNeE9JVD7iHiA+zx/ZCKeuns4waFKgYkh83q/GGpn0YtJ
99waKSbW15N9Av62KKfwCGporgpYFQTpdaDvK1qCW2gP3pLUKZQHw9LcV7mRPIHe0y6kPDoQ5LX0
s9qISdtj38JGSpk1774K1YuNvCgYArxVmN2EL4Q3Fyfwc1frHY6+3CDG7lOAozmlpvjHLMoszTDi
zZhakVEmv1R3jZp1owKHZ+9zgCPel/seme1yJ6QKrLdHAIoERdUqSNycX9M2oCvaovS2ZeylGtSs
vTQ8We3bazYSyUf75tUjk2g5VzPun94CXUocyLoV5Y9WBv+JO0ToyCxa0YvsU49BTA+8yzGNOOcB
zMI9xemT/iFhsHnzD07ZdL8yGA7M9u7T59jQshw9Pz+yM4oHwBbTaB0r0lGpzTW51/3KzAc4VeIf
WuZuf9/ckx9dNGA0qcGDuN0ViFT05YtE8ks/XjjJXNKanTs4LbrD2JrsRRkNCom+tQVHgXtteX9N
XFFiDvaFA3oZcWtqee2h05u/NcPSRa1ILJdDWHbGVXpORmxwdpd3TPUVRkluPZuIMizU9tNfyDeH
DjPBCickjqWpB+3zx/J0EmctyU/H45TO/5dGYKG7AGLL2YQl2dfUWy26ZSZA3AN2BPUGyFYqK7G4
30O59Yh4maQ4KUImDfa31yIp5wwNd37ToZ8POKLp/IDmaLP0TNE0KT9Ga1PRxNkSxIJXPuhF4FLl
EDKDEbC3pIOJjRcnElEFWnP9sR/DrMCTuLdi9Ud0aP1REWQEZkmTIxpPBVgN7vD/pVVpulIuaVfZ
U9VFjRJzRVvZ5Abb+00wofCRoKyrkcnvV4g+fNmJAas9B88wPpMkzGAtUCiRjjT05N2NG+urCrP3
L143v0Vyojk6CZPtvxOx7pztHuzd5YDYqLZH38o0X4pdVGQiv9UpQjuEyEsxJWx7VGRSSclTFmli
URW2e7zoEKBfVlXcWdI5WEQWcpwLMdLMcVB/eRRtSnGII7ApLaXckliPAa8O1qDGYnVcgJDe9K16
uwnAj5sJ4CgQa+Qf+zo1X0lv2vg6L8DA2pawLjrg9Zg/F1b2a1oNKl73kbokCGR7oFRKQyggngnZ
oOYK4wwZBskQ4glE0BFR2Zmi2fSB9Y4IwIIcVHhMdz7LrvH9YbDcjexjJaQ2VBChq5D8qbVXYT5F
549i+V3OWsi/CLRalbOR4CRIiBkbvzeNOZJgPNtyp0za9F7prTtEJ42RNK4ieYSlkySiMgmkcWWb
OuNRoGDA8B81NddIRSnRLEMp3ubIDRmavjzWWZcAyKsG1u/3UjCROHYxYeaBQ63IdF9XhqHIJ1GM
22ptuqGslmq0aE8Lgibq/rGPhv7pPTEY7rG4Vyzp2qnyCjy0MIuZspH3QqM25vnWEbH2ayrkdfRK
/Wqj6ClZQFBOJU4BLWIfxfMbtcf5jrmtZRbtP58uMW7DV7TF0RhAArrUnDSsU/1+tcziM09Jjyxu
JAtdztzrRqk/U37TzmqHbmUtDQ59BCCT7jag0vFzaHO35lCb6uDAzFcuE9x0klOHazzbzCT0Hz60
YtMUB23sKsUJOuqs5wXIb5XKOy878uEpoN6lO5CVHG9oJRhkJvaJfms2mbhLHRN/tpRFKqMUTUwI
Cr+vRy46Qiu5C/POcxL4EmHbBY/Czdr6LdLpn2hwVafiJRsyaNPdtjlamFScZGwVyfcqJ4MrjVlD
vIJUwVfpbZsc8ACODxDsPff0lu+6/eImRbjlMR/ZOVnWZp2SBp1thbD8XEvdQAKHyrOfKmfWRQ/m
CB/3aKOvRFtEeBysLOyZJNkakbAYO8KyO2CtJx21Ghopk1zSczaomQX+TUdqbvf69hqg1wUZ9R5n
tJYRSI+0NeUE43ipAUz3bfRKmotBATz9eexbRv4rhMABhvVluIm9xlj2iGromrzFm2fdL3NgENwd
3DyvUmletVMBlMv1Q57TJaY8G+tsOo8BKy9g3shLbl3yvmLxvkqP5wTOsr4Rj/rnX8APCS5Uscy6
/z2MOVjAs/H1pllsP2yc3sQ9Wa929uXtLznGm46V6hIAp/CDRNEsaaQC1G0bL+ihi9sI2gHFckMJ
AxtQDXcGAVhk+iaAJ4wX9/KLeQUbf/iIxJbNwfzmzmV3ek+0RHSd8x6dPxx31udmQONWfIis7ZEm
0eeJHC86aDkcU5ZBbnuqrXy5vxSl56B3FXv/mlQBbIbn4DwjtDdkr+kilFt7K6Cm0FNO0w8twQ3G
Pne0xKivlNVQFWV4i8XEEPmKkxH90Pg5yAZNKGCYnmkTirEnIcGtYtLnY0vA5PidoOmsqV5OmJ0e
EhyHnvgrBVXFcuEE3EpgXxs0a3JgsepMm2dbjiRAVvRqbqFXYIrzJM3n03EqfYub/jw6daUpfU1F
x+4GNEGVi6OyYrWylezSYJQoGVIKImNaklSEW/wtMAGwWCm5SRh4ww1u6kzd1rRVAUUt4IbvCFIk
UCGhzNBu8v2ksGSw6BDYzwUg7wKqRn11YUQinQxLBWZoJurE5Uc1zPH02AEIalWwrjSAxRY9WC0+
x2DUd0NPVWWV98Rys5KpLPsaljz1btJnJDBb8Y3FL8wOtliK4A6me4wsaEmaKWPAyc0QKEV/Q3K5
DBmyQYNaCvR+fmo7RCjf+BFpa5rl5o/qpjffKE478IGoRO6rdVWy1qCGe3LZHTKDIgI9ua40kmx2
IIovTkt1rSEhXtA9HCeziJVivUVosU5TjnvLdP5E2SzPCJ1UpvJXTjnCto9s/t+DJV3nJl8GfPfX
Ln8tmayZmW4dAfNWaI8NzigcnuC6Mvn9NeATLby1/wfvQWsORs1If7JqyYJGZOrLKdFBd1xdIwmz
SC+vcyr+ZEUTkiRxfu1HdK9S30VatBBh7Sfq7K3u9RiW1IUVkEFC8aO1ArkIsNI5DgyjRgLQpQVI
GZ0Rujv1LrsWlONmJDzoWhOTBLS5p2jWCHz0OdvGb+xgpwJmF+bJ/KwMoeZ/FVoCNODfSosJ/rqR
wtai9CGmR3m5v35knDZk3DtpMUkgZ6s7UEbWIu+UDX3QoTaWDZIllfx4pgt6oz3IMEI+/GhFuC62
0ViRNcZmJf2mTD6sI0W4frfItrmX9F2rcldeBy1ihhO7Xg65lkYSla5LRQ1ccnJciVLeMJF91nue
ATQrWSvWSt17VXoP54eINXC/Jw73H6mcstzPjDI0ET44D4Sk58qHyZZVNDDlnVu/kFW/24CVkigj
Z9ZGHlyt2QJ2rvX8JP6VC56imI0EJ7Sk48O5LeCxdNkkGYjtuznyiJaqnyhyx/DG5Upkhx0I4u/q
4m5Dvb2X5LN/WvNrCT/9qWI+20gREVfYabc4Y+G5MrnRhQWOvyOm95P9Il9WMCoRxHNjNovKHuZc
scSzhURv1a3fKpj/2REqv0Qhy/Ui7Q8LWHCr60nZqSFqmxiXAVpM/3lDZ+lFeI3zcna/v8B7XlQK
NR7CcFpBMVzyori7RtklA4MOYzpKT3Qb/hLlnt10W/4O0ubthsQFnUQKUI6vf6bHPZmIPcycCShj
micrUjJ//8v8y4MhP3abbXd5zW09vK+x6NazyBOe2i0rvE6sp2z+NNhL8ueo33qvcdyhORcf0GUm
m4y3Gl7tcnfTfwN+BZn8oEduCc4VmsotJyj50eLuaqAwPwCtv5lyQ4xTnZb/kWzLO+u3Oaoo62nt
hIvCpqUxNyME6B5Q9RsSveYLSEtqwgOfQmrc8yCiXjVwIdsQ97uIdgWR2c8gWzvU8b5sq5dZNKp4
BkSGFk/PaAtPaFiZxJQxJvpVJ4EluLiw9KEavnYpdDJF5Zvw8GB9bYG6l8YqlfMAiGNcehrLh5z2
I0ecdKrkh3l+pYSdzIIbMOOn7dKY28RedNUMONI9VamFcLi522GLZSlbyScqjKm0nxVjQtpXpK97
It+suofwGdf2lwo0NJdVvh8+u/SThhsQwdTWFkYtTYSp/NpDyD/07RYe9f1ixQHaBJuwees0Ke1R
IrEdro3Lx5p/f3d9GkRg5Qz2SgolykhuBtRg+lmlbXLtQzHvag97PB2zpDLp89oQp0PDAGKgpUdn
VisX1YuB6dxH2JYq5ywLb1L6cNeKiitgK+09goEuaJZNXqPf5CXe06IYZ8Y3XSUz+NY91rnz+5GK
4+lLgmWAIn79UaREmhzMxR6hU+PAJsFzDWiJCaHroVNxoTD4wo56bYWF+nMY6EQH4ukw+HIsl12G
jp1BGuzIWZ61iDSIEGcdsXPyXgpF4izhZzQ69cVm9gD1LBzgSU+86L8w+GXS85pTPHoOrd8c5xrK
oaN9HACkJU+29Ecl9x+FS4WGC7KBN/arkSTEl9PmJ8CEv0GY9PGAlCikVcd6rFZLZ3A7fH8jh1V4
DZis/WW0M0QNXyC80QciyFaNZ8Zv/LE7ebd8VlEYJ1LGJoFmzGew5iN4vdl2ffrdu0fVQDF8QTnN
yk9CfNL7+eu3rZKG8Vt3gLk2x+fkhhOkdisvxWOiUTW4fFUxmdgbfK2ZJsiDLUIu1oWfEJC5aOk4
vm4gV9w8kavHsWpjtcupAtG3sATwycblTFM+TYitN6LvuUUR05oUmrjZor4T2L4aM/vR/zAvieol
GOGnsHEu+e1Z6IOXw24Xq1chZHHlQpDcoTL1fopnWYmRxcUHtufq477QnnyMw8VNIsdn/+hM9fof
7yIOMuaVznPdjr9MTW4N+vmUBrF7SeqnifSOyw4NM5wfNxDoKiZeJw8CDGKUD1VvqkQXPDNP64TD
/uNfbSeObSVWOw0mk1LEfl4MXlhu2xz0/cgJF7r88p1cOtjpoV4kctVTxiTgMlz6/4eC6p0niTBT
gpcYfQAy6s9WEfbGNWJwpaC6elP/kS8KSX91hXrXKBVbIx6pEbrX6a8bwBEtoDNW7KVspAjvpHCZ
X3w1TZDo9CueSyfQ0Mo2iVzEQyvPVwRyBRGfWV0MSkX+ziMgZliWevjaL+3hFUDUqQCYTNmVr+4O
vIPIXcwQakx16pVxyQpAeZgubfEiZOMxZXTUhSQyhxMBU88sQKkKi9QVh3AQxmm5WamGZpdgScRx
ySYQZiEtryIGezKmaw291kz8J4Wym43zeGVNhzt1mMjSxSWKOFD5g7QyuttAY/a+UDljEL3kY/r9
mUddIm/95ZeFdlW2d1bUj9od2G8/Yt7Y53BMctCID/iVVq5rvMtb3r96gA57+tlT2RVRR3JAIb6M
PMd8lCO0zosAYzdwdc+wDEHBBE2lVQIdlDekFBtevnYAYKKe4w5wPGwFz/NJVsjvoQfqBIREfADB
fitrCIRRl+oE2GJ0+Rjv1xwolik/Xg4dt6z/Xorx6Qv7fn8stvIQYOHt1ZNYOikP8oslyOMQyQY5
jmjos7hd1J52tblFLNkshMmgnm7EC+kFsiBjUHw+YmBbL+RGo3gIoBfgXxnFCVfi3Atkhsut+5Tg
Njz5tul5xFpXmBYfeD61YO+PFykV0Dcrio+Try4QEsX/MBY1jYYTdv2ndab3Anff/1JsMNT9YUp7
fjxeH1+odUWD32+1yRtFKRodSC6YTIbidrUiv9bcP0jIopIjAA8ON4LAB+ivGAG8zh6RirxG6bzd
K+QUuMo5GHQGnvhhBBLnvsy/LqPVRDfLX2Pi3F65V17Jx4FnimO5bEVRugkU7dR3o6oRzXzgEJ5k
g3ZHnzs6rc+wToVSyJwNSRuZL+ff3SvRjdP3XVG4/fn8gVLIad9r75hyK6W6umvvvZMeAras6sfu
HZIIAtd9PXjVYvXnjBMZR5kTIAr7Gp/dR64TJRktbKE1K3yrrmy+4PPoOhphq+P5ZlYg2gjVFiEB
ylj6Nn8zXuhTbPDNxxeVLljJgpsaxZ/UheJXksDoLosWmb4aq7u7Gn8JbWNo72jfe1yze60eIb1d
24Pur5Ih9paC8lngEh2mNJeai65xvSHMad809sUUUIhBjIes+PZ1usctIlnwXGY941OjrIrBdh4F
qG4k8EopYhMGxAP1n1JxFSqCOSeok2Ubfo5p0WjkHhlL5nE6PNvo1Mn8klL/Q5ghycno6iHSiRMT
GbLilJLd6EvQg3K4a3re++fUKTAjIb00+mXUFZEZYe6Wye6jCS07pdoiYvEG/aRgnZvoGpvgDMw1
O3ozYDUNBmlsSvP/CewjX50V2cG47adfe+9lPvHJS+yvCalsvvkKE1JZqai3nzbt44MTSramfRAF
4lwG8bVLMrn2HVKP1oK+pMtsUrMP6LNMlcPYf0hjGNJE2YBPLovB1eKv5Ukrm6kqRqysVLQOwKdf
KFOy4A1ynhtoahgzk01ZXVVRiTKk1SeOqLpl8MAjMRUYhX/uiynYd/S8eD6HFJef8zDPGQJ5ifhR
AqSjpSAnqm2iLIBijb0KbgIVmPaSk/8H1YKPdRcwpXFrOGjgcuv71WWxrld0r+zvYwX27x/wJmyl
IHIbh8JrPp6MvrayO5mNg+sKByovlR7Fo/I/yK4iWXZVz6mJqKEvZBeyNB4nIoUvaFKpa2k00Itx
Rizj/09fgaxNYyeCSToP8yIUKypvPYKvSJ2G6TzFTLkaTtOJSwI6vJV0NTA7Vd/eD34jtCIVqPwS
ZLJjUWQhQcOySFiESH4yzGYETCbDsjj1Y7l2nWajkqv3BTlCjIAYkaTfB9kBvMu5rKc0TCOZRNJY
OXZ+OENWlSwKKnc6TPKlNgDiBWTsY337oiDiUFllNwhFRU1iHxm6YDAThoz8uR8w59nGkAF9fE0h
iwUbKURTxXqA0Ghr3topBQJQPq/2gT+BNDkPe8cRq1QPO62Beb5Rglbvq6WDgoUKXbunw0fb1XHS
DKTZj13MJOJfgFVulKVi0JGS3g5qy6AYObjJBGfvQdwWubGq6vBrppJwN+c1KHwN/yl7xVfS7s3q
O465QTt+GkIbFMvEZboEaVMUuSHoAs5Er4xAFeQQp7lkckNKqRGhaPyVrg2YKrf1XrszqU03Likj
hgpJ6DyuhhRbnz5BOe8srnSMR9t/7iA1+cThimVizDNIKJbHj+vPulvrICSQLsptvjFjc079+Bxn
okuofxSqSegZpc7+1LTV+lmufaRwjGBod2gc9WsklgpoXZ5A7HxJGhpE8SdJPOw2CEu925q+JkPo
EXGIUjKYziUrRe7JaiMYvWOJDoabK2nA+4Gw8rfNhgImJtneFdBrhemDZ7VKfbowq//UsrB1Y6ZC
P6d9HLng0QmoOH+LW8NY1tRVAffDxQ5Mww4El8KMh1TzblbDB6ibG4aSFfEsw9P+F3uLN6MEZlky
LU+GVBRTnNx7oBoZB5zo+A6c8OHzRwKVInCivumrHaJRuryOiQoAEyFoBgfjtaaT2eJvdmXX97gP
jtt1gXNlCxl7lUGXetFBmqE1+vnbO7GixlLODcMjSmsxmGR/54swto7DJuAtzZpl07pIvkIP4db2
mIn4ORexg2tNccKi5KFYKQ3z5hR5l4jRRRigZFDBfquRfxd6goQBkKVR9PT1uxIfH+4CO9dWXg6x
EuS6Urv708guGAHfnruZciTUII5wkF7MqVPiBaL6qyDZ7goqCbD8ReauvSxFFDJkNZINi0KnmF4c
y0NdT3uaZjrF0N58bzYXZkMbomll3XpsEfJVzUfbiv6cwWhNCTkDCO8PMx8hJd6xDJU+U6fN37v/
3mfqLm/1xF/0B24cqRWukYZSRBSZxhrVAS6C0hVVyv3sB3AxQ4ZXNxihPZ+1KALpcGxxCtbl86/e
SnljGAxafsHlpct1PgVrmjRAqWn3FWdmZuYl7KPk97kJpgZcDxYdV1CCm6v+FTnkrO5TxN1og4QS
cQlZssl7In+B3Xj/FCY7qA/VGBjho78EJiEt7etRHJzMEF5NPYRrePpwv2lUbpDHfzGAFPlD8Rjr
HXUT454ESsOdIUhKCnFPKbCbdiYmoqmzcZj5HpIDLONcoCg2PDSKOkwEEtfdQAratTzBHquVZRFm
I3jIVE9DjUDie1GNhpxT+5HPwUN0GbMBSL2wNqPN/3bKNS0xbojLC7qLnHOAG4YmkUFA6O/qPoEi
amIncUW5scviZ77LJBwlTPfJoxsA8FtZ+NUWjEdj0uqhxt2M06kzEWOYxQtXQWdqQaU6z7C6QKCZ
dRV1fUnWvznP85xIAniB+30LtLa00MSO/GRnAcjKgvWG9mEBmsLoKZL6NxTxzIU+eCmfoNfbpE3T
aFk9oB31XGEXy4MlXkHGKZ3hTW060XYrUJlmrRkB4l4sXwyFxHlwjBWjLICPIqb+4sKuINAyQBer
GpPFIYtEh9bKqM8nbGIr7uKeQVL7yI7gvkuV88RrvnvdWT3/HwkqNqN66qdqTC+Sxez7CznlTHhM
HlFUfRadUsSrzpumgUTVTOi6VvQWo9V7Q0Ii2pICl1Y9B6Qc7Vmk4tuDkXRoNgjiyP0Pcf9e1T4F
PKu4mwYdyg0kjqyjazLUgMTOobjpyAVuByeZ2H9OA+cvLg7UwmWSsH2dGUYOdSi+ObQiSRmwTE7r
UYr643yttKZ+eMs5/wSol1qaGbsK9c6X41uahfnt83Yoq3mmAjhm4KDZ2eygIcNnNKMjy5i0qWWv
XI3NVIZQ4og1DuAfCrjxCdI4EmwfpN+xmWRh+kUNJVM1uUeeIyzkye5YRCaY6KPu1DozdiBJDrad
xPxIVfM5FKoqHqYxSEtitoHB38hWustapi9kBLMJczjOles92UPcDPxbOFgBSO9lb6rmNo+a2gaw
bN/RZIPENCyIi4lkyf5ywW3z64JY4y/cb8t4SPGZQWd9OtFyZI0lpJx6JcsurZpOSkon+jfBFzF1
EaLCjE0RNaJ3X8xRLhOFuvkiVZm2dJdfta3jWItuFKeHrKlTeMRUCyytt+ieRzy7O/dTOtBazp96
7u02EfVKj39cSr6C5yrEqFhcHFApd6BNMfK/JqYOb/5fhtiYBM0AwXR+5JZP9AqOEilVKAGP5HDR
wH1xHCJwD1JSS39QCZ+d22KGIijp31CHCXjJx8sKw7z6K30jnDa00b6nukRLmWmkbka6E0GFaeY9
wB4Lc/jpEVUGhlu3RtmD6fLfPtMoAq5GnWa2UaSzcgZR/fDY99qRgg22wHOoV13UeLJlsTQI27ly
dgosdTZ+5XptOiEqB0yZpaXtIhmRM96o7ZGvXdvhRq5DSQXPIAVt3FzhhLrqtEN5yBvPwhxZMdTg
xeIM9PwI5Zu7QGw5uEYa3F9zlOaGZR5bFE0EmGFERrorHd8nzwuP4acdepNbuDn8WYLHJMsWT83a
nUpLMRosVKxXXsWUtW6qZXUUr5uvT6cguH54G7ej0/nBeVXn50MuWNJ6pi/tCGemXb+cDnW06ryJ
Xnx3vcfOrhIuAX9L6KcN+a3xSBBNRRK+KkYMWzM7QamlQo9sZoQhxyk2QYNh7fsdNW8ZKz3wT/tq
kCeWncKF1Gql6hVtvuYJ1D6o/L+BTWiw5O4uNK7GGtjXabiLl3LQody1Li69VflUCso/lCxymyjI
IRVNFGpFrDeCdpVXW0VtNrWPtAF+y2tVe1KwjQRHPZbQvqL0/XUrAyoloGiFZFq0oEQhe+p63I3G
4qMHrZcoDGAmrNP1yznXsbH5L5tsB7IK+kRxj8IyfuYqj/DoTV4R37hezEFuqEurZc9JFHBfnRSG
XwS+4C58+zpSVCJdICuIP+Y8zYpqyNB2uXRnVtSG2qGO2dpr+zFZEH98A61Pp7ttwj0yq+IpuI2p
JRSL0VrxnkrPxSnciDP3Kc8Ehpz1p5W5IzpmjYJjr79OeFSdKkndB6IDJjUrgkRpuYCWt8cBCCvB
BhZo/RqI6lbZQ7Mh3PQWeNC5ckt1N6MOWdk7rncIEu3NMDnV8rV46wkO1oYImxmaU1IKmufScP0e
mS6Th0fonp219du3Q7O3UZahnRDdYLcxq86entCdTRHEQGruBqhvEdnExvQYYN+buVpTGdSVaCWG
FRb0xvXcuWESie6GK/SDQoznl/ion9Hu64PxQ3RcM2tf3JJo9jUWFFqURDH/+vPFfjOTfraAoRIQ
ZsSl6SJpttDTpALg5oA+5nQTGvAi/tCfti75as2vXn6kqBRtJMM+AFA5ASdxg7r57UkAGwwZ+A4A
nmS2rtf645EKUlhecPLo5kIAyoEFeE+ZI75wqKRP3AHkHaFbqPDNruerGIq7flG+XAx2+csOIPpq
zVxJDcje8S7sqKY5M8+E6SyJvFBP9/2Ldy/BZ5ohvbrOeqqu4om94JxgG2MYSa0gBSdAJX9QXHC4
FFv0WtNSi9/LhYBxOr3yxPFkZKk+wk0a4ObVSYEyEnR8O15yQsjBQyjSFbyPdcTrPCZXhaMs/bmN
5/qAI2lXw2kN4iKLkmiUNVewzNRvZwEWtM4aN52ZLt0uVL26s69uiksYB5Ag7HwL/lVs5aYyYOXN
9WU0qxw45jPOoTP2RRvZKb9NocAupiZJkfazl3z9Fz2taS535c9gPAoLe0W9D5Yy9KxLC86lF+pa
j7Uwewqw3yazhbPlVz9bmfLXfUN1PV+my2Pfp0E+rM7h46ItCVmJVWZBs9Pu5zY976ZTkaZVoHII
63lxh6kHrcGQ7uRD6D1+VSJa1sMsOKgtoPxbcqLpZID1RJM5/iO+eR+8jMW7nMnT30Ot10xsaEQd
Gtw7k+w8UEkf+Sovr9mXeFZX35QoQViWMKgZQ8v0S0U3fljPcG/w3PaAmEXR7Y9gGlWgWO3VxopL
kK89UMUNy4xOx3sIYpEIuFwuw8RGrGDPNRWkDeqN/PmVstii8A97jYqzvyBgeK1mXRsjevhutRyM
znh0QtSAxoH+QcPsds5mBcRAyGHoAvu174NjjWO83e/ojo5NNFLUmApMBUfzmOdxyKJDK65b8XBk
65KRPaou2E6FYnlCsbbmkDahaf1jOxPwa2XP/8B/1qQLt5iRpfGrc41w+7R5k1kBmK8go3g/Geow
x7DGef4fcwY3XJXxvsxnSsbJhoc5v4MwmWTdzftEBIdm263T0TsJM1LzBBvoOdC9ITanQqZIS9uB
8oHu2gAdZheK+TBgmQ46ZsvEtMmjIbRORPeT2NtZVjrubh/gK/3xcWiEDnrUUJcMwJi6tpjvz5oQ
Pq36PvQfjVlhIyxcNGReIPkZ0VOwVa8zqKFEg/NzDrFBqjA1DYzNdx3AN4wdn5hu7WsroR/TJeue
gypcHPI8LgTO6SwcexJHCo9eu2ia9Lu4y20FQ/qB2/eZblbpl1uUH/PkgdgOrShOf8NwgxFN9I+u
R7ZNL0SRc9QaTOn/3kll0yEypquGc4j71SMSiW4Gy0+MoZoKbEs1Dptz+G7HGwjEDpHuut4sOJDr
UYmRbZC/bv4oiLxwaSCfRDy92OiuVC5mfPPtaYTpvyXsQPI1sJRd/6geg/x3ttWSJ4Wm4p32Korx
HkL6s5sp4OSQmD9jZUvVzbqh801TiPQGLdkH3Oz3spHugvsMq9Ij4vPnLJTeT6bjs5xlZvRdrzlM
gvRiyxV0MdXo4sZkq+gzZNwFxiaEpDnvDUW3n3VE+y+YSdi5sds16l61mmMNXgOEpwDyu4DkYbLT
NCeIOi6I/EoQRKV1xGNUAeLIyGSzAPbdvmAKqf1lfNLh/PwjAcXbveN1WhS6p65C+ouQbcLHsz1c
55voHki4BJUaF+BHUnCpfcrwE353wa36OrdbSM6fgl5GiJHTPwX0RTZFPC49chRnRqdfQXnGSeqe
IqyqEHM8aVu7+XLcHTXpM2TV6v/GYNdWBQ5ozkjVV511yilBKJgV9O83DoPSMC8MYV5qQThCPwpK
obBhPrKlJJTSeHFqrYoCh+MjS9eucHl0Yr3i/lk7VDzOc6rI6Jk17tShntGI4E3Y4y+um8gybuzX
jPp6WzJ3TzocT8XPXKW3KzCujU83rdMT3soInkXrjNxH/mUkAkgdGN7V/ctXvXiGcn0FFWWCwf/d
TUzzhQX7CX4qUgJjdX8KkpQcU31+6uDCANmoTXrwQ7hQt06+JYV7XxxraIwV7Jl14MxbZ3sCqYRX
8Uju/tQdEmGtOI8/iiEHqEZZGhrLwstOWNrRPNTpqX78Zw3vU+WHZd5SkaPlJs3gUtIlTPOdjUNZ
QxA3hY60032mAKPLOtvQjg6XJHLZa9LfJqet2lXrvgZYaAnolN7G9BrNP7xS99ljilXzHU+Kajbr
h5DbXBKT13EhlbihdD2k55eH0sqRmIDVFSv6lU0NHg90KhshWKL+GRxrkNyaRJMudJ91bQWtAPFU
3KpM/S4f+6hts2282RjfOaV8H4XAc/49UG40ogalaOSSNzpB0oomC5dzG6xPp71UnQX8H/+fwvxO
stjwHoGuIRPuLSW2vADSRsx9QDel9Wnh7rxjBTmMAMliULl1WMNq3fdC+KWG7w78JywsdUOOl9ls
Gou6zYuJn3dVlxT9U+s9w5izMLbPFEfgo3CUUdHl8q2xM3axEkbzUpsJC3n+uwURLAZINyHaJHH2
z3JZ9uHthlGHpR3+6TB41yD6Kg6HBppx/rCZ+T+i6Z1tc/ScUmpf7khsoD/LovP4jiMttwc+tAGA
XiqWqKtBx1yp9sq/KBqqOStF0SySZ9bFBfvoGiCZ1ai/xzas+Mb5m7MWpUkRvRwz3eULEnIUasoB
wi6Of5ruo3BTmj4gg+yrhuZ3SNSLGD4fRVthlmBqCDr4f+rq0rwgCNWjZDNhRWrsMydAPLfaRcgO
vSRErgmd6b1tijFGADqR7l8i6yFHSTLkunB0ClloGlHxyCCtio+3f5BcIU8ecb6fuJf0y587/nkg
uiPq+/DCcgU3yyMYNJdRwP+fPG+6uK7hV231XfYO5T24k4KGzfTEWNucrEhzMDfJvWNoCwOAmo0m
cDEW6yHnDrRvBkUXkR89UhZQIH8Z2uigE9bgnqOCe6i2AFRwAKDQplojQgkXopc7p6QCCxPL229a
xgvMrYsghY5NhwpKfCqNZB110fkaGZBY+7/fDYFvMCjRiwmV8Z+soaCw1JyUi6WnOMvFU+imKsCa
EWXDsfvaKvtO9Pr3ST4db0T+af9HVjRPsPv2O+trHsxcEKfwxjHq4KzKgAqyaUMQojNsFO0Twz9T
ITlITVJxK4JzEbuPeCa5dVy5/zRIoOW4UxCFc/Ld7gp0DUIfnLiyhbnZfzF2iPMmp5cq7iPvYH0+
s64zrAP9inQleDou7/OykpiC6r3upSthWhd1nVY6QCQioaDP/2DXI8vhKK7IVzn+//84/s3NR/bb
fp+N8cJSgJM2kQxf7VyBdlSwPbJfFPlKRVcqx2UKgHIlTXmpHuiQlQT/csT/ubBKD3pptWp1gczP
vus4ElpBQoZ1zmiQ+cHBeboLCyZTMKTkoGPGGTt4w5NF+sBNydSLhUVcBKf78+SbkL2yY9vSBOOD
liFKLWTKog1EoE4MQzDnCwKFsRve7lXTCRXAikp5hKTJQzROyXaQ3iTE5YnkngHJ31mCCp+zAsva
lG/btyFzdAgu5Z+kGS4/cijRcMd1tx8jPenGQAZyJUZ0XfDRrnGL9aJkSBr+wGfd96sQfDBWlRYW
z6iMr0QGYoBdBUD35nrLy78IzfRH8OrwHFWol1mRhCUqIpmWWk/0lRxkNGfhHdNStYXMsLl8g95t
FaNKRurUcFREoVSCRmkp5U165SJdR7fQ4sMWPy0RUYLK8WwDCgoGGCWIPTtuxz5qeWXV+vOpspVe
EFGjtD/DrDnP7KbX3a2Ilx27obwkLbIZn5nPGTkvrSvGPu8HykJzsCgShspRezlmcQd/myZTLWgQ
J8+IEYHsXk7L1WZGp4NX2vzW9aYunjgDwP0dRM/sRqeT0Y5GDJtC7bWXM3oOVjYgFfhq3NXum1AF
y5WqOwlqyGW2lLndDnki5CyPzii7euGDPkBDrRQ6OeFTPUpD1pzo5AkRVhXZBeCy7ejSegwxSnMm
qJTQXzJ6DOxeuNbqN1Xd1cnvleeN3giRTp6CxUk1WZx5Y5gRvWZgn5G0g5NHd44PkS4staoEUMGU
pNgS0tU7bgWsiQZABYhr4n/UmTmS9W4fGo0EfcPiarfhc61RbTPFda969BdGAcwRXTECea0LgCHt
o0qQRdjh1g7Bk358i6YnmD1h7OYQHqOe4aLWpvBevuulLj6h7FMkocbegqwmPJigNUv3n13SmgOD
tz8eNwLth4DYn0qrrIa15Ofy11Rf3JMTGR1eyMRmJzHvWrj7dlrZsaZOM/Fyh49cfilng9eiZf8H
uS6yaLtFqks5DiCBqiJ9JzCvg/nW++Z0x0B6/vLsguhcRtB58c7wCusYJ81btN/I9zL7vjXGRJbE
XpaYsF/jdlcJoeIcVIIBzyaOqUL2ZAwvffWoGXYLLeSjawJDDqY1Id1Q4FKEHB33D+7ekX77m701
pQHwfIaaqdonYMVMRZK5EqawYrHRtUtffItij0oOfcIJZQ2Ptpf5hiT6/0ZF+pjWW5QnxP7hPt3V
GnI1rCgiMR9O9atehYIRwXx2RLMPya9zVnAhfk9TfVGhbT1HqZamt+BxD4I81m6+B/00ZaK4Zb4c
1NxR5wk1ucedAnrZMjWhYYc/+fcg4+CcrffWpADuZFRaXoBo4p4vUPRPds/zXoQsSfDeV9edRXmO
MnQpTdxQe6FSCfUFOcSOMODpyu/JKf5S15W5HJN4KCvcjPYsoGAUlOmSjRdHI8fRjSw+OmH2LYWg
bbgNTMi70SKUkNniWEj7nQnDAY3NlsEoA8ybjG15nDtZy3BHUc2e698Fc8uod+5swbgYfQDQrscV
bYvf9ITkWVNnRpUqqenJ8LMQlbjLk9SzaxE6iKtbECxGaNXcDsxwoTrjQ0ZLNZH9FvitKdzmpyOA
olgLfAx2XJBgI4HdyCvqJBg1B42+jrO7ETzXAZxG7QPPxIqmHihBnj/hVBkG9kU2M3S3LRDhLMp6
hlp4CaWhngg7ROf4yEFIjG+Thxbu1RlK62ADnDx+be40MwYH79O9O8W4H232U9SH85sZb8vOjjGj
ZP7BGAW3DWI3CyuwTA/QTtqPlAkHJcvG5RZG3zUN3Df4Ng+sdAoNpiwU5Gv0PFdq05/eSEC0kiRM
zzuTNItxBHLkgNNVaZ0AfFoP3612D4CHBugid+HKt6gms9r1PrVvsZHJkcJFUq2Ctn1lniB3+KqY
OJrSnTtthfsJjOJiVnKJHBjSiyBXumBkgaSO9WOvV9QLDSWbegbTQUdbeL7WqvdFmpVkzFLwWwQr
FQUlC5GTCVER72mKY7R71zbTUSz+OMWOTnBvfB/mJlmFuxXt4kIyHnowgNRJiro9/aRqePs7plto
2vW8h3kFGYRqxItFooe61m7x7i32VOf/sQBu0T93UrUNwMpziRxqp0MAbf8FqUiCCiqLJGz4cySB
gCW0t2f4iKpnwR4GuSJBRl0yYcI97ZcgiwKxw7/hBartbALC4d3MDbau5PwQKl/OT8eiYSs8Xfs/
oesT7Dpf2wWUwzFHRa9gGnYazZkEGW2WDGdESLkqdRQ6cVmfqepy/lMd+ABSIIuvCw76dRh4W0rE
zLpQiEx31HcAYdvQEUbZFTlGovKslSaykwdqeSE6bFmLaTR7VnX5QNk5tsK7/2HoTktlGR5/WlX8
uOQx5KQNmq7yLJ5+2TjyUfPIbDpQTcFM1yIBj4ILxFNB2KCokBrtoGHAHYll+tvprh7jVj//gpGa
XqyScMJAce0P0dhKgSY3GEOGycap7jz9amSZcf400kkaMViR+Kgvtc0ZseRnCjZxvIim1y3qm1xI
gx3Ud10rEDF98TSYYUMHB8RYqCyHCIYUVCYv6ZLzyS7j/VtLGaJoAaLtCfHCHV1aQcOsHfAeWGWN
hL/U3nhZjGX9bjF7e2cpw7/DVY3o0D5QhbaZb/RERH37a1+ngi1rcaJ8CSfeY1qXpq07qIjqOL4I
tuL8K36CldlPgSGexFvcCnfIM4XfS+OSATtNNDvFHNTLB7rneXPlvn2LGeXjPcRmaYnOqDy9aB3j
yTXsRTU2f0cyLIMNAwSMMS1I52fdp/RHlVnkgHosgermKigF96t92ipwCoz2xysmEyGUJpO85rLx
hDC3RrDI1Q4W6a/m/K8LF/STR1GMCS1sR6jibzH6aJsCrlYHl0ysDdKXFmPoH/ME3jt8YZFzmknv
DDTaZeyE/B5KuxnYK6k/fXjDytwwb819Da1uY5HD77vqKG5buAZoFj5rSchZIHBKv2kc18N5IfMz
6NJUQ5orrxL75dQV9A6ReTPeSWtdet0o0WAwwjp408TKOPnxZ3CXyBKv9PpgY0880T9bR0Ae650C
hLGxQ+gg8LCeSiyPp77ikJ2umlLisZSfUDQzohEZniqjlaVff/4e+LXUYroeKsb3d747U5EML/qK
6GgCq5pFeh/sRsrQNE/oLBFC2sL4h21Ei9baZ9B4W0D5BxzuX2Bc7eMwgyRrG1L95x045sZtqjG9
wuq+N+xHYKPLYj/pcepNn7JB54oWDlbchMnmbyxPpaNsJ9aE1Brmnx3CRa3rssitwcquC4dnDClm
RK7LQiBhzfZ/OB25dr41siHpWNutWSURfxblgbVywNxIOdwv5YNQVXNssFrKpg0M89hpAluQbizk
I6jnb09ZVBo3q1C315P+ZpQmTvavi56VVEA6MlSf7d173dphgloZD7Ehibmux8olb9/SqWlAX8YI
R01xvbTnGdR9GBoWJBj3FbH/6EGo9c2f0JuFeGtZBtEv3dSUFpRH+1GrSnsGaSZMB8ceEcRZtUja
QNySlQUD0YaW+jh/kWQkT/zWzd80CFTKsDi2iXI+ieFf+Erivpm79Wmcy9Sr/xnY+KsOZ2guizfh
4DhpLsoAtbWSTz2fgEoOw1+Q0UHshIxHYsAy5qqbE/CE7ir4sqa0Kt82lFaRIDbsdACKMPNrh4d1
HY4XXJuRioBLIA4JutwCO7EveA/kBPoidTThoeOaBIVd/72QGpOpPahMT6K63bnOpgcsTTDeWpK4
6Ma9+APz10tt6+83NqcTgs4VZFUdJ4k5e4SjN4nnAqjZWAq4aLaFAC/lXod6jjDeR7a5MjE+0Vcc
W8JO6/ag7SjzjwNFNsHQEVDKJOTtU7Sfs0gW+oQNj/iAVVLiXAcVmWfohPbkbiOjcvRXPtZCkNzX
W8pnx2BIhf0wNEuce32OEd+dWCZT1iKxNqp+01LCR/DIWQiUWkry9XhBw0OxPld5E64eyHRA0zVx
8dBqUtawUUsxyvHkTzqUuIqGu2AWJdFcMEHkajUG2zXj13gLqD8E9D1JdVeYEu/ZxDoCxegXvajU
K1thvB/wuc+MUMPt2nr7pP8KIaUk6GLhixZcw/GpKEEgZWOGEm4C9izgGYmqLPaz8OAOFM7wS/RK
fRzEnAffHM77f4HzRFHfVGXEBbG/MqWkmwTLFdE5peNINB+20ppaqeNHTshBFMk7C4hc2JNSZlgy
KDwKSpLIVI0uRzUpzfPoH+Jilw4nr88NmAt0yMRr0cKJbbTo0XMKFKmZ0O9tG3T5Jj1vvUQb7y51
twZ7zNziWRf+uxt+HY4WT2L1oH+ExpZ/IR3YSK9+YsamEJvS4HWVKJPzEoY+jGyn1T2DjMtdOUL/
jyAtyh2vsGcQ8C9snxG/kfgJiq47iEDG8aFdvqtTVargTXxDkzkwpE0IZm06vf7424qe/ALJXgOY
gDsUmQj8T1PNdDaQCUfaDMVwqg2ZwuprIyQDDLaQzbJ5SmlEwrrT9ZG91WQutBKBHFdD3rcalZ0W
b9ep6U9voh/tJIQP6olEznEwqMKCtCMplZLCX/rcoDUL/aAH3AN1AbqtAUQ7ks/HjUGWuz0jekrP
OetUdw0RBTzXXJn/2Db/8OUtUbsdZQiR/ODXC5KugeS1b1hWylO/MNrcPq+GUK0IUHTxKOKBlqFj
6VGROsLuIbyDB15JC1uJUYNhTWvLZbp79omvlWvMLkaQphUnm9lvV/Um9XEnrp2PMHVokLRCP11n
rcETLiWt9wKH3G5/5T4l/TxZYDh5vi0sGanPdxIrW71DgY6aYwOAYPjYFckU9Pt5MpvCOET4GNV8
qq+/beRbF1BNnxmE3LTzU+AGkceYHZ2+lRaz4OdIuGUmdkLp+vj7pjHb7wnb01Bx12anxKpldgjd
BR4xu4ZJjLo2OKSkiA2ILkNGnpd6re+MfSYbZaWQRUS/6+sSPLP0+BdC1+9udlFyged025FKQnxT
zk1ZfURzAlFk+Tomkz5FQ8hlHvISXgfQUigX6hOygQ9FIH506oVvosDH0GxxMNdsgK4o5reVLlis
VyKSGujtws/mpkI/n7DgmOlAvF8dmgHa7vdMmFzLMFCeo576WFuLG5gA6b2COS9YDu7OCtx2oK6U
rANsB9WnLPDZn6XCOo+WQAFQMgmlcrXM2rY3YZSMUKHJCZFvfs+oBUiPKOYAbeycz+uzI2E5wppQ
AbakUgqpo5rytxoX21QInM/E3QhomAKQrT8AhxTKoezcYEzvodZyBd6eAmlVz+znWRjK8SQxiAET
rfV0x/QMdGwldT0UjoeOmN1ASM3ccB9qlRUTsvZ3Hjja6vJrz+ROwoJeWPHhhObsQRjUnvttPq9g
zPCQRfUitkNq+sjzDJzjjunFnWR+qq7l6UQtZ3eJ0yWkg4uvdI3apbxu7Ad9MBaqxlqfrKPSRVr6
RMIsavxw0RWHvF3gjTYheLN7PHIyiiyPd6zjvZjDPzt1hGz8vTsO8tTFHngUX5ni5sb3MRA8oGrz
x7J5oeSP4XXMtcESDYSYNaIzelhUi6RPPw/Xn2/Xyq3erCIVUqhIDzKIaH9BQ4GdHzhgEfQE2Gjd
Lyvag0E0fus08+2Z+D8Ye9Huft2PQHICN+ZtpkK9kPNlodnfzRpcp4Tyjb4Dw+inCW62o2Hk8e3P
WnISmiSyz2J78NcEQ5tzi8ISlQXZIXk1VeVJvu8hTbCcz7/M9QdV+vIAxMnByKkQyMmkfAc07uYq
kbPYaRlW9A0CwRNcONHQJtHvnnFRn8rgEs3nEZJAZWb4a3JsIksWpNB4LEc3q7Z/bmaTYuZ6qsnB
KEBRiG2mhoiBF9YYNby6/8JxLEmGQI7JKElERA2H3Oh9fZz3FTEtZ3jA6PVn1TqmPb/nA1Ln+MfM
AyEJHm56j3PKgesWA858ioUN+Oe/EqArUYz5J/Oay/SP7WeLmgCmGZo7/5wEXCDP9k2OGQnMpMVE
QcNvKb7ge8u1N8T9KGucY+SJF3t65pRBObmCEt+LuR6+aI03qXbjBUNDDXyR4xhUWQG4rc4w6UHV
c1mET7dAUwZjJznFIshics4detMg/3U5HJ+PROowlJ+8ogm48HC+L/lMFtUhIM0uOIyNI6b72Lf7
w43oGgnX474oYLEWavcQPMpX1fRsu/3hPQZ9JS8GoKmATnIyV8PG7TMu3xcdbxAL7ta7qw2ass5c
W4g5TO9pg5saP5dtsX9DSfZ1A5eUVwzKgyCBoBuKsMRcJ5FNLfFbVY9hi8NZWxBG6rfiE8wNfhDi
8CijW24nMEDzxb5A0JRwJKv6TkQsusD38fI3YiKqQix55ztXcelYQaPvctanvKKi9sxihvesYdQ5
81m7vUvzZ/MaMSXxYJ5Xx6JvAcFB8ka/WXg4ufoCY27WbDa7tG41mlJ8bHSiAJ1ttc0HXTcccSJ6
snnkOaTU7Tm7YLB12tHGiKEgT5PcuL1ru3tK8dYep+mXohULTCbvYcliBC9SO7xuOGYx5KweI4NS
oBYEKpx/m7+WOfRsUoTf8b9ufTDE9ERQ37nH6Xj6JjjB7lb1iKt4WpBshV4VCRK3ERflpbIst/PC
RHwi8Xfatwwh/7m8bBFq7LhveybYsqYd5gvKBA+DgzIX5wSjIijQGzaTN7d1zr9aq3zWOWsyNyMC
f67OCEI3D8jx3WmjnU78xzmVWzjvKtrkTzaLbVy/P9fNaju/sGyWprGFky9pRWRHd4NMYe/sKBv5
VuhLohdco3KGXmsIzqojk4lSU3UmWTJ8azOUgY9n5LgxxO3iPoPyiPWh0bFd7DunyM7bkKcBqlcm
E0rArr9Dyg0aV0joJ9m8iZVAdXwGlNds7Nm8QRkuyEZA/A0Skj4RYtIH+11KxWjEgolaxy+5yiFv
gO/tXslC/F1KGNKKTsEexnitBekXIcXqQm1uK6VaJ/Q1sVO0MlVNZh7VoZIb5tTzsBmBfeAIYGX9
cmbK1nr2NM2thcYD/XQnJHk9vmoTWz68asNWEL5Afbh70PmOOuOjYS8HfxVNklOPY4oYhXQ3aIil
KRutAdIAuAyEJv88CY5Zcniucviti8dv6HCk3BnjOrxAwa2tJrZm3Ivmh9jNW8AYHsurRRsuo0YF
/AO9q/Z0Np9fEUdSpR4BE9Zn71nPV8IDWPDp/ASZh9auFbVLqoPBGKm/nWgR9L9IkevQLTruEa5P
r3NFI1KQascTa1w8qzVIjL7UunCyXm91dSgOKLQ+xxKorlZG3GRXJiSalYyY2ztEBH9Jyoecbo+3
RDep1zTgRgEWrxa7JcF7hnxC+7pDpTwKZ1dVU0q7DqSomZILIcoVrkKD38SqqU96hPgwwC+8vwmh
qua6pnwsSqRvMM/DVfdplbhRgIlvz1qHWE4bxxo8tc6fZZnvy0JhTHtwS4B6GHx/O3XSZ+qEh57e
jCKarqO1h6N6fS1A59ESO3oOeXCKS6UguPUretwt9Ilhbrhed0Wp0WCNKWyHN4gXpxfW01qq2Aqg
wLx35i34G1e8dD7/qBXTOsKWe73frQrQAq6qqZDUX/6yvUkTYVV9GsFPSsgRVq/x7oNhFaRDyoIM
TNm3XkflGI3Ngbw0z/8CezHA8VbmSAmrjm9nV6hGCQ6x4u+Z+LpQFol+zYcqDpFMyrnR4IEYN2fw
lVDhRTlKnYPFodubdCo1QFcCXESMbp+3moM0xfiJkipMVoZpFhUoC8mm6vhAjnMmM0xwr/PDh22b
35Vi5DbPR9h4zwjcR6fK34gGM2uSNgUNxbDPOXTUEvKNg44MSrV+e4U5+IU4o2kl4Sx4WvEvMW0U
3aBhbVVPok6/jwwmkpWocV7BvszReM6PDumIBepVC+nIoIU4JwPVHDKpAJRTaPR0Bx9TmUdGXOv7
q0+uIvrrUAHd6kbaOkC6LIrqneNhL7a/3+bJ4aQcoeBJBTie+Xxo6lMmM7sXsqhbK1Rq6rBY5eRw
lUM/VMs/kKqR20BvkfH4aDbcb9jKKu6hT48HTISpu78vXMylngpIRi0avVhAYBgA+XdU+Y764OCO
JnH7UU7nx9/vqkYTIrL6gXUXNnSAM1OvyfM/cOpDblAXqRoFTKZJK8dNprIydd5/DhtO9VjEw5qO
qH0VbhR903Ec/HLzvG7Gc2+EGsMKBt/q+uxSkE3XxLJ+fasMlSHM6l7sv2isAdaqr93Tmt13aK2X
C9cc1bvfAbef4Kxo1U6NStXNz33FIjdd141TXu1ceFQE44K5hHp1J1ibvyUiKCgx7WHgjFfnfAi+
oKvJC6DmCkkByz7ps5xR3VggwShpjsnubWuFuD8XUiVruOZ9bwhCbX0KxiNOl9wcUy7GfobpmQst
2ZvBUoIDdmRnf5iJ/D3QW+bCNb0awkPcHB/0e7MAwd4pnhUClnFAIQurN6+b6mEj3CSPnQdM3oIK
aU//IwGNaqQEZrn9fbaxv1DVNT10BNE/JYaWX/tFWEj4zqm9T3P40AyyIubmfOUq2iSKtYAMcrgD
8d7BLUdJqy23BbE5l/RX1Sw490KPoR+cIyc4Mr47lrD9TQ/DyAbcv7BxlPw1uCMEf8NpRLmW/+Bf
7mE13sJ3bTOXdIglOkm5eiMa6KdARX/174q8nnuUqXrgHl0EqgsShPk7Qt9KR0Q9g1fKdPhUOGjK
XAc0w15/y7R8SMyo4zSNOPzx7GNFospxlV2wjkqhzoW5kfJNK2AhJ1Xgrhs8lMna/F2wnjLJnThy
kYON7hnvTlXmSmxFFuVv+xRMe4pgeTnby5uauXj1MAf2SnYBL1pfZH7J+BwvnjtJK8tnM0Sj9f95
0iGpFNssmSb6iDPcL67tsAOn3HoPl6/K/gkp2N3KmjJ3XyrWH/0yABdjkdae/o/+U49VAeSRi9Kb
LhZb+Yq4TZtdUfJFCxevzE65e6jTYzGd1IHIwV4DaB6sISSF2qkvSohyyhUTGjlBJ93yZ40iLui6
xNgnck84UP3jLNrAPhxeUgks3XZYfbZ7JdS2N3j9k+Okm4cjlaQv1Nni2t1qc5fqO8lnMYa/k5WW
aPRBPSWKO8xyHLORruu432s2Wji3GqUXesPHYvjYhVDZ4ApZ3ppo1aLzq4/rZXhjuEDrad6D7eQT
f+9rq3Lhl+yVJFPAW4s7rTGKVhspwjauIX5mTRiFF+8yk2ZUQ6YCX/xRbiGDxrR3dfbZwnEVP7Ak
z+gTwsUorzIjHOcrURiujdDNfbAU028+f0NVYkkbs+uZL/DVej/N4mYbRohnlsiIRh7wrz9FnhSx
XfnoD8fPJHe01BmChfEbGizIbze8ttozf5lswl9FnyZSpvcn2ipy4+g64HezXQ+5uMwmuS9qp/KF
9No6L4YF6VOwEjtUyvn9K9czm5FQR24+95b1StS4yZBirUOOmkFlfoYd33em1S/vTsdv0/ZycdzI
cFo9+jKzMPaYO7VA+g+e+zvOGlxtcV1fGzKCqzonMVejcsAuujYrBLVGPtFPDLCbVeXY54adiop6
oyLcpmMVX8lUyxW2OlshuAikmkkYH7iWNLXjPUYCP+UHZK5R2ftF6IeV3x/fLm5WUiXsIOgUJKoP
lAeqAH45GFFNfO8YAfu6u+YXcXcqBR/1XPudJnoXAA2LMuP0SOXgxj8FxrLVdpY0UTNzyOSYPMoF
ZGLt/4Zoi4kp+hoNPFDVmkKz0Xi8YdY718iY96Z4tX6H04jaO3MY071kYUr4u3TNApncLTDDdE8n
v5euUtEl7QikaF8a7Zkk7QLnQErcpeEMzCm3zj7yygbOCk+pm4wUXEfOAoOYTU4iBoDVZ9Dqhy8E
JVFemzkG6kAIXpOQBQLSR6iHrCg4/2Tfa24ohqJbTDwf7aHeKDx01CYbAr7slIt3WYW7yX1GSRO3
24EoJlqLs9xPJh9nRuwstEH1vCN4YWdHr5LUyg79qVRwIsN+SDvYfTMj+1dLFIIht+XP5IymnolQ
Cy0kqwAaIRvSKrDFvKe+VFvrVEyXLBoqWLu+RvzZcGKICQP98L1pSrYNdTXjvvc7RoFu+Dedg58F
StASCpIgBKLog5OGnThlAa1jFymlJllCqIABnFt0gXXiTgV3eckyGqOt/adkvm4mWgfKDBo9NL+V
Sfgdt7TVEI368eqsP5JfeIy36Lzram0DKmsCwPSWW2ByXPBmqtvif9aPY0HtWzN8DgOn9Zs07CwI
DqSPWFnsDiIbn/dnmE+KZ9Qc4dL8S4BQ9ml82rkSUr94ysRm3G9j5zAo3+9ax8SydOAJPuZa8XiZ
AC4xnIquyPQ6IWOSmAWuIJzZhDQNw+Uop3Spd16rSu+k6gf8HSkCin9p5k9A20WyI5/ei/iQ8bi8
b3Isu0wjDws1lgKYNx1VQV4qlA9UA9/7IaLuEjLCVIjUuHjUTbrEaIgqMNK36vWZ+00Torbhn5TI
IHTW4Op2A6oIEBh56TRRFLUtr5mUFc731Ot4JrSv2hiyLTGk8HXYzTmbncjk3VRYIi3t6vEdx4nU
hi8PbZFGhiFqkJo84YHXl3KSI+5lLnvY6Di0uDABe8jAXIjpEBTASMeJcSZi3j27BVVmAp0e3Hh+
Ik64bnw/IYD0Ht10y2UyCd3Q9VTkQMlZ2R0vz9EXhSwuuFkgH4Eqt7cMdNi8Wo5iHdfRmUWfLNX8
rSYWrAiiXh8iFtjhGjury8R0twypTshZf/PSaJOy3BId7b+rvoPh6uq/iDnUwdJx66hRgfn3hjpw
zPfgP5nNBjVMAdUeDXBlioTJPh8RcBlxj3ckIRPfvK/rCav6ENwXbjbWlgl63z9w9aG9emchIMQM
jUssfm8sIQLZRP3/sDtEsF81adgp7wW67RiyhC6nrFH3+qpeyh9vhy1A9eUdTEgO+RBHiL6Qok3K
3rpK0STJsI9/7MSUwOCFlWeCI1iLc2haa45wsMlaBXsgb2j3PBPc+qKrEzx+03r7jDz41vJIFwJN
O948OZgfmFU+qoHgyIP8bKZPaFKO6rHzgRl6B9eqPKpd6RsIa+cvTISAksGKWQ1amzTvlCk+LXKF
WAxVsanpTPW5wBWq0/sCOe8sH0nvX/euiZPqiSC70O27QCbyY15V+xaO3xy/oJhioZE6V1jCv5xP
JP12z3DnszSgIooMUNjC8rHaj9GP83UDHn0sFcPY8bYePFaOAksExNvgorKhuViKhqHQ28LHWkUZ
SrmiOI4wWyEkY/DP4tSFrUwBln+Tl/A1qX7OXuPH/thvijA0fQM6iFkJYiH8og1RY6nsY3nFXBHp
tOwSCfvA26gvLtSmT71aXpIUcH8RML5pKN8+J+ZIoa7LQWtz4Ncre+fEa1gHlZU0g2JBJw9fAunX
r1+pCcHsUcEqQ9Ohi1my3TLU/RfFiFRiTtWDIO4nKciD/Z6Ko3qphdQnh18M6uoHDcqp3tVbaoP7
5OrnIQyXl8TF1OGr8UYbqlsg32eZnAXyeQpgzDjTouIE5JN16JhiLwKgiyCAOSjCwHElmWNQ4Wag
pMD9bCTDdElufLFkTt+Kk+6e700JJxjmfCncyk76uwaBxjcklyBVbrBPgOpdwagMPDs9sDEJC3ij
x/DqNLazCDJUogqJqfR+rQEcLGzqh+6cuWQLBPFvJGVuiHB6eu2M0euftRc+Tr3k7GmfublAygd6
cP+BwnOT9QIEscavO1tdjc8Xv5fxnK9rqG/BbZv75PZ3wf7aA43bHCRevgBd4tEhc1aWsVSsddWK
t3IW1/Jna1F4Xy5V8VbQmiSEccDK2iaSZT0OtOapM7hX/8EUeSYHzp12Rd74rc2izwzfn3oewGYE
Wpv0+n+rIzM3/KhttD+4bK9hcxFax0ELmCYdiXmcFjG0E8iTtYzwrFjJN233lQj3Sdqqs6TQOr8D
mRI6Rf+GVSPgyRpnywTIM0YdQB4BUlhFxkjoKOiybHKW9nPbxlL1RwKAtq5RLzqzbd4XmEhAYPzp
jZYxIZ5CQJIXTVZACuX/kufEGxeRyl4d8uq1z/ozJiUvPYAO2qNYqbgVJxkfwDv9zm02UCv+ddqr
1KYGlFGAvtgQID5QMEYYNNQPoJGDwdD1fbRdX6ykMBzsu4EfUMkyTkKj9wlgo31VoFZZrXnFgQqA
dbR1B9e3I5pYDkRMr6Nm8tnp3QEvVHA3aRcxd08twx/51csZhL+NQXnYDEDYq1QFXeZPEO5M9YPC
GUtex2BCuBUuSMaCEa3U45OqVk9Cn16dd5xdM1pwzGDBqmbzZhdPfAJ9oyUPD+xshCM+acmfAI+U
QU2/OuSP1ElTKDK9dg4La+Wfd5vgTce8lrK33R6CQ22mzt4tKsuvUkLOItjB3yeREXbBmmDPTGb3
w/NCFY/ip9Ep9po+ow/q003TY8CZ6tCBj5z5um01OkkjdOvo7dX+8VNhXGJurwX4yFrU6A2V5pRO
fgGbz3rUv5nSf/qFuXW8V8Uxyw3YZXDXaBeg5dlX53CYFJYx9eGODHEKD95cDKJ3cADZXbZSIIJu
jfnnDAePfLACmdCuIXqEqxY0cs+EMTc2huYUIhQSv3Q/J4RwusaCd58g7Cdib07boAXh2e/DjK4c
fKqx6tafW3uyhJ6F1APAF+UHxQim/X4/Nc0vK2OqTG2asbumhqgK50Zrb58cXSUeipSiBhObX1mM
WUx2+F3blT20BwimavNSLXoSzd+qbtCUWnqnhACTEsu1QxC+0q/VRupZph9uDdy7avx/f/AQgH5C
8r0iw2SAvzdN0arJJD7nrKrMEfqGIryH5p1YdaGX6Egp72T2ITWPos7USZ78Xfj2QUM3q8cy5fYv
qdMzyhqQivgCBrDz7n1nFM5Sh0TpNwqD41Jnkyco8RjYKpp81kYtTR9uxTtkTm3kJyLLr+cYVrNO
ffVevV1CIm1pOaJ0sYZi2nCGQ6bapnE7puIjBIg+BHBDTuexSUR4ZHHdhr3Ny8+QfZaHGRjUz5IK
KSwbVfulzV5I8cEHmWIwS/H63InVNYGGLv8TREM9CkKhbJICsmJCA31woE5bwJKwu0kHg1pe+WAH
y9RG2pimbrJY7RBcVKa1ItQSUF1Z5bwAWpJD0foBrfyjJISJUYyJAPtCh0JsrWrHbECi+a0wyejh
+QnfBRR5rkky4V9QpOBjtXmy86kXtPbLTN+oFbPMgS7gHY//QiFzzcfGoKnKMdQOQMp3OXa8yBJB
13Cdq6iFYof24/3KNaidza6OrgUMn6UuHMHn8uW2j5Ukvgb4jd4pF9NGIajF9yesKiw8DzswMets
Qc9OI/5zvDRmldTn0msAUUgucJnaEgSd9cRAf1noWkL8HCU8J8QXtIrTXsydUPtlOgGj+jjFcEZi
EWojKBhOFyT/LSaRsrBJKCpVny5M6h7HR+cjFN0EEjLShf5QKNaKM1U7W9s4d/LyuHbxcYi6+64h
pE0dYq2ZqlEXzFFy0FtwN/rnB5Vaw/eae+Gr+ZVO/sD5ifqShoqyBGHo/4xiO92PSbuUu25HHsf7
Owc/xgKADZ+hxysazBlCQgl4ydLnW+fzJDVAdzSMQdev5+z0Osb9H5o8CExJkbz8tMoecxKo+dMi
oXS+JbA4MTfmgHgVm5r36wsegx+eta9HcrbItC3GQM7O1mWdVo7yJjj5nchgCznTxyKTWSlUxJ9f
jwvNY3EpwjmVsSygs9mGwAQmkBClXF/ArPKdOMKutIIfnH1VkJTSX9Bon7wF8pDSeCAc/XkYQIaO
dCseEbPVI2DuEr9W9fpfxkLOpheQFPs7RxQepmVFcyE45AMFndb3imiRopO15j/ODYZmDJyx6wDn
P0pgqczbEBEnJI742fap/uFdfotB1FKY2fdnH0Bi3u+Jp2zccIsbyizNbGvsi0LFzA5Np9hL4TNw
En4X5T2GObqELNyLqAeRWi/0YJOeUTr5bfM+Rxl+HnV6t9Fhge9dpDcc04rCD+1BQQkDDLSsxrbY
AT0pQSwbVhkL/K3ydXWnyVomwgic7P4rnTYZpuNa5+jG2BmnLjgY2/xcYnT+6yS14ABgyY+VtPQH
YWmvNTF2/mn3JYjyrg0Iq5ZUqX4ovybXkoJ+3s3mJG61Gs2OH9AGrscfEspmS9TiTqvEtX9LYR/a
RUZVJNTns1563bEtZ+/+RFRLUFivBQaKRFX4I0C4uWBWas2F2TeHBGAMyGwzSGwk/IbAFgAAmR6r
JJiwkM4Ugg8CD6OQrmyvpb0hoD57ymMmhwbDNFry6LbQWeo6n0BZTFElLffCj0grD2oPm36mLWGC
ktrRo9KJfFZjWIrkrElpPIrkyR222hdpmBN6BhYu34Ot7gr4+9j8PFzFJ4+tP35T2Mvco48SsP9Y
nrb7Tc8H+O1pBkzOqYFvtvArQwfbjvxyHnLFnaHE1J8P0SqNTOG0uAkwJkzBRYmwEqOZE2sjNkM2
DcYSRtoS89x47tOdupJ+uN1eSdIEZCRH1ux2s/6pFIdvcp1vEEboj4XAgpc/qbRtbyWmWLMFgEj6
nIdQNHoLX6j9Tqme3aRHKA8ZRnFXGH088pGKP/xNN8YQTYyRZBQiTaw9No9QGFp/siZUMzMjiUTe
oMtJ1dA2POqnT2TGhlL8ho6COfCiMdcrERDwzSREC8+MqbOHFkiRjL7CutJunFgZzlNjD+iyzdEK
JZBbHDQvH+BLwvAar8ZtTnWisEzp4Zv7N5JmkyllxMJOXiP85vBzRGkWRBl9dBv+cA5LNaTCNoYN
d3FnC7vd/tXyU5MMuW1epCXsreupNA7M5gbWBEeWFnq1+GF5oyNqQ74USLERTylHBGQN6sZS51RA
svKmKLSgWCzvWfwB9P9q6DCkE4wwBUPFnNRw7e4s+jK5Ose/8PHMjdSsmnhp5d+eGAsUrLkN1ORe
VAJUIlMJkaJufffI92SjE8/5kKSgH4rlObGRBzA+0eW0KFrk8AkJtw1323C+hvy5eTn4PXFf4CCQ
IMn8kihtbUgSr1hmm3lvzzUPs+ID5u1hwp2m5Npum/7WB4NFcUYt+97dqTUlGCkqZLFTgf+FFfpm
jrom/sBqqdyRqvZwKUTVO4ooyRK16bGQzTkA6ffKWgpfwtMywTKq1J4f8sFPYAJTVMKbVMQ0a/Fm
Cqp7k/JFqqsabguMxyfQHVZUmkhbD3Hr4eAP5Yl466lyUdqXRgyYdsCISZ0dGAGcRYxRz7KWZFY+
dw3VDrPAGBhMLsqHdywf9w9TcaugSVSf7SQfx/xYomU2emjrENJKoxaudBmtlpVqy4rrH0Kw/qIv
lQRi6AbbTbTvCanGJWzi/nAJCyE5MlD0tHZx4mu6cuHT8eUIaeO1FdLgWFIxcTR2VzzFP6Q4Pu77
CMGvG6weFDcggNCD6zshtRZttlBCnXPdexE5dzgl4CexvvQ3SL79AEKbMKUqgwezTFdZarFcK3Hg
08xW/kU2I7Kq9+F8L7rK7EqOvUSAtuzMzxrdnQfA+yyTFZOlId2IKNmltpax0NheK11CKZBFdLmc
s2pbEOr7++eWdUZ/vLgOiW+xwjqMmlipG5asQwT6T010P0TSLgd+55gjJWnowuFqBp3mYeqD28V8
XR58AYtw6UijE4lzPi2SpfB5c607xn0O2oZYuVu+qvCPKU2LYe6wGwrWgzBBy+4+zJhabloioLCA
xJ5uo0S65JkecmjhGQmrowS1fRlYKH5ZStZTRoEbTUz3UQr0MYfHxP0XHRQzTxlePNVc1d9AOMCQ
2skv1X3SDUgvncHNgkRBd+LuhsHiXsVMT/Z7FKh8kjMLz5gWMwI/eOehbkH/P3Wib3lKGW/NwacF
hmGnZ5XPF0vironet++se8wICBKC+iPemJq2Cwn2YKoL/l8KSeGfsUwKptxb59tAodF7EU2Zmr7Z
kOuGXywRryo2XzR/r+9niFPp9wcgZLXPmv+Dh/95W8lW7Uxz+pWVMqudk9NRSuP4QoHevLqvXWhQ
hlZSk5AHPjx5uzsebaL2pOY2ZbBXKq3KN9Dy4dLnNy9YPnuXIf9zhvwTtF2zkTiGafqR6HNoJJus
A/Oy3c0lbaJBQV3FXRVL8xJMpmHn9wmYH3ehNu7hoWYDKdEN39E7Agrps3DoEhcI4Gb1UZZ6ScQ+
Sh1lFJ/fUPb7gaQS+f4N1S45NNxHTS4fIE2Sa4+URTqG+0QhXxp3JvMXcQ1MGnIzgi9C4YCXtQAI
VZheb77jI6+FNDJkAlUYnw1qmDYe9SN/IykWTPMkDUK250BkdV/aQ6lDStYqLv5bk1k09y50UadS
gxRfxQknVrlre2cS7DJRbUazeWoY3jPZfyikZ1foQfTMGUBGHDLjKmhAnlftYBGkpEba7zR3WuQn
6hUCOHqFTaf8xFiTo/P4MXm2IYTkHTRwAYXZGM8IHH1rOKvw/eJya48qtMM0AiCqhEY2D/h3rDZ+
sOWTAnIObfEFXM6il4OKIoWZqOCx2di8oGg57JNHig7xNjbmSZ5ZrQ2Sv/68X+mjIj1cvdIeGovj
UZN0jRhamHwRB4JZOwpb3/DeHXslTcZm0noJYw3Lk59BGx1gwdnnEK+jivVSf39oSqDChcOckX0a
QGTSI4n30qcHpVpqvVCHWYDcGqDEYObOUPrD+OhpQ6k9Juld/dj7FSrJw2wSABVAVuyPpAKr2o8c
b/hRHjcGE/HIRurE30okjgT5RbPXdcSRcMNzzB1qFcdJkgDEJdnK60gePrqTMIgXiOw6cj0+QpiJ
UJKzlyDR9YlydtwEV/iiSQN8L66OYVsk0klyYrtdWoZMvM/5lQJR9t3yGQemkxnFiU5iGfSy4Ilb
zso4lLlhvvudbon13XiG5oEK+QXUwqIeAjqrUHrc2in8DqHATcqnED/CO1/UBxOciTOgPQzB45ss
4MNGDbmhyRifAdRJSHbfKmzDbheaPQTEvFYAiisaKnfXyyK8HraDsM8CffFSHBGdqPMONk2o8BSE
O57zG0hOiyVRN5jECphn4zuce2LtUAFmVDDRzjxrW4tk0zW5xxQnQdsMg02xryB5f/DJ3AyT/w7T
0z2fkVbKlqij0NHyT0aBVlA+W7GcG4I4IoYUrQNNIUjBi89rMVC7kxCGvAbJPL0kQSV435bisbcX
RuBCq9IYZDzE/3U47ort9f2Ze94QXUo2bLV6YYz/k8llC/89hsqZR4UHye7qZXOfxNC+noLDz/cM
pwIg+fbgzejvNzaFaH9t2GB71mt8fLSJk1zT2p3cr6UeYE5Jx5UR1GnnGaED//ml2gkXmZ4ElUG6
3/+zIeSHAp+OSXa3vhtU5xmbvqfZ72pnWb1IxE6CBwYkBncOn4w4I0jdYk9z+EqAiHvd/khfSny+
oy6R3CMLcEi7hbQmDxqY/+6XXo3Q2yMIzxGPn6zEufFn6Z8PWwescCht8jnL87SZmxUNcb4x3rII
gjRrfwmeJlAxhPaNsafBWB18vY4MN87MLdanutLx2himj51osGM5wNmHVBxgJZuQ9XrGPBOhQwYo
ca/VU/EEKSnYQ6si29fxuthGh7lACvjALJ4WAyjQ0RxLHK4t8I3V1LV9T7yFhl9otiVHBePu/Zv0
di3+M/RQpiP34XxB9t8MPC60PR2WZTmTI5Ns+n4jTTKBfZdLim6gHDJgIbLgh7LphIddNAtqHRsk
Doew8HS2X/98KpV/utqMHLebSGRtQVvox8qwhpL6XCMWKRlSDoFYMkzKSr7e8gfKpDACNwAzDjyp
KsEPkAVy93tZfD9NjqF6rlQlxOastEdpT2O+f++9l07YwSj2RUaAz1C32ma+NU7Y0nnwsETwtTY8
NfstD2/h2XxCVBESWEVpjEbrYsFmnO9k7NBtwcEElvHdSqXvKeHpKC4du7RFQunye54kl3Qw3nEA
hcNRbjJVzEuIm7+vxrjkxgZWJjhhz94ZZiQwDow7yFQ5U3Xry99dNj5EMellsxdV7ogJomu05L3S
V9p6wGrH73JPrN1xLblEdW/fQxcYdC0mQusBKIdptvSCBqZ7/vPg5clsnSdV/ByxXwWdxMJ0cO6l
3V4Bun+VTp+jx+lIv+edUWs8lqaUcnb1qeCC61xaTxmL6GJ9761eQPmns0wTEAG0prgVcE52OExg
cKfAgTobHEQugUS8uxVTxNRzFMkIVSUTShbLCASlAhMLDsFZsETh8oTb1CdmDR9SEWUa5PyMNDRF
a1jxdYZd0cuPSNAcDX88GgtRYgbW/9LetmSurlueLXuOlzx8cbgDZiewzDgpBJ1X3G2jdScKYLzl
rSYbFYrFawYSvIDqjcVNBH4qtKXts5mbgbAv+2cSfoqs6t4bSgM/zu9vjzZxbTtWHtGGHLVQeVGk
hO+3oTO/1RuDW9RbuZApXO4Hrgj+HEdj42v9cDJ0vX6lvw7EcNC/NGux44C+PK+CfeSdWjUdp0A/
Jxhp5KVl3jO6VfCb7Boyne8Nh26PcBD5gx1853s3z452JkvFDpCOMnzeQ26wx1q4mnM/ckYeptog
VHZ5hG7KIki/fiTuHtH8gOa9g5NQ4D31FfnfW7kLwUIff0tef3PSWax0hTzaMTJlGQMByNSv9Aqq
tji1mwQo0/UHm3N5zsZKiShi6wcV/VE25H41itK7ISbb5DQZDI536e2lU+V8Qa/rFelBkZS/ycdg
vT7AP+d33OuIbLbtuBxweHm7SFxObYWfVC/SXVWpUuHLkLSa8kAgFwi+t5byTA8tpfh6eAGYHSjZ
YA1VmYVNyMCX63tPvMwsk94OypD+KOokWoX+I2fQN8/hg8nPKG9xQB7ySZz7wKKafmfI3kt4wv9X
RAzTOlDPms68g9+w7v87Dyc9G31ocu78dCpD6d7CWgOiINHpiHZExZvQOtPGshwryJGJZHdUEumS
VVDQ2Pr3LQ3V7cZIpvp4uPPPo2EiFinwgalqga+XPlg8TfOxTyxmvEvAobATHjlfid8khm7ry+BN
4Can2ePqzSGAWinXCgNCBWiV2+x5l2IN3QqZUtgjW76xGkZvaYVx1s30re2P12Tux7yEvfsEKhG1
KL6m2flY4FrotbjAZPZ9QG8NezRc84cn4ABr9Zv/CKQ+C4CRTNeq7m+2ibrYt4cGSKknNUBE3rB3
BQtRv5g6+aqNLu9CzcxZtWailtbX+XJ7sQNFV5tl1DuY69KDY2Avtm+YJZgdI+sO7yxcE2qFD0Q8
zkK79pIycAM1dNl/K5XBrXSA/Dj6TKsU0LEgw8/MvwtsYR3dXnlEiaFOY0t+Vtsq4SoitknNYXgx
T4lg+GDNMx1H/Vx9GUx/kbakCvf8C1Oi2eFaEolhXVUHshDzdGJGOSpYNy9TcX41z6bs9/cHIlqs
hEJuViT4/MQQ/LtIyLBXpiOtbjBYxXYDgJRtSL9k0HisZJJn3wRh7TIRXVQOTryQ/AV1gEvaw9Mc
FniES81nVZ8rThFt40I0KlpvBh7DeSyzl0WAssmJNq0om2or748/HXzO7qnDkDmHhtmJ9cvnbSI6
ouxl1ANdQIaaP8S2rgTdGVQVMbDOPKJZ4IAEvEODwZYklOvP0aj9m05t1sb2DvoOvx3hGRFc72Ci
FtBIBr0yNkMaj/oSRc1O8NjRJlzzlCJvbHiWF1NGnKVFxPWZ7j28oJfgCwhuSKCVDyC4acnyj1VW
GKTmg6myOy+K5JKlxOJFnQZCrGXlo8OGELfZtqWb52/G0lPiBFacRkvAYLwrFhjv373czPsuoO4F
U78okinUXaKcJ7lcKGWLSaYFLLGXonyAnPsfVG0nvgRcNzewIkmr+4OArr57X1Zx9UlmeWfv0uy6
RQArFjnCByQrFNpNLHJeks9Cr1m7fyHB0tWCLZthpAu06mzIP9e/dI55R5u3hleKatK+uuJq9don
R8FMID7x1n70xOHUoK7wIBX/nrjWq+evcZNmuY5FRSdf6f4Pzn9UxAHhcC1QBRshaQF0KoQH9tTe
mJjlHEXVVdL/cl1VotSpLnoO8Ipw+CKoC3g3F7VxUu94i/rWrq1nMsAviYmo5RLqlH5/f/ZsAahd
JhtlDlOXwgzKX4pnEItdcKYRfBrRisxS7s+3EI1dPAGleLRt8vJapgAeWiNtUI3squov9xT5+FO5
rh45bLlJrkD7utRV1+DJnurinRsKFDX00qkXF5oeg/Qyc4+Fayl89gEItGWbdNSMuuoeLKy5vHjQ
wt/8OWYLMnzbAy5pbv9aO3gZOXZOWgCTWAZvVs0cOwTNl2LurxRr1u0Q4xx2R4YQqVdsW0XikNXR
FHFFwuY4cGidUu0RdK6DO3jvtDdjDOl5kAcUf+QRobqvxV5yar/mzqnYclLk/qRgxlJn7YCEN1KS
shiCWx0nZn0UhyLgr5pnNZyRQWpx/mW8znXd3oY6pQz3vyFynbol9sSE3kGTKiZNiwxIuES48S4b
MfBUVhWOhActlVQsvnLzhluxkM03wcN8hPElHpO2zkdLJtrbdUjkEiXUGcdx/5OvDIbk7lau5SjE
SIcqYR9Qiu3i6zRdA0mjNb5NAqrcmANviZmyqm3F9R2utl1J/RtI8uXrPVO6FxTQqspWDXyH7IXf
aL/A4jJU15a74I1f90sPg//Rq0zTPFx7V9y5wz75bfUCoxBGW/WF0oTDHJX0x3dsCwr+wc+JCVSU
b5/9nCZXED4nzzx19QFSaRAHIvJvbKgya6mSZj80b6RDOEz02lCmJiE7wqvpwcjOrEteeijEwIwq
7KfQ3WFCzU9azVKTaj+ET14WRwNVX10+tXZ6Qhy38Sy+ZJXb5/Urdmb/CUcrhWWPUxCNpTUnxqED
f4MBVf0ob1RMA4EUCiT3YwYIsUVgYMHxfz70HObcTwXW57o4lY52E5sdcvgQ60UIBCNLH5+mmh2n
4kWp4GpGtRkf5VVZzlQKeCQNiZvitzcqdtPZb6z8Z6nEsHum/0SjEk7yHLfvJtmK4JTUjE/Cjct2
QmbwOYNNQB7pCCgzwJs+x0kNCTgjl7qnel8bBykSEmv1M9LJwmuXVNee/8t2PiCR7THt+OhQ2gwg
p+q9WW9U8qhnkDqtsz2iSTBWwFlnCLb901SUuuUUEpDLxsbqrNCO2qr1pttDmqdgZrR5yAXBx1/c
EwVeSgRTWT/yUnVO9Ne2b+ekH7RHkFWeasyZpBNphIWVknHaNNIbvoUN+iyuEeRRY0PmQ9nDMT5d
UZL2OP4ztlMJSWeRs0OLB77Q4cx94PY3y6HBRtKtRQKZDFKea/g+9RNlyvtT6dVqLoAv9r4gH2Wx
uFn/YZeITMPyuQEEwSOHQBLzLDKp3XsB8fNrDFeEXvTLzG1cZMlmPnC+RpQNuMmMT+YUZHv2eetD
7FfEatkLkPAv3r2PBlUfPc1icjM1RxIwYcDuXTLS9/7ZQLPmHcaLpozNJ2M4WvNgWMZIHyzmgq4R
JR0qim4MXyuzqektEFNho2XnVp+31/rvsL7lwIAG/gXEaJFoCqR9yZixgYmGFviSjqPm48GqJ68t
rtKf03RgTu699UfT7aiRRPsCR+YYSsYZ3cHgf173S09/bDlEDioL5WyY70sg2wvHreIXtZq1FSLf
+BLPp9HM5VeouIFFJwM5tZdYZAJ36ptvDG9AOMw1LRZSg+QJdq/mCc30mlijcDpkJBL1Rnx/WN5A
TQ0Cp4v3RgRbodMSq15tr54UR6no/QVg1BvAdeCzdseLOb+i6h5FIQrO6UKBuHC8RElUqxBtphCd
RrwQYuruINmsdR6HwAlpwZDrZnX53kdESRpcMKVMyLCRBayQCqxUrtCNp53SBLIu1LQVFfyf9FaV
9aA6Cg++/dAMWkqvj0wJdOX/MGAw+dTgL3mv4k/ik0i/NIYjnsYc7DiJsFIygJalzHNPkBS2ZUui
/lLKcRMjytGT+6PxVPcTpqf+byJEgeo9K0A2Qw1L4CBOsWo8LK38UxcsBZfjEoawLEG712XnrM8G
yeRs+RM2KZvA71EKXfibbW9AedKEDRv0J52nssH7WHWe4+WbB1beDWXGK4+k+KwbZ83TibuQ4UCz
JZKfTigxGKy40mJzuZU5F16gn/wtscwNQXIwtY/JMHsc4CIxuFE+Q+WKlsVMzQSfboUkLEJKShbI
8zRuApkZoN61C6P4+krHYe5jFtv+0Ic6uZSyuK/63OjeqskTNjFNpIL6Go32HBvNJTRsk9g+crSQ
ZkLqrZeAmtJgxmSm2OgGtiX+wKlnUXUDiaz5jz6OY3sl0cX90DAULbUTsmjOMMKOEaJmTlCqLUxi
X8WIINbMNSDDKzHR6kfl4qtopmytXt125WPZttmeKPV0M3v5eGN023NE+7uvISWfxDI4d7FgXSR4
169h43O4Ne2quivHcmTfilUQfTXSH8+2RozlAaF2dcD+Aq+VlujkSZUyUFEx9brHDttKWZpGjrKe
7zh+82EwseLN0N5RCSQG8V9qJ3jTpNPMYbppLOlyaWM3xUfmeKTlnFBNozQCU9Olny3ajyDfeRVk
8E91NZljqzOSVaRYsZIv9Jwy626ZwQvsFB2DFPggoO0QRUsotQhgWzqUepUue50P1xmSB7mF3XHO
VLGw6MriXSQGr/X5FE44yZ0cX7Ybvz6Ukt37+97MeTgQXswpIoeZg7LNgfGBewZ+Zly1nPhSBJQj
osK2JLzTVsN5PIsSHp7FVGxjQLixElMd8dGwkiPaf/7aH+oD5++wUcMELRAjm0vnfqZrhIrP5A7m
pYJ5shXMzmW9D6BMjSRPLwmAU7aZxhpt3q+stF0QBr+7j//m+iChztr+hWCgzQb+lpULrCvRDKda
9sxsP9HLl3jNngmBZo6u5K90gHFbQvGDbUN2yeQP9PBtVQgQocOLlri32E7jnVG26UpdwusPh2Ns
LGk20/l7P9TMhBYS3tlmm429w/Ts59mXbtviFQv3qWziFrdFoeZW5CbvUdByveWPAC/tLofI12Gt
UKEjURZifcsi0gmB+pPkCjLSDUAoRz1PZLxKuDvGWZab/31XYQETIiJNKFsEnaa0r7FYE/zqBjZ3
sSATevrPpFDqoehMiLwmSPOdnOlXsGryw/eEkIvGy74Ljyu8Ua5zuKFAfbtX7NPDBB4tgudh2Wf9
5vE48gda9//glgD47YpiCasiQJf4vqjgj9CWkuc0kwjDpADXJzSyaOLNzhl56RYjDSlAJkHKiwBT
asmewQ68d//wod/s35ObGf1PY3zBQeCiUNrz5ZoU9sgYeMQ7jrDg//oi2ksWv0WHQbmUWMgJLveH
xhXDFmkxHxGa3QlJy6GvvNg5l3e3hozZHXBp1i2bQJLTi+4elZJdAFHVz197fANYIeLSTodzb6//
UPs/16XIG/9e6972GeWD5ObSNaEme9FGj34F4S8k4MZwYQXufywvXD34UqS8LxjOWbaVor0QdB9b
7eCktH+50CbQAQThye+BWNIuru9VqEp6Ul6SWvJ2a87aVlz+1Sz7cZXC9hZDkjTc1ZB2TsXvGh9M
ySLFuGHf08AHVuGIc8xb0skD2GjVVl5aaK0Z4+pWZeYMdKezdmKY0vwIcB2xAWfcRhZMdZejyCWI
2TEJsdHI6YdGWPEcFyL8sXsuJEeIVIULvFpnZNTkVEBk7sroyA1Bzcp9kVdYDCbCjphQaRbhPHLA
6dXErHpjD1RRCYqy8iYB44CQk5v0qQe/1nFYPRB6sMhA3jmH26Wn5NO2qFt1MbCt8caA/6YDKNf+
Ip8vBTo/YWhv5eYQN7QuQkw/iIEwmFthT4f9o4mFAwM/WC/8Ebn8Tb2itLOhuSGvSrtfyEkpW0xY
hOqpxbHsy7Gew509EC/3w1aTD+aCz/PT++Fzs+gueqdvOPoEl/fF4ae69B+h8DqoBSO6bFrP9mcU
dmnpJUViOD/Zfhutr20MCQgLS8Q6J/bzBamGB8gP2uw9Aa11Ntm8kgtIDhLK0QGN+x9fJcNsivtW
/UcIJ2kyQszjWNUBvCst0Z/ikgG/iescGlvSZY5af4CbhOYRJlZr13U1Hi4WziU4UYvMMYCkGSXC
jSAF+nDDIbWyKdkB04Rfp9WdCHRhsER+v5EkajPfLKvw+bmqk2XybuYBUIbnuvPVNr27IkuDs7LT
1qEo96nN3ghKcK0VQny58szKGAXdwyIJuqV860wQrYyEnxBtAB4zDVbNtFUsXIpFPSuBZqPCzQk1
GIUHrlXasYONoLa6Ipyr/FZ3wSGacgxz91b204PZjlRhWtq46Q2FZNXhdoFWMdHAvzFNNvf5PDvJ
3GJ1R+2PhLzMlapUvF2GTc/hOmRO5+pAyT3303puCcG13guuVcRJ2lRFjJXdEXc528KSqq/FQtFg
U3yZpKI2eDEAbgL3K1bk2khbOYwhkXew8IhTwQMvdNX/MFGjO/zUdylyiC3VJ1HiK73YwedsN3Xs
HaHrZOsC+LtQZ5P7rzPl16ZnDe+AcAxRq+NAMoeDtWUKZHYbQvbIYmgm/CQCfieZEh9J4Vc2M7zF
uPwxUkVW9hq/WcDZdgYC6ktEcfm8PJKQ+8zOzbTudSBfWvuz+NA2CiFHHXZLFYfJqpbA7bg3a7c0
JRpDvoXufkvelG2ZULvdJMP7mwB1jXf5PD7oUnpPv+P4/+pUKXyIDwCuo0d6MW+4sJDxNhvDotnJ
omzZzmYU/eBSidu1+NQwmmQYxkmOglo5UdI2IgVn/s0fXwcjRnhIjoKcmHsdydespa9IjQ+w+0rt
QR7wYdJAH9Ngc7MBN6Agleh6V36UsI60ePA+JrcE2KWNH1FqxpXZ0SWA5gvr4rAYAHt0prb9BIJ4
I+Kb/HaoQbplOEu2d0cSDTISFUFbDH3gN2rgbcCmS2We0bZjZUEMfmgwB5NcmR29MxoLgtr8aePY
DhlyVEislkFRSjFK2hY0Yb1JH7ROIZai57DJ/0FkhRb/3SWefi4ehER2MkYfEIRYmei+g4SHH3Uy
cLK6yhfHQ//dQYOZdREE0cSjeYWuQuuxQ5q8ko8LRwyilKxxf2ff+ksDYFZSHnhlgvvQcNFBf0b2
WEF570SmaKipM1SmA/5VNr4vIdaSLrTMA/fCjUJmTJW5xK4b/Qklk67BNbSO+n6U7l9b3EHA7OML
j8cBJrIa0Lw1EpswtU59dLhF58jULIsb3wZs1eVYr46yYWnzM7n84F2oAREWUXOzOhOXOSG9b6xv
SbSNW5lkwUrJ1OrrdxjMlDAIfStXvZcoj/K7xFlw4OL5gCeD2Z6LkQVfwOR3DQ1rEYwNI/FFVWaC
8pUOFGTPIqis0aBhtai2x9OiUckwzgkqqMC4B/1CcZsn+gapg/IUICey767Qmx2pvohOlHksTvhV
udGlNjDCpqgVodNrCGm7jBMH20EV4rtbq2klug3Kh+sBF35c3C4zrvubXlKoSm14tTgvhWzaHA1c
Ok8vHZRj9FBVn2z75l8gsLQgyz0hItv0Pri1o9jvX7B8bA3FaP+Kb9KF+lsITOmR6z3JJ6GjTleZ
wXpnd/gevSt9LdsTQqDI63yoekbL0LORZvnDEgoWG0X3ffq1IU9ONQunXIZd0hPzm9ny9X8CdHA/
Gd7LULalg9XCc53x6iNF5+AZL2E6SKHdG3fT4BScRyRZfS7VUZ0XYAZZM9YNMBbd9jDEMgal5ej8
JUPusFyrNPQvu3K6p/c+qYcSt7tY5Mnv/NAAe2VRxzMJC8jHqPomkPH7LazxOARsqo+vfVhkdNB7
lJ1I5zJR3qePp8rO86gYlkIeZg6iV1myIdhqrDtd5vsHDwEfvAvSAVhZrIc6veElWbMbYoN5nEkp
6CcHgSqGz8rjGqFCN4GJ4Gz/aISSz7CGVTvxTxsRI9uFo/6agxMZzvcYeaygxvAbzFJ2rMqRvD2Z
012A/MlyAqbGLmueF6/wnTjkVddcHbFW9Z7ttlGN6gf9VHHeFAlOnLAcG3qGfJFUaSDiQBnqbMbD
nPSpcj1GBLLmFA02EBqiDKWm54LG5tA7wk9l8rndSH+a68R+60fwVW/iI4vwkc5GUQe4baGcVaKm
VfSt+c9FVF1Txy/m6q1ZP64CIK1LQAXSXclRhnGRk3acqBKBSCkKk0unQspsV8AwkReqAfxMLb0d
c0yXRgO4hqW7XqX/RxTlE/rkfmVahJa2zfVXexK0XvspbwYbeAkZEYE0EOt10zuoecAHfiM3YjDm
QWZ+54PR05u9lVdBTZcBnhiCkHnGj9IIZ1o9/FWM79KnSrnirDkrMAZrdWcu22lV1K2QtyA7KYiF
5U+utdtMW6QZiyeH5s5pYr1xHTf98UsyvFyY28nm2xcCF0+HfipdadypmO4e0D0yxRBHIxlrtJHS
sYpfnqW6y01Ugjh29hlClwEf0Mj8gS1WQ++ZixvxN8khm1p0zx8TR+zaZdN62HaGxkwozZDLD5qw
d6nPRXt0Y69VaEeV4Cxawd4nxZVtNC56x0Wt0Nxs0t812To9xq7ha6qq4UCTMmej0KuhrVNF9lej
axUp0LsLpj58ZZhfFoPDiFXv2OMvgYyH6Ifphs8Fo4J9zex94C3TwGmu6OgKNQ5gSG5hF6uf3MO8
d2Rd956WnfS2TmfWK1CCCK4QD0imByYC3d4fa/RMEZSjql4BCCsDPwS0GFk0EbDUIWkSDQFoE2S6
TLqJGxVdMn1nLdFlTYBn7MZx8FX+Z413ATp1HHof+Yq9thgWUYSogsHXJlbibdLyzeNBryLn1v/7
wu0gppoW6o41SW02wdghnR4yLTB2xprVVGhLDEIjjaJOflsvTy9H6ByfpP8fJzco+DLQsdINv0wJ
GY4ItCpvr2m5wXcvzDT/TpMoetSsTgydYnKVnOlDR+tk+I6XBBIWSwgjzHXAIMabBUx8ae1yFFOw
+uIBfS7Y5o8JF/hYml7dV+/p5YJPpo80as4OTpMFN5W2Naehw320Pxu/30V+un5B57iiSkvdU4da
nNC8Fk+ilSo+hvMkqghAtK8MNuGydpay+lbWG5V5nnbnFjasZQRSX7GDdUFjGm0qnEFjHiYPfDYt
iSxTYkM3kpBY+PTt7lcpaLcVJ2v9ZlnbdroihxmvYiQNVf+b6d4HwxZEuXU2NJtr/ImuTBXW9ppc
miL3FjeoqNSwWOAPh93FTeMEFHXJ+GH4P/2rvJFJjgfkOLw/oS54nybjUe9gP9u86w4qqDsSnZxr
GswXfJ5nCPlEhOhg6v114PTJVIe3uQI4S/I2wa/k4axBcJU1I2MJINsIIDKxbrnVHLZWECEZphMl
1uCRL4JfCrw5zvisBYCiaEqCD6HRPicy/REy5OK1gDu+u1QL0HyzGGSSYk7CafMvCIXt8q76NRvp
7qf4hlw7yTg1Nl7FFJGZEPaWeH/bYp543h5TUZrBHjuix48xI6Py+XQYHXQxOfZawXU5kBpAhx9J
l7zJylZe572mthLat+CSUsf5Hbx42Dywg5KCNz9ixnWjy/ihEQ9SoYGkY02radasIfFjsPIPzOZn
w3ipaB07NpOrw/XVFpxWw82OVKZCbkuewein86SiYAvJmAphddwABl8gxh+qHTxBU1wqyLuKw/5w
32LR9oSQBcu2S7fUaTXFE32zmWjHgjtQ2VgjP7A6pPPttW80+seqj/USp26q9jrl8dQsFm4tcoT7
+BS3w0M0L7U/kZoW6g1uEr5YS2e7VjAIFgc5HuSGtLpr+TcA7sFFM+jEnmiev7xyiZWXf/wM6VUJ
36gRKSYpzrR2iYF5Xt+SPukoChGAHHnlQ+RPO0NP+kRrLDw/Kxae3T2GWBdjcQjhm8mcnvd6rYuG
tD7OpEZlEvyb6P1bJD63SjtSyYJIq6I1X2VV87kvb3Y7g90WyEGb9bAkreGOyiZ7DRYHj8QjIaEo
/7U1MoK9FT0fL+TLrtrfN/bcUUwI4rrplmmT+IFhKJb+KDjD2HXek3nDT1TBi4ZQXjmCDkpZPagh
1l8jpttE9hm1MoauNlSfxlJ7Oede/9LhDemZD5sndGXklrcj8RPE2vkJo0+h0fTijeK7ozQzqFk7
VCNj11sOnKpPiQXhi4vUs5iYO/ULd2fnq4oywt34Oa2T+iQih9NFSi1FrELx2TvMT/XQTmvJlIEg
7BvdDmPEHvwAweFX+OpE4hDSojXUBIgPJYS+xAaLEJ85RlS1dXwUEn9SFNLVoXqSJaJmead3bFHd
N3t3Uwl1Wd6z2MfXGeghYtviQSzc6Vn9DRGo8vQTOK6LgFpIIvLVh3vkiEHN233OQj80nymytxZM
bTwKWk8Y2uWGJFDcs0/aBeYrKO0t+qyCN237aQlV/xO7NKx9C0DRiqyVYDr+TfdXlTMlWPBTFVg5
R5RSQx88GP5x48OFWiC/SHAkf4EjkjDaDwJ7gwoRrsY69j8Z/grS8MnOkZuzEgL+Pp/x7yD7HN5Y
KK2emZfVOaIGt1fFeRmKns9C1Yor76onRUxshVR7I0l8pCrYaunOd7dCBbSdXAKiR374RKjwDknC
bilXwEO5UijqopwQYbXP8cwWDeQPElJa65i7J7g6X9+6sAh8VIaajKADXzSc/8agBfmoJlMyY9mj
ljm4taI8zWn9OC3xbu+YRz5Cq/tZaqxuQ3OarUXFbVhrSK6DYNYlyXFNVb6R9mBDfcenKlQZJc2r
hcdUCeVUd0Mh39e+thbsWL7ihCNBuMvjNanrCLR5mfXlYu6Rtj57k9mM2/iGOZlBjjMDrqr2FmHo
aeNd/ucdLXaKT+dQ0rt5IV28lwudWnaHX5uPIhtIbvb7XkbBqjYuzGCRjQ+Rvii5AMlxppfiXog3
KyZpyBcQ814s9DIF58flhPI1Ufa1hg/F7XwGpi/YeONNfEXZgsJ/8ZyfavXxUWtGvJZmhfoNLb7K
DDOAhr2j1KmdV+gHP9ZSE8QbLIHeKJ9LOwLIYidsgNGTCjrUHeYBZR1nknZklIj8B/QgkGB2bqWT
K4MwZAwjungRmIap33RF8IfdDVTKap2Yd+R7msKKWKXc2LLQxTACEn+WhSG3znl1bFMqhm/zLL3u
RSeGwwOil0g6CI0OCzPsEDua2Mb+xWU5Oeu19IqL1SUspPa8AJps81X2gyGIE8Ppew3JLRcdi5iX
R/AtY9u20qbK74ALZvAjcaytNerBr5BK2+Fm0sAKq0R2sObBus5+pPyaOLMFXG+8sZf3k2IMhnqD
9GhYCPdFpJjGIqie5ORXCqdThXarULTNqjo1ahLFQ4rNWKfx8zBArVRvs7JKlg4YaK7l0bwUqgjH
zV6eiClxt2Ce2cDkaYNVSfXW5ygDMiJU0W5doNFk2nkJUnYxen2EB14EBB5htEP45QQw3jEvSVwb
QJTCuXrjtPG2WryeT4CiX9xcEmLQnuTVLkozBOi1cdDDWYfPtNzSVGGMK7L0MrBwR4QJFODquS2c
vroDnYfZWyqDYuzy6gbNGOPki2KNIdtJDMvmzJMyAbfsi2uEOzf6AGhEVVaIeAOPqXljF5ZVZ8ts
KSirK/Xc9IHgH+BYomTjeAmR64l2A9ED6odB3nujg6CxECFrEQIqhLX2cKs38U9sV++cR6pEz3xh
O6Hv/wcaKwUkXdw0cDTWiVlBQG+ej6y9MZJhryJGnBKNHcKH2yL7baIaO1DqlN8ft3GEVRz8sg5n
aC5A25J09vtJl1QITmGXd5qs9R+fiEH2M36yOON9RoLfFrhucVjmDVsnyqw3t3bzBehDc4UMbWGl
4LXvrvlc9Ky6J1+N0uRzDikgzE4kC655VEr2eqdfK+IiBu7hUTWtqoXY3zC+aOVRIlMoNN+HU2B5
CCFqc4dsJ6wypjukS+0ZXtmQ7rCSBjVNQnSkJfpI2NoCfYUdmI34EFwb67KBriqiwX6761y9cLa8
e35wfZxcNxwiA7YnHMdL7BCmbeXbXbQpfCHyWmiqpKvxolb5CqH9hh9Y8o0HJb/tr9N9qlvpAsKq
T3e7ZC6uPYwlSdrgSY7ZrnBBaAausTDnW7h9HQy7/R8wIOHj2zNdMQ9EEx+ODggmRjymSL+E9N8T
D+CdpT94q05cEIdRD4BWYOnQm5W2zqQAq3wvPQisAB4QVf4N9J9mY/+D6vEB0slIdX9GGRDBn4zq
fMOqbgQU0Z7k/4ob3oY8JVO8CEALO9WR2DyqxYqgb0EenOZzUw6M5jwtuSVkNGrnmTxkEt3w7Xrb
9AN3UElAwaXNvRt2x0uLfiDdASeIPhPbtCzU72puHkJ/C9SnVkFunJddP2gZJ42q7meVdVapiXRt
7OrthK5SHiSDyP3cGvHgS+SZ8/rRiqjlSbhljVugaIJow5mY9pXAlxHbJKqdY7caH4rXtFg/eRZs
PRuV1+wp108Srk3PPu7d7d87JVFctGlkb9FnHwNRYDJsljskHQwkqVJwfkuCGR0pDxbZBypS/hbh
t4qgtEoZShtlFl70O9xaqtiv46unM0bvchRcWCyz3ZvBUeNk0Fr6dsR04UksTsE/zxgLN0P0p+es
SbgW6eUrQQBQ8lmHSVj7qUL9p2DhMAgvVBkjpZeeaQJb/2kAsphxH8kO3f4fTEUAX6QEjomc+099
9SWacizZR/OXbjoPFXYFeh0J9ry/Mq6FGezWaborE8PWvwOc20nCZmzBkkw1e8JwVyZnVxjXpkHT
i8A0pQ/NvES4gBe4ZIDA7UbL5Mt/4k45qXbkN9jjurQbJDnghSm/lROOasCauKcBwlYDcBtzGN5t
QCkQ7AsM8epjAYaoeqeX6rx+TL//n+pQCH3d2bx/AWDOA4i/Eb7JYAVVH4eJgHY6y5riP/ENroMO
Xvhi6FqqmrQ95GU+5KOCWMxQlgs8Nsv1SqTVZb5V+muHAyI+Y7jMn/k7PYegd5L5aW2LQndVY0EJ
BE1UmszYzs2+FUDw5A8aGey7mIvSwJKS1DBlQ2u0sLImD7/9Pbbj43qMWQ1V7WFGCAMUbJp6+Kvd
DPeNtzFydzxvtNEiC8bsGXXAz6OB8mDxCWTgMYiinaYOmsAvLKIIdG0jQG7ZsXwo9UGufKGBOfRW
M+4t3w3oY5dJ7uSTgFmzEwuHp9Rzu+nugmtK2mhnJQOFwytg3cc3jIKt+lJZnc5smjQGMCxWta8l
9ZchcCHjcuoG3qwOgvhzw5XcRJyJvhH6E7wouHc2f7sdgOVvoBDiGC9t1vHXJZoRckY6hvCXgSdd
17qwWsM27lEsFtfVE/yfBsqfR24fPRE7p2q7Flmyq27Ir+OTYbiLHnq0tZXwSxAfZujw7boANx4p
lPWjAqenk8/0mIyiG/azHndRMQuALkmnqJADRoIWRp8CNIvDW35aaocWsDNC2b+CBAQ04YZqpQPH
en4xB3btavM3yrof0qpD4+HPNQXOSCmtD/aPoPaUnqI9PdDLXJkteG6ubJJfIyT01HXDjIPUtOgP
Wn5pLEiQOJ6s56tDFC0Qif7nKVhPkFpNgfGmj69VHgyGDXUW8C4cHjRRKxk5/wwbVOAg+8DZcV+o
v+jI8PZ2htOlewtcW7qJmOvbgN8se4MwTczfHtXj1Rb/Sa/RuFpOlv71ahm1WzXY6QIgKBdGmiYw
HZ1W5U5NRoyhdGCOIGMN8HAkhYsuFtyYkgIuwKfDvUxFo+RD//MCC5drKBHSZn2WBjdgtafcnzJ8
6qE06mZUtnBw6Fdp0SixALCXINauP85+XRR+KQ8+FfNXwS8WCk5XFWeZDaDvMrZL0JW4DrEoqHGZ
X9rD26XzXjzH6h6C7FkUKhBnsMcXuHfvIcUno3wRnvimI2Q0cZ/Hgc5awEoWxE2iQCDrhYlhRSqR
vYbk3lbHU3XkqAIDwO6biu8iq6hkXUodpRX4igO894jxQvJYzDcfQU0OfFFjHpiHyvn/vdU8Q66y
uipNuK/TbzkBl5i80thbhKAYG5XS8QcGAgO3XyBZEed5aEJOO3Mf6oXQnjY/WQNZXjjX1f+N0BOj
S0iExOriSk8GVk/evYYqdUVySciw1x9FtLr1GFkmAkwYh2JLzRZw0QTsvUJZW7Bi+cP8mc7gNNJO
IiI0Eaxqsbb9YjW70HUKSRUeUpSxLp0PQvOSFx3awbMccXvtovAaJyb8ah7ccZU5GRHeEABZ1ho8
bR5antRGGCpL+40dYxLmt713sQqhFwKxLjKjUwSkj3FbHssJMk7nIF1ONi1cYloRU3Z9Oo1OL02D
3ApzdEWmeZVWMTZNkk5qkCbFCBKF5GE0WPb0PBauTH3uuh2KvTY1Q1G0fAFWJJZG2RwABsGCYJ1a
xdEBzDpDbbf+ygpI/B4UQpDm7/KWvzkz1V81uGKxEWSCLvapi8ATnH1WDzmYp4Z39FDI/h0jLDco
Yzk4rKhxqQ7UBe1ZAMIunXcasnbEH5X6Rc1mIcJV9BuwLaIChsQxK5z37E078IwuHo7DxF+quqVz
2ADbT/7YZIZDg73Rv0viiatc+uaOXJ1j9nzmrn/mvLi+VXsjYuwb4/3wo6M/x9nZQqMcxyt2s+6K
k9FFW+pM0Q3s0Irfpcm0ZtgU99XAy8KPHQogoY9Wzm0HCTqTp5B8G3z64JswCL6qPPrSnemcCajz
LEyuaQS5EFzIFw7Q4HFyp7YwVUVssmGOLK/n5MAhuz6QbgKWCjoiMDOF7bcTlumFtBzrYyVW0xnN
163SVeB4EDkFNs9VUrjjTlHYtOrvL+E5H6+tfuX36XYbjhruf0ATGPDzMTcWa+sDeSdJXMyaLMzB
/GFcj1eIbW8paGFUgtF1r7/2nJjzb82f9c1vXhikQbDWL9oRKy/wOCWVmC8BAs33Ati7gbWypfrR
6j4MfGOci1lCV9VuhJlanlgnx89VB7l4L1NKUvhL7UeMlvjeegiflUMq0RsPoVvHrAt796ghjLwk
nmn6rHu2SY7vsqKb3wouwgk8WDKJyzvXuHeDSHSFmeTHug/+rn6gbQ+YWzbawZc/iB7ox/iWCydL
5QMlL3R47ZTsI//2xj19cun8Vv3rI42x2pkSM7qeMKr9kV0LivFUqKun45Q2amsOJ3+bsaJRsq3s
0tfzRGgtXOKqkMM/uB2+/cXxCA83YywfptpcmtO62xIQ91JouCeMZrlr83Jc2vUC+wmQweZPd6hW
fcGPzAezYjjvuPkXw7jnBaFhK32G5nH+J1yFHQWdVFjuW5WPV1B5DpAanpbnrBubQf3QPT1tA6yE
itS5Bc5HqmiCJ3eLj6gRJHdfmkej4REv1+PtWgg/aXBiTAG91tAZH9Mno3DvcjXvBw9h3qtru4LG
6ZTCL6Gqr9IhPGkVZX9FmB1xoxCScIkUpFjZ0Zpwbt9HZmSiM/eoRxXkifHSeVD33y/ecMGn65Zv
XVCM0QV1oJOfr6nytHp/mMBiN6PO3KVfpuD0NqNXuLax6KWA4HhRxXi3C2TQhXZ3vE7iKeHEgbji
3dS/v3Uz6pBn/oC44rRRMIk5yKwkVe9G6HfD+nUDSlsHZEuhH7NQJsabs8G4Sa8UgIDuZmOZNgCi
uWYcV8W8CxqXhYlAeq3g4vaj5zndTVzjARHJrZJem18oLnVM+4sWyNLiF95IKwCXkmcyayXgsK1v
m2hXnYKk4owL5vtFTDwYxl45gEhTw7e16Q+KTACESZiS0jbXvS+vqTeN501yYzvDdexLVHq48ct5
nh4R4HhLf9nmECBjuLZYleCZzq97uLCt02ZpGGKMAFfwXyiObxjouYC8TgOSjsMRzvk8dOJXCP8O
8xxkdp3cQ27uAokmqeRt/zsGx0+nJpPPgR1N/vKkedJQnk6w4yrmEpndHC5Y7xBSS8tu3WxUquFd
XOHUWeOCMw8Xxwbv9Dul5TZUxOhsWu4xfSWQk6l0aXkHISV7k4JSgWM4RiMsI5v3Twt+wubgXbZ1
Io7ukLtbPi5HYJkOe67p2GqhZ7Ly28Lnw6daMjRZyrwrL5FCupctkGjIX9BNcsh7H43SvfTZmU8X
VMVKofjUqCeqQqJKxV82yZc499L8KWW6h1amNR03pQF0uy+ZH7zGqUnhp6cnVOGrizOuqfaMGA3y
TMoaDKet9I27D769TVPj4c4k7pLxVmdxkFfpjyvWYbDhVAZvVN5aFQ18k+Bv34dFDse1b54pX0SF
qYInMY4QWjoo0pVLh3LoiR/VsgQVP2TIDuIsG9UvFGBV2q1HUeTbv5ZF6n2Q0IUVoYWj52YB/myb
Ihv0UBeqZdzeC1TWugImnJYoGkpcf4trYT+ETjig8CgtCBjOoj5LMJUOzK/I4C1Ee6UIVJFHirrU
UUY1KxUSHkbFaTTTbwL4dMgidDqNV/7rGAtxHRJxVpHYqiuW6FoJ9MWZ2i0iOh1tVHagu4J4z9Mf
VpnnikMgYiIrVlLmZBhTu/qTuRI8CRwjckRkXd29EJeN7/qZkG9CGuUON6l7nRMa+65ykFeQ5xre
fALbVMw5bXmyMHq3nmNc2JprIpCzT2PBTlyrXLnRRWfZGrgCaIfLvwtWW09rhLfLWQ2ecmIw0Cb6
KQwgIBwxw60EPfrlzR00ByBvuA7a2Bzt7a16XJwgwMBcj/nI8yAzgT3+LRebJo2HXySRwZxYEoXt
PmIP/c3MqmtKw72qpNekO0cT2vAfLwks3vgVSG8jc+XxcTODjBYi9N5AXptMAG2gYF8f4tIPCCiG
X8iJJYD7mUUE39aXfoQmbT6ZzU/nyVLaKjsQVsdLGup4O1QeOWGPhQQuoqw24QumM1uX+QQU7THF
d1uPRMC/mJi9EhnxtK3trYggV+WQug7OldJaoLYYUlDkQSzxHZIZTKjV+J+KzKFaWNVIuAJIsHLn
pWTM786PQYlYQPDMNmpPYtA+z1KtpYw0fKUa+UIlR+rO3H2csE+BWkC7ramU3/T45ECLqJ4hXItd
J8SbhFph+97yQnThhryyaYUr6EmSrdHjoB4KDBa2DbwuOfYuhhic4bGj+WPJP4yfYJLxkxdGCs5Y
KB1l+6buAN2tnjLps5Sn3oAJASlPTpjMA3kQdJuWvfx7f5PRtTaKqGgSm+y1/HkeiIQFLqjJbhHA
SpvSVjAAf8UgVlu0LzugRIjQndt9sxHvP7wG2Jh1o4+b4mXgAVk6LNpWh4abefIjDghaSsOlTuqH
USSkYt9mjoUgjV0Ij4D0qEcaSLh5KcYX6TwUeaQ4CcbxhUlUhibDGyzUAbWOxBX9zSgk2rIxZac5
KZ7I8eXqVbhSsQdWoNSCcysV/6eViAEvxKSKi4yMAqBWBv5AzmAdSvw7a9GJsScR6sQnpDO8P+Vb
Z76HIOR+iQp0YcCiD2Ay+47RV62RwRIKal6lgnZ6z4hJoGnc1lznHzNN0+xFZ0n5bxzpZUcnMhyu
s0rvb0e5yLZ9WrdTzTSDPmeSjjhWfYcH2fN8AjBxsyys4fE+WM68CNgyIVwYQqBgEpb1Y36R2Nk9
nrQYc4as1a95QimtM0LTcqP0CRtwwdBgAjFi6FbDb2vGp/hxeIuJ78wz1UYrWbkLy8oIy3YjsM0a
bNgQlvqfg9PSm2s2dP0MWaQzWKeKmoE6/vwqBmZQSh3BCkS/Ht7tPl8dL9WKNetguDtiAMgbJcVF
CFJSDn0a7FGERpI/E7BGBr1fBZXRhudnFlvvQbAE1KK5G5xWt0KmkaujuxxLJ5KFg1RR1/miBxM0
3Y2I5ab3xeToFWf33mkkRnNm0MSlsXVRNtM2gB84eVkzDp+GnP31JJlq/KIalQGEKIeS+i5XCsAL
/3DeIWnyPhZY6SzRmh1Hhis1vFXRSnEodXKlIF5spLL73ZbXUvjz3Q9EMb4cg+4aSGkS4cz8WTK4
XtIobOOdx+n5GLQu79PjdeHll36SP6OTLMusfhpNuSfBAk+tE9OdVOeCQOkDRkRHFwre2kutLrnH
MGn8cLEUdwIIUKs6ajf0vcjbt4QiqhEtl4ZVT+pGDszwA5oUjU/AauM/wTCFk3sQ+9wNQB6Bn1Xy
HQDpgjbMhRO36hDCm7rTNUvLAWtAawVZQtCzoik1K4nTxjvhmYj8PNd5U5QS/RHLyYndinztqnGU
5vcFEoJ/C2EUXMs5xtrZjMiZDei/GqXJIuBtRozfyucVCHNajN9KLIzGe01Iuh8Rd8jZiepbWSQB
wFgsYUwTJS21t106uMS9xop6o0x6Yz1MgGba/lWKLrrlJN6w0Rf9FPMQZx4F+VjsskQTll73+cQ3
Da/pq2ZdvhfNotUuIIQmKDYMlGMfe8PB4vMVBJfLxKuqCkrkxVdwPGrgp6fUvLT7n6+4tKNvgJQc
X3yV24RIeTtVTlNeb0S5xyxJV4oGkyuoyG7xGQdGgyeyYz7W3bfDnMif+naeL9Uehdhi9qfDBVHs
gso2zXFfnQRe8YDynhPmn04uT6tPrn9BQKmovuDWyd/alX4sdDTFsPtAX5ENqbImqMRlgyFb0FX2
uFfQzbGVqqzdX/mIbgnnyijdIf2KX+XAiH6ZJ8ml/9RRfQpTnixOIZqcadZT2QH28Uplaw8aAeMT
gUIVYtTISFT8Ukp0yNhwEO9heXUyVXxV+rO/+cRRaRKDhGbytuL7dK53gUs0dC4H4rDLBqpDPNBd
MvwUnOvbWZM3MQChtAaeujgha5Psiik6KXXhb0eNpXDjokMUMRQfM0rRDLArzCj537ymDZHxAzN9
jyHQjOpz3mHuIVpRzMpyf4GZiWYbHn0WR+uNSx5VTg9v0q8jcP093wFRutVafxoZr1yrBzynjdTR
54n67JK09Ifs0YBuTVAU/0p7U7OWs4odheYW7wjms3AQbmkwmbpXin/JielBK8aFCHmNqqG4yvwS
Lj5wPR4A5uA0fP+Sck3DEgC6vHUofP/pagM+sTOSPGbuYIm4H9B3Mb4BS3+QJYshtkyDQBXAIowG
CA+qq8VWOQY7eN5zSc4EtR8TffJzcQG8VJkMaTQDw5Y/Gny7XqZpIRwkLD3VskWR/d/tC4ZMAsbC
P4U4sqWpM4VHjfFdVsv30j6mcjsw7OmCevjEMHmadTkPJ9cNu52Y2uP+U3vJTKf2oqy2YaFw6hT0
/nRtmZFBD/oiQwwnhtoYcht86c4Fu9E/gMO3El6cWLcRn6jiTOHO3ig0LN+NTmdWaQmSzciNgmIP
Xdg3H4I0jbkYGLRdpW2NhsGPUPdax18UZKP+EN5XkJ53YG9pqR8sEV4sfZnVtN0Z3zXG36GXrpJH
nJ8xWwR2zKhUQuU7ZQioSLPtIYkJvQgXnC0YnimV8teRfRuBturA85P8wrTklgjjUXUH8fkYJxDb
JC7N8J79Tuvj4hjH6BaZVA9WsRC39tJt+AsNb9ETn5KT+/Gdwsiqw9XXS6ICPr2yJtXtCF41rLnr
Tn5OYuT3cyKXr7g5sBSSCQ6Fh+P0SZWwNKittTi9f6rlNQ+R420QiTP90PmlK/StF7kXWY8XQ6hJ
1MphSnajGtlUJReS9zCr4dqU14W5kVfTxqcTYMQ8TzvW1BOQA9eqADKPKLK+CGNG8OzVtXWW064v
OhCE3t/Jl9NJt9XnWx/GA0Te7IurAm6Ds0wyrtDNa92HgoJbLOmvMP2XEexdDVYcc/3WyZPnVYHf
jUU5vIPPjQjh4ItH8azC3ZWyFGUKNq0TKuf5fmFkJEsBa6lXxlfpsHdBuZTOU6LewO6QOqh38eFO
oLASQiXUZJhgLhH0mrEob36ymKB59bTZuTqja0VkZAP9mU1WCivkYE5mcQ8YtUGCyEY2xlZuGVNF
cLrg2WGnPG2sCzCm7JU7aLJOh6AXHPj/0K36TuMq1OLRcohE0lqP/n87jGzZiOeuGi31AJ9d2R3Q
rSWx9DJrd2mr6bkuKDeZeE0bRm/mKF4nKjtI9kjzeLe0WYOfcVX2/KJ2z4UK6PUxr3G07iJc4OB8
9CAoBdsX1EI1rfcUfneDHH8XNPJxbqkwxMVN9Lz0/oIf6Nbz2YHt8mW6WRWwsEIxM8VOaJ8Hu6tO
JyFl2564oWtrJ+mIntkEbmTu2BGCGX3ggteUiMzL00BjlS0rzRiFx9Tn/S2D7JXLMmB6Tkin7whP
Q98M4wdV/SjSObhKl036Goqre1spRlw+xaqQjZtIFD92Swl9GciMU0icLP9LMuYzHzMTyHGqumFQ
kDiE73d5gNjmbMgK71Qd10qh5dFrf1RAM4GiFGTW88EOiEcC6T4v2vjdLCX1mX9SBDjGVglRxdOv
C4fP1Yh5W0O2hOaKn6h+Nd6ETobj4mxhD3Xugc5Ly2bbgIXNXZLw6tus+KIVkESTZa4ADcD5NwXr
vLFg6LGY6BaOfkd3MTmU7GOJJ95n5s6gKnsaPzhnngKIDVEeYTQ8pmgcWFCQZgSkn0eQcdrmxAEj
fTzzqReffxOZIXrTqUiQSLZIuKd8ZGhP1YcXish2uWPyiRt2Z/sJkIyisr7VfmDR8y7TsFyptI5Q
Y5EumkLVBBTT773tKeShqi4wGrGSQaUgrLyC6x3OfD8kUuShhYAptA0qzbmnyRiFDqkypw7DX0yr
+koOALjFnJ94u9y2ebDQecoVnygxAwqGJm8phItVkphAPnM3+9QbPsCgR154gxfEQ9R1BvgBj4Dh
35JaLQz2H+s4tye9uRU3mLRachsviQzglmmGlG2DYAc2rNgU1vTHKQ/kSQVvtmI+jrYt/OW/yDDV
arAcVKjI0pYwEqQiZIdAkd4T7HtkMqeMQLukqcfdXIHu9N050+3xkFFBwbgAvm1MJ2SsHXMoPicg
dyqw3GyfYUc8YC59gm0RppbfAaZkehMy5BkN2+vNb+tZDDcsNKJiXjkSWfNr1ENYjt2IzT5dDGVL
gOVU7i1eDQ+3jGWjQckVaNkqoe14gblxcgL5Gqzs/L13/ZDFBTk2XkFYU18pVTjRfLIn4cHpf6YD
UscEWa9MMXhpWjGXxn3CuWKp+DT8aJtR0IzvUVmbYagQEpKTmMY26B59BnbLIFJs55GDGdvL09ML
zmeoy3qNzxApHJzJU1ZYQxXzh+yhRBK5e0IQbWiOsETY7Qip90vZI1YvKVbp4ej3nhUq2t7Ns/OQ
L3USsMA1+ul7hu+dZfwnTlqtjzZHZUtpmLqvmjgfKeKpXjjhs54q1yYUhO1eTIDvPmHpb9XkJ8yY
o9ca6LJ6sG7NOB0H2sklruifSYKdCCG4HQtscOaENireT48cNiTpMgbEFU9qHpEqWXNZ19m2bhyS
wqfc0e8znJASR8/I76+yJBNnJkFMq63f7Rb+UlVqzNBUlIyADYpQ/jA8AcmFR2jhYIuH7hoxV8fT
lIKMMmwzDNVpe8+remMiyxs/x/6qMpSodkAKM6eye+pXbU/SLUseSM9oASOnB8cEbYxoQ7NJGTK5
eAkKWDtbAlUrtA7CHJY8XELGuJIq/Xfge6Vz/FDuFdl216V23HSq+Xpp6J5FtN8p33Uoefuz+WA0
4Q8JW1hGMUJg6fR1pR+YZO/AyKeoHuSTN6hw8Pi1AmyODWCNzedixCG5lYJ7XHQEUnWByOQOQBqM
1vnuKqtVM9ep9jFSOg6jkE9+IdmyPNZyWIz9zFJWyQ9VkubtBNjFFxtOGZTOd5O5rpCw2zLox6tA
SDSKtXLkDDJP3+/lizTyiFDj47cENx4rAa9XElonpht3yAqsNwH3oVL76TnCE0yCpujloUqG9JMb
ewB8xbzcBuxU+JIgtm2Y/5y6COHRbUoAfgorY+xjS6NSxiN5hPzhOmkXEw2+Iu3FcJlKQhd0AngT
hetLgZ570zAeIFD5amwFzlqNOvkLdcRiIQAiqGE1eD1Lk/ro3yp7zvJ+b2h9f7NPulr1wJM0MxAy
MbXwqmuqz0TCDuQ+FneXJSESCNQ9l65x7ntsqQ03sKjyqj75Q5epqA51/4LmFg5BQeIhypaFEiyN
zh+tDZOvQKEyoOoPteaXWFrDAMdgRQ2nGJXS5qX6rjur57lNQZ/kDs/BjOOjt9WBYqDoOL7jFYPt
LK8ny/yoG71kOid5OzcFaSyUvw6XS2Ntf0VdwGQY3096Vg5YCEsIGYMAKAZQ2SipowycIK2OYsgC
H9KaPVSXSO5nh2nK4hmaCFogiBsmx3MEi9tRhUVmzyG3TZOydRwlXL6Xg7F2E+h+4E4VBbPDDkTX
WdhQ+gj5CQ7oAkkhVwozrzh/jSXdxUKviCKy9L2Ru1T5wBQnleeTWM5yyNJZIJ7nsvHKo7aD1iHE
mCFudei9WSAOzW46ky55Er1nYO4lwxI1/fa8oicIJeOajBPcGr58qHTG3mXuCGmLBiE1/U+Qk6Hv
RHyaXkhYRCSCaag1TOZu/vnnse8eNqCF3booHhHXsksxz//WoAwoD3y9iWQe0H1lSewZtEFdRvAy
//fxN7T5n0gJ8EV7DBMz0Ce1vGtysoz8xxyXkWrC6zCVj9anRibbmu+8mhgjMlN0y/utdmywJLG8
qh38cfBv3aSPtrzIQFdVCQEV6cTJl+vgv1LkV/zu+L/QAE7XDxtSc+pzKcUEGe6csRgHT8H2r+QO
Y9A/AQEA92kmDKXrqGFCC+NL9vfwf/LtjfV+AQoJCyhKBczv+Eqn0DAIgOBnJWcDon/k+l1dKoAO
xxG9bicJDD/ko2LC+aWs0rtBLr+7+YIgAK8pkxUl2SKSfFOPvuzVA1YYVfr8FOKqeiBqkJrzpIzl
bqIq25fB3puRvRq8xiaDDv3kto73zXmd0tb6LtdElv8dqRspndklOx4snVaHzNbO/nWdPBN5gbUB
7U3rOM1KKxazupJO0tFy53GPl2/721YlkF844SLA7TyzJmmoOxHmI1wSxFSNDdP+vMVI16IYZT51
JHSykVJRD+w3pXhXAWiayo6uxxMEX7U3LnbN/ThfIgOPFajwt7zX7ilfus1EMzHq5XMxijOZLvc9
jBeJMImWLPvZp7XdMUFngcqsBVFB+r/wyI8SCLXfdD8o5Z5929wlwzNrQI0HTvFK/9YNmC91pmtx
D+uzNJ9EzRRC/jI9Nwegh8E5iPJHazGgsgnWZy1n0GFNCgw4h7ntniLQL7Csvxv374p+3CVN5Wj1
jFH/dUMNvXt/e3Mug+o02whUl/zJ1lqKvT+QXPilBZcNZr5kJLciysv5a8YewbG6ebQwfstWhpHo
QieQ21saAsgirCNNn37+eGqR9j1DSNjhCrn3ktk2Zwft1GCBm6tpK4Y7H7DZGiJuEhnTHKJZXp/d
b5c4uR179lCeYM5C3JRkE5mkYF+ccrduhOh7nB49nQuqqdB7EsipsAGgY2/cCG6Srnx8RwG+hcxO
XfrmDuBhI0vCB7j3phOCdKe2UFSDBIhivlQP5r1tEiSqE828tTIoED/IAcErxqRyzg3scb939oXj
wULBtkLfCdPpzi42w/LauUL8mvwAchW49LBIcf1HKs7EOWttIupXARXDxS7QzclLrLWWJrCHIbbD
ByuKNOi9TP6QSzMTFVZrHFNBTIXmUZFdkaWUVz6uzuqb/j+Bm8nLb4wvs1DBn/30huSbGt4Kal9u
KIqzNCaIeSqzmoEJjisqgyrrK+4EibcrEgC0zH4UxJ5cbmgIsH+0f499FtXZM6uV7CuYAOw8yBzf
jKP7EvctJhTkspMctYAyHh0JbtbwWFFxo5G7fBJ4psoaqHsmiUpPPXJ1daC+OylJ4N4rWPwKFNHs
juf7eeNdDgXNA3UBMVnJ5rPW21I+fQX1P77Yg0K1wDfRqs0jMzjwjlVRS4S0oWzXV3iHOPMyFM9S
cnQWlH2pcazFMpqN2ZnLdNqrx371400FdJAP2yHArAWo1OGMmYrKvoLVq+n+33Dx4OpQhMqZeSwA
qlE2e/N9nBkQxzmfEmHNkTFRjEzcSenQZZ8K4GyZd47zW3wcsIspxuDJAQ4N9zJ9T2DG+cgOMSEd
dTvNToC36AJxjDf4Nn3kJTSZn3U30mBoac1QSiA/ut2SSUIGkVx4nXWPvNpFntjW7FeVVov9qaGM
SAsU+qjimQcFgSChcYE6Ij0er2vRTA6WRMhkDJUaimhFae0H+N2D/F5oQhULiMzMd9lG93P843+F
WmIh7XCVzITTMCHcvlbGZLD1JXlajAoa68yO2RcEAd+NMOYe5IfWV6bL2egt68wI5sKGZUi3sOBz
tU39iL+Oxxu1/vJKwQmgotqi4wElIUwvyJY2B/cjG8MUtFq7FmHZC0ZE+svIq6R+vA8/JAxCUbZE
PYGuA8Q/KwdMeQiV2Yuds6FNkX4IUtRmrQTZk5ElHWDxPDEwZWVHK7eQUXqiJ1nn3biztpONTu+p
AtRGsHl7r0PoiNBW3rEluvZDcXlplN62CNhd8v7KniJYuMLDoy6E2JbxleqbONixEHIRI3tAGOYt
wqiaj3f6QHIOo+UrrOC8nRc3niOkqzXZ+Ozx0HfSh5hf60KnPn5S3Rz9e8Rx48h0xn47sTEguaag
3IO5MH2dYGj27tNqltuAHNE7M/WcgsiwfWCFVivUOHD9zgIjVL4BwwZJpUgxlqQB/F0s/VA2l7gI
k3SltUgRQsYJ69aIBsamYAJR9r2BKKXnK6w7eeJ02D55vMS47OD9R/GHCe86p5xfG7NtsCX3zUyz
H2QHygvxdUNe42jr5Fcvwpt5HanFCDvU394W4JPiNNT/GyJMDVCfTKDHhx4Tgr456k4FKM23eg87
TsFIbnY3lDqzeXb1dfSGllGHDCXIhyhSf+pnpbCXTRZvmthRKwiLjIrTGgMTTlgcRnGeAWtQCOkV
ZhgzEEpAeAh7AzuynKEc+D6LSXhAnesKRJtwPnDFLmGBfIzxpZLaZ+AwxGVWJrn+s2yvfmA1rFZG
Z2kfCloYE89eWoXyebDz+EBiRbXuvaABov842JvaRBQjlkkaAw9aU7y/Ki9GeKPfufqyI7JITZiD
GoFlIfrTr4V11F6FgeGb6mA9CQ8A8N3C/08giqJvYIHVXT6gCzy1/20Wt8b3V6DRCpvkfo9gH+v5
uPL08f7pzMrkNZXif3Zw3zQlITzDrQZ+g+t+0B23l//S7YZZ2qPnvGVfsMRKXzP/UfnDigpiwRkq
yomSGcapModk652+yzhkIVsoKN1R4kzEUvo1/4a45Ul8PRkKSjHbCFM3j95veNFYS27XWHvtU/HX
A2tItbxGX1c3gd59KkIKsKT1nyZ8FYKXm4yOfjRoXsjkeyS5fQvG+WnRcZ8aIyDiJnTobm8y+cdj
IspEK+VSKq4Yv01sbsAMv7zAPlPUP/Q8rCNVykEpOKEl7ZAan9eGnwlK12A30H1wPgoxwlIHYF+k
Nl2A/7nG1btpZrStJGktItY2HCj5/EU1hYSDK6nXBH0J6yarV4aVFGGc3LnDMdjTyRyut0ID1y7J
Q3UbnjDK3fuAz99s7GkVUFTXdB7bheLBPJJZWG9l4v1fQIcJQECtWgLivU/73206/8FZGr6RTXIW
0NZgikh3G74pgaf/jKcVfN6sYv1nh46KOEONESHay3qWuD/o4oW9iHrKjldlmG+pPYd4rJOQsfqL
F44Tog8Uqee71vF0hD+iT+wfX6jduFku8L/v3uMHpFGCl5agBhkTaIWp4W2NVtjAIxsJZwQU3RDv
yXYSQtb4Ux0eaRYIAHHxt9eBaW0GQB9vtSfPkDK2GJgrgGDap6L167XRJWN/6Y+KUfUGEDp2inGj
eBYsTKUFvYVkhkHiQ91DrGSpY95UIiozkc6PAsAp0mXvWt7cTQ5s6Bxp6Tlcp7dwnF7jG+you37A
/eHvqpZsAf/LqSJCws/fAs3eFphW2lUwO+eP8jzWZzKz6zvsiYwY3tvPzkBDiA+ZYW3GpP3urH8T
4cxUhcu8UAsfPI5BUA15QIe09DXtVapxd/VbBKDSG+M6mVeiWA67Vzmf5GEGu/wSkwzyPx4c7Aqc
pP5xAs7EOX0lHXOu2KY4byYF/KgJWZwccaTx8lRxJmJbBfjUXe/plpGmQMtnCmoVHEJ2NDjjwVdg
2D2np9JYcIZwdBX+Abo+GjJ+ysKmScs9Pw9lOplyrHNOJoX8B/BHYugTxXPLzSVZVNoPPOzebVMt
2P+TgVpMepclQzWo1I7yj/8bi9AyyhIJppJW91+ztM2IIWWJA7mJe9Qbm1aTcMS3MdijnAxPBXaH
72CZhW5tk8InSlyWkbyRxl8a/oM1AJNcvvjVdLZFfBv0HTkNYpTUVF6/Qcpytb8WE2GZ/274oIaJ
sIr82fO6iA2PnCdzQENYJWWDqCydBbDLT0PkFlfqxEJS1MR8ymVeA46cC+xN9qT5Rei+pgNRniWw
Y+w/Un+ECZN9pCpFRlXaMSj2orkrJm9yl5ceXYbeU45Cibxa1bSHZK0qF7KLTo1HiOQJoiUhRpS3
eW/bNDpgNgyryxpQcyDGQhpOTkEbCNh+RL6OVu60MB+1kdenITYa1J4u2wxDBF6NF4oU/ED2vDfB
S5jYtFPDdcUpYgFUlgkV4ImA/Y9Y2Ty/rn5Kc2fZNrv2nnWTwUJUAks8kC/Em5mczegVgBKid7CW
mmOuj6ranad/U3GkdKNdGVseTT/NvRRuBRfe0F/leXwDxLPO5kStjwya5a/BeivIiU3DR9PNF4Li
t4nIJXk+B+Bhh3pEkCyBvqhEEED4GdxwnGsuroLE75bQIBOk/nGzUDCGdH+e7QCkRZ7FL70SqIxO
wRDj1Yt1awi/d5hr5jLIg9wyiTISZ49nc+Ki8HUYrrXvdU/RwHvEqNgvo/1sJRgfG/VGUGRJh6Ri
aN2SRNlsbBTFYX5sBgUyX4sCvy0HsZHn3IdESlQmmqjEuhSBsB1ccynGb6DueAWzjrTqzxaZsxza
xpPxuFQuL1NTf0xlXP4trRgxjupbm6qjCCOjXOjuA6ouE+tv8ZEGuaWbPFT/yw7LSdwhqj+oN/Mm
DVrxW7UKuPJpnCwKRciIn5vFMs+awnAgjqwXQM6KWVVgxh6IOrKM6KxirdzKUgkOa85ih42MvgaJ
GTjyed890yN/mh4lbt7/LLUpOYNi/eaXNVeTYkOXsTKnDlxarfVLo6NyTSoChmce+s7l+DFczCFk
BQi/mN0+yB9/R8lpx2oQhXaDCLB9g08DpolMvzDU38uXGCsGortlgeiFSBATU9gB5s9ZvEoecRNe
sofNSAgGHeZqh5A/H+42cUONeeq/2pHORApoi2g1Oo/97OCHjOm4cEmDQzzB+ZKyeiOjlxJPUV4l
I3Jsn/0Ih2pDh106KuQ6hvE4iqMNLQG9hiHKMbGcdXrXunxpJfE/qe23EcII7eS1cvhpPTFOE6sy
nDivd5B4dmawEbXSPFKf83IQKzO4HWnvTLBqmG58Sr+dweV3W1ujoNCk5YyES1q947G4Qh9J0Laa
3gbt4PKeP88TTg7ZXlwX7JXYObYezdPFCdlcMe5gl53oQgzTHS++teXCEdyQI9nrs+a3MOmycXTq
0SHNjm3H6DJhn1g6W5XqcvON48JtVXtIa1xp7gnqrtcx8VqQdHUGUdXXKhNyL3ZM1WLJy35FvIVt
SbYWk5rv0bYfXoxFoMibPaAvTVe+4EXaRT81vsfZQpyphhCxV/zTzbHv4WiMkSAfU2Kcusz7bC+a
835iCusWC7epntzP2rcyDO8TNrjEmKhrFwke245F9y1XDR3lVBhZQ3Ie5/43rYcAyR9fq3ECVHTj
yqbRAVwhTfFP8v0rc3vtDj98iJSRT2ieAuonsOrUu4el9bYsGdOE3pX7AVvBEpMdqJAGOPYGYc1+
fbk15aH6MqCCwE0+KqNRHRkgWYp+wzS+i5gQj84cirIM24Moxw4BTkdC/pj4c1zN/a4LekteWy3u
JlzpSDpds8QmhO/Ds48RX1pMxT7qvWvWSddc658yL0i90roO8849HCC3VQcmLQ6o64x9ep1aYbEB
vJGI5KgvyA/NBAfK+jM+aSuGGvLbKjUgCZ33I7Ct8+JlB/4mZp3QJJXCHGCRU13RkQV+AVDtUK07
tO/bnnz4gUqyIk+YQKEt5tBLZcSkE7Ae4xPXQya4Ly6Xf5CKSyHHrC4/Nnl46uL4fRt7ZKdFs/L7
bboJWBwpQt1+7nwHRp7SDjoOJhyZaOFh9d9uwUNZtanen5wSzjJyjC//4k9WcXZbPfqwQB1xc6ms
vHf/gvy948379VqjWXrlk5ojGi8MV/y5epn/iqPMnRg48oXcJHJbe89hu3G1io00vQ6x/zrndL7i
dbI+tNmSz/gJeXyPdKTKX0vZB4Zgp2COT/SZjWiNhatfUU0FDx2qKqMV+9R3uwL5P9Iz+6CUMeiE
jGyOZ4ax9dFpp2rz85T3QtsX0vsHyAhFoqMPmBS//yb8qzOgfQjRrBKsBhX6z5NhKwslD1JiCM7m
+JCabCBd/vUIh/A/GcOyP5kWqg/L4I1yKsQ7K8XkgYRsHLkgJ8CgqQuv4ZSB/B/oX/oJdlWa+DWU
iD/v81mUDFOtk4ZQ5cSVCvlhzXIB+vzdE0XwdXuPprC+czvB+blNBvs6eZTydS34/EFXNpe7F0LU
IaGfoMkYkdvqQYCpsgx5uutsfErVTB4KPP+H3B/I1hvznE1/7pVNoIoExSB6HENOr6vu4o9R2INV
IBIprJxDIguT1UQqwjl3W6LEivJpqfEEp3RfHPXK5khnyc3xNsh6f6zaELzwq+Gr5yhi6uJfxOO6
+iDiWi0wds68UvyiuuENdWWd69W0rHoVLVfHMSg7g/VxdELTqPHGFUnKfivWltrxudqV0eRS7ZSd
W+eVQQd9tc7Ebi84/iqVorYDvfrMeezvTfUcEZp+0nRWDEtCvypZWIbgnyN6fAHQzHXnO4qBBsF0
bqdV5x1KXTVkFrOfDkXCNilSloT2fEB+hjMBFmH6OJIWgKxQrzSAqjTKfuC5/BE+pL9ErzmKh4LN
D67ktAq8Rp7R7bxVNqMjkPuHnEb1jIIBfVa5N3k8IQgKmegZhFwgJe1LMNIBGgxpfr9lpUeYv4hm
LtaqtGTrEpllppw0YoGrQBWbhEj3tgbCdaCew5m5HS4nzkhrxxzEZF1AUS0wjs9rdy203qi0bkRU
Gi+SZfP3Cz+NPI4e/TTuLU36mcO4gywn9NSeI0YkgV9iKZrArFcPEokKcNFr3IUq3KCUxHDo/pGz
nrmUXmeDB9iskOqlKBBn/SxILKXET0STQOLjwWNxlajnaBb3Crj48bP1cYHQ6GCK9Z8TCsFYPkVj
ATbQnFvRKfNGlyYyYVK38F7DMnQXUqg7ptL36Zp9FBIL5BXYrd58rxcLLpdmXup0BzPLgeWa0keJ
ud8JFJljtVj5/DPLGQ3kFfU+YIRTX46Xcjc0HH7clcruk+LN3/4VhOENZ/wVr6P8aWvgFdNVNE1v
l1GdFvaQ/4rMr9eTLohis9GxsEygYrSpqSbwVJMwN2YWCh/nf2LIUD0AZehsD0pIFIhbBUtvdboU
a8tSBUM74w4z+hIB3ys4UpDrCKt9Sjl7iBqJg83mPSMDgifnfX2iJ0Sa4hAFc1uKMor1PWxiG+A6
74oSZ2Dl0hHFlTnPCM2fEfJBCk13eHMx/VWoRqpg/VCP7gqEedoFtuHU/HkBLpklPC8pkCY+AsKh
NrZT8wFwPwwVv6dgLKvDJIBbyx98CC95iQ+PtyOwnAqNqSCiKfz7CEUECMzRJebuHp70//9eF47v
1S9XfEWxy2xL1WNy64sUFthZbCcN/AvI3AiOvJfbMJDyXwwrrKdAnaf6dcxgm+rtO+6DY9JrkU3g
876NfGB+S3aYsKovDRPk/KbCwhplkj1EBRN0VT6Muj7dt3KR7kP1anWoKgI2UYEmvs4HVMITE8bA
RtiOs2YRuFmVrYbYLkcUk4eGNw6YG9vwIbbWB/LIW8miygSxBw5lO264sLzQvTQCnm1pMt/+FvGc
Yv1l54LswmlYfyL88NEsqRAa0JQlblD4hFxU+af7bWo2ZldFxd8Xb1Ml7KlIyFcrE/cUqCdlIvLF
7m88OgDEPWyMWERnReYG3U9TTBBVRWq+jdBl7oDbXB8zSAl8zgJUOhBKPp4pC5vRTKkv7+anDbVU
Dyur9NYgjJy+4M+VZli649ix7wjp26dKyu52quThqEUm7VyaG72TNLdfQxtug6659RqOkW/JQ4FE
px+/t/kdUQx/9HA+1rxPFSkH7Osw/O3/nCBFoTAHjhKmNKjRpqGTHc1e0k1nQJPLqcUgX5Tpnuan
szBwUHsi57RZPZJHvZoGmWknSfYyUNS8ksQQWkTW+LqU410OldygywwbIX9khXNCDSv6fFLBV9xL
FRyER1ZMPFr8xPZvbw9Ydno2w86u4W/RWRS8r5v4uKj3Wm7p+SoLVa1FU3rlj3oauKYAAu3Y3Mh3
yk0ymlv71LdTGp+jko8Jteg4wEHK6pRb6VqsxiU33cMdvFJD0KBH6hTYEvKmBfIq8cxyMJyDPKbx
fRguceEM/OoxNpf7VYmf6x2L8ZLlESZGf3pOm/mOIFtXbCeu0xZZz/lvd9eb10nNUBedokOZEEdp
aTwedqywX50kpMijjQGkAXZipjpmLYsypF+//gcGJt3D1CasVC7avStADtFnWRsBcKSPZUvoBFDg
GHJTquNJXQsJOR1XMf+g/7qTAOaG0fXBXMcH0fBByT/8uDWXYNMhEwoFsrAuCHAwM45qlgA+QtJV
KbFL8qgr9xxJqOhdE5AF2BMeTyNrAYxQaXS5qZZpdPRV1S+niGIAl/xoHLLCKSst2gkm1Nxx5XDp
3llZ8/eOWdwl2CKu3JB7PCi+DJkGaYdwhmwpZCXeNZvjcFYK1z7MmzzFOvhPudrQgRfKswo43J51
tOClu9hIK/d4BLI20uoRBRIixYT1nsnyDHp2q3S2s/A0Vz59vW7jweok9q8dp9s6LWLTXSphf5fU
xkJuwyTQPUMS9D8NC6eh9ia+O8a+4V8ovHXZRExAQYPVeIjO9NxzIoTZYK/PzU6fqp3q793kG4UE
Wmo45muEyVDp65/OuKy23scSOUkVoCJzwHOIKK6iTzmRdtmhmNL/ug/IpzpH9T1bjluSM4eJNq+r
obQQcpMuRqHspLej+qdxupMbAqgTdTzFuA27yC37yB+uyjjnd/lO/cm8QS8K/D7x5uQtAKQlCgcj
kNKLWG6JI2MBXjr2VqEndDDzhhjvEybSSTCVKSJImLpLn1ojNCVAhCxoEPgYL0sx6ik5w4e9mK5y
pOQvS3Je4Vdan2Koz19+2rd2DenA+qF9YmtyN4Li2wt0FVODBjsuqi1APF4MB54s/mEvhO49f+XE
RGH6yS1nwtZRGZYY+UflQ+DH14B5dg1ZA3QMXLc8hC6Yzk9SBfK9N0k2YT71E/qcmnBFR1j3VcGq
YMQQgB/RYysYNfRb8xUzuQNyx3b6+jkuQCCfwRNXORijm+mlz6ENDpgJ/z0smfDyESKCYPu1tx5q
A7PO+COvwYS5mL23V/S/N7VnX3RdY/wjjxENWjqMNl81mhKjWCOcI7LB5sX5V4kS0zQ4Qk+BocOA
bydjqtMvTeVPssFb9QQQTfBRB90ONcuRjeqHJq1iFNUULXoelgWEnmPTPXXVaZeg/Kx6Jre9mxRU
x5H9YFNxawiuY6sWjL8rRcGxAAORLiz1kLZ4z2mWZbfAbGFbLtMJ56m5XJ8J2Z7ubatCiGzG0TDp
YHZ2C2SQJW6qRm8OQlbwp86zqjhSJumINo6EYB2hy2J/kPJ5mkrvVaRddxmr3XyhX0sG8VTj11lD
dUBC4gHouqyRP8oFwOdCMDYI/bNk2wCdEAcjlYfiMZ5MHZTbFvEojrfb7R8xz4NDWWnqUb45OqRJ
I2o4zfwMz6HkLWoTvbjdE4Ma6xlIS/ZM3KBHUWfO6ldSPcv2zR6bbEF6feUDXF6E01soruwCLsWH
rdWv9l7a+qyLYpc66hOmtsmbbskHJaGF/2euSdURk2O0y9YXEZHMCY433Du2BWAw82Ty6oQUFU9l
wzVsWWa8jxkAOF7y5e0yg4TRhZKO2hIptOyburlvkeXwljxHEUvus5L5IqbtVS6OSopQ+2AqhEqB
bbjYjnRTIrlr/Cp+m1WPXZR9idHmq72hMSs5uNbbhIFwhevdCIZoN4w8ps5X7GE5xdp+3hp0++ys
8w4J31DmjZCpp6eRs+JBRiBt8M5lUhg5ddcRKnelm8DptQq8mdbLdmIeajDclp+B9nWYXEzEnG9l
qNEnucYW1EwoEn5+q3bno7tq3vpuDuGpMLAa9P861d56SGAnv0pYAIl9PK+uN6DqazQGHH/u2UY/
7+PbKqcGiVg4paZpBErom7GyhdQa1XjkrWexQEIvU/JE0jyS5/7ZyMuFpXwirlYEpKxAV/33bcCo
imDK7n+qj+pcso7pAoC9m90r0TP9E1/Xa6qMXDSojsE5Z87hTDaoCLRx45NrsODeCPCfCwgjGDvi
8KxgoNjLUxDcGk2Ogfh1S+sFJOyUxOTsVw5Vp1gPkmo652I2lhXiwseuSZlHbmIYTYUNZ/kqcOuU
kGtl1AGW1wbwF225P/UyXck1zkW1V8PkiBxNn7f1/RxnxRgDxsbCl5KzdCoFFsgVpdNnd1Xd2aPy
wr8zCtRGQdk8FiE52c9zvCCqsTA22mXMykyX/1/nuuII2zawC6+bLes14Oac3nk4nOrULk+d4IGb
bsuTbgJ5G9iMs6LX4UGZweqYC9N3z1pc4KX/JsMsv62muhk96rP6eUQK0/MzNo3vI4YQ74Ro/rPh
mHEqq5yJ2qXJiLwmhFGa/C2M5jieHDdlochHgUYSYDZT5m4t2tfegHSxlbh48W250ayPHDxvtWIA
gYcr0354PV7nvBtEfYMd9i6jfnnuSkEnSgEwrmASE8kc461M/5e6XLL1xRBr6E+wt85kAAt0jyyc
Mg98d++3zErMyJetTkfSkx36GhkxQDpyZWKVFjjOj86rZ/pNAtFxZgBM/oUfDGNCXsiSkzln4Ici
d7LOQ7+Vjnsgepmwt12BG2Z3WFYECSZgPaQlKLGNPJa0Hd00rXdxW/Iio/81+tNDB3UJ5zkXG55B
z4+voXBjo+QTte2L+DlDxc8iJd5HBxFhUrTq6hUkT7DpE9W0dxHzMSigbFAsHj4BxgnRxM8MvHN3
3S6/u2X7YCUifNXs/g8s0lMFHz6MBjjth7oWO/ZP+lFQNO6JyPs4W2d2zrn887LMrbRtpMLMT7qF
JjIh/GGxLv2W/LYJZoL99+f6Ki1N8u9WWhQiI3nUL/CjwY/SF3jSo0Kd2AB+Dy08iEjhSZDyD2vC
2MJT3eX3Kbp2cfd7L2M3AmKtJM61y6uz1P5ovBGjF6sGzh4ksjb2JJ7J7mx/NHg9W77LMuTRZx0P
fPZug+vxfg5wQi6oF86J/3ayLfsrDqfFS/+IltCLrVw1WpGiNbEDIpsA6UN4x5hfPcupT6zfmwMa
VvYqvzSgYrfxwB9q3hZ1wo3nNitO45BXK47C0E2Y+j5B+paCQhvg2YchbpFuReFW8Qu727Q31ouL
x9vNiIhYubHcFo8fGmTw5uXT9hvLHnGLC7hJuv2geC1lAaRUo6EGmxWGeX+lFjn3ThWmyume3GeJ
mzjtJuaVbje61nDft2pHIVAdf/E27xmThdMngbSyyVw8WYEcPlOTRzLtB96aHteF5rXNPcl4FmGQ
Nih5LBk6VtEnS+3Bs8PaHwjVyVoYv71nGJopY5woHjZbv/9+dpYjx+XBkjA7nCwrJtSJmH18uKF4
CzxTiKR1ZLtKXBgrE0DSs1ZxusM2YxwpGcFWjkH+vBPavWnMCBkmul/jUGu9jLJlsowKR+9MbRor
56XCSacoeeGowM7rAOGB1asdTCD/5Dut9fRMGDupsT+aueBhMRdN7dExdXbxLZk1nBTj5jS+ndAx
3LPWul2zf605r7vh8YSwL+4LmWTF1U+vTMvb1Dy6QMbdz0N9tTNPG4j4MEB1q/jtmbdPWGA6TwUj
4HFA7C4t3GeM7G8eSV5EBTQZX5wlucf8pCjkUv9hA4TUVfoOylZwYxg41Ag9sDabHIU/yKC5vx9J
dcUAmYaVRf4PteTc/vOBRqQsKPkgzLg/X2+psrjX5xJ8o7qZUruY2uVbLZKb+VfEe2DmQ8T8/6Gl
00tTE04KM22e/nXICixNy43aW1Cxeu4J7Mzfnz4xKMftNIQY+HDQOf2DguEYqQo/4hY29PvP7bOc
qKH9ukwrJHLtESIq5ChQBE9awD0QLn2ZaNJSmJJVOY3V37HSvY+/a4rN4VfGSieDmLw6lmLP41hf
HPEC/NupTLY3i0zm12QQBMykuv7yQ8RRv/LG0+/+piky9G/PKwT33b67f1ZxhAfddwyfttPWzj06
vl87xVzkgr7KdIgS7CNGLBPxMJrrvFb+39n3pv9Pd5KJx4Xp+KukJ9Iau+FVJHSsDgPFdwR9+pnJ
pZfeoThmOp5D0dlZjLJuPPwQJ0LNIzQ4tSKnf0J8cyxPMvXcEIPUJTJecvQezdH/DAtQRhx2Ffbt
aGfv0XjN8VSsICYpFDyOgbpSC1FdAx8tNiWgHVkSfXDbit6mfU0ivpg9Dgemg7z0k8le8iflnO+3
qehbkJ1qTcQ0l9Ve0tyHadMS+NZoLQO4h9vLy9WxhYDDFThCubJ1rXgFf3IKlXty9pbEvuZer8Nt
s81ZkbIlB1QdTI5d+gPtDO5/FJkyno+Rs+A3eqKwcu/tBSvtbsk63iEJCTuYYsXcB+RvsumOYhWb
MuVmgRTH7t3bvhfVi6qtg83xcN48dLX+Nr6+09HuKFyaijqsXvAgdQyE5ou1rkJJDxXkGUB2PD9J
LMrfdiwDsJY1LIgNUIf1W2Z9ctmGCe9XJD+2heVM1PGrgGV+lPA6EC8k4FSHXyQgW51Adfu/VBRv
PBIZkPBZ+ACw+gSjgkx36dQVK24AOQwDjK3CBoTvk/JkSFuVlqiv4ibb1KE1a1ZuuLNdS4tGLo8j
L9govRRJ6drF6/FkUyj/iaw6MOm0us192iryltZoXVZ3jTZhuyuooAsjRV+UpqqoiGRqqGh5dx3j
lYpqLI3yM38SElPr8KKTlxxUyVaNxqbHQHvESh+6IG2SjwIdhVFyogJOesZ1/RLy1RcNpBOYy4AZ
IBLxFk/wMJWQc+Oy3rda4xgzrbehLI5nsQjFcoVQQWgkFajNTirwzNmQmEHGVW7WWQLiZh4fauyu
RkAdPFR8CfJHidiGVC8vwUsz2e55t1DXW97Us3PJVAjrzT2nHcpiqN0mzPCR6DpALUGWzeFaONME
n1MOqUty4oyKK8T7vKvdDymXC5JyDKgny9n/RxCwNDm1jeQ6c8JGiWHJ/v0n94U9+7tP1p3CC3WQ
e4kVMU693iBM5ZpigyI6BjOxljtAiBjDd8+Y4svPfiSyUbhvstS2dgeduPM28uAqgJlZEUDhmpGl
z9+kglqoYQ/2ByPdAOZhUyC4ezyjzpKBnh/jK/h/vUFnGfxFr1Ojzkrc33lnBC8/ANypjPny8fDF
eshY2l4woMhGIC/R8iE3RydpdksmlbszmCyM0/Abvd5A6pEB+uTGBsnumUXOXvvg4gcCutz0s0Jh
JQuSdvqLLVt1FURzJQrsodN/DWskNRkCjx+d9y6enxVztPc1mlhzJOZ5FnZHm34nZqvF0tdU4ARn
CSMJfDIt647IruKY454ZcgULFCFLgYjKQKBdVMlmZHRdpvfBUky9D/hhBNLTaowWp9XT2GlFz0g3
eOGcmAy138+OSiockpocxFI5hf9CEl9k10UuHJAr7NRORJxEcEckWMbwrpFuMwTAJOMk4/W9MkDS
ROEpRBM6Pz6t8gcQzGOxkUQWoq8lXz5ymEfLQ7wBQtHeGHF5juot+hr28gw5IZZSY0crDLjItb2H
dzLmuvgFvxdwTNXWRpfLTaqgrqyh8Oh17f3E51XUG+MFtXjnSTXrjzKLJAwTIgjYeyL6BRWX8HRh
QMShefN6PjfMB/Sb1lip4nd6zySEK7VeiLe65f0S1FPdArARVc73OMjdZk+J0AOiXeCqNBBF4h93
Vf+PfGFvLWEqV1buHSE60UEQAnnYaspogg97P9qG/J5rAdOisEfG5xuCEF0qZ/Wj6GojpSp0glAm
V23wKr1RMFph8Go6RLfvFcob6cSH+ePFQdYpOd/Kt52fNgh7JIhayli4UkLj7pqRCYZx6vhpmh8B
xmRz15tBGa2jQ/NgKUUlTtiq8uImCPOHTBJXAy+Xs9SOBcklL30RTArD7rMEjhLSfnFs/nVnvBNM
4mq/ocwYDCtY7KJLHg2al9GcafXhE3MDjHuAb+6K0D7sfP5SEdfU9yRPDe05zKnShx2BKoeVT1EQ
LlAhSGwnPzlpQ01rrxFjcNZ2t6TYi7NAZCSP0GoUt/R1AMwIhH25pp9SvTZNN1/+RXrsR49r6GTp
4cSHWGDT659vw8uZ2DPaxfUUfmh4Ms+tY4BbtsqnfJ3AWcT5FnpYxZFXTImfs8KSXBCW6a8FIGe6
eZ6fjcCIeTQf/fLllOqLBSqIqqqtDldXVNYnDCBtN/2dXabsgxX0XDt31BPQwY77HK3/dxnwhT0r
7zXlxqkXNxfN0k03Us1AJRRE/z3DpEUjOZyWxAH9aCX+wMss+6rEQQ05cZD/jgxdGJ5RCpeeppPM
CV4euR2KMX1xCR0mcfrMrW6a0XMI96oPmfYzJV6N7ecMBl5oSLcK00Xy+TbjAiaLPuhwAHo/NMcA
+wVizc7EYlNfzVBstMMZhgt/DWPZlr6cHNW1C+t6zVySsjubFWyP01LL9BuuiDPZoJ0wRlAOeMgD
wtcatNTQUzM6B9dOshKsGxaw4XlfGBcbElKY1fQYLchAtQ66Y+guKqEWqTIEnU2a2MZaeYWKv4zZ
/SOt3u7eTIkKINqO9D/s+6vHitXR2QTtVtOQNR9qOY2z7Fd2DC3XmQTIGnaBP6ifoX9GftulWw1z
B1jzujJN6qwvC6Hb6O3HedWxLDXKuaVE6LYLzLN8cKD19D903e9stTY3p7tS1jsHhp4748bAg3DA
62Ky43PbFFT2ZPOqouvWQDuE1qhs9PrG/QH0mz2aDXXN0v7Kt5GniqsxH4ah3TaSlzg9r+2F/6fN
7vussknUkMvs/mZfeEw9Be93e/eR1YLDpxT9VbSk6nA5EWgHrAs4vGapTmeXlNZnm5mdRHYlSDMO
HAU9FA7+r9eV8+DgNtacXUxwRQSMxPyjQ9XohgXo29Rf57zijlzJDbUXjedh2eqooFfl+SfC2j3J
JCeGUm/9QHxvKPa4oXgr4uG/df+1Len29Vq9efrpWvAtK9f8B4dGBxvp4i0OymodZVqWfB4LjiXm
BiwlkrFksLiqAWkUYBVXOTb25QllXzzo3K4CUFt8KX+SfasKxGL8haM5r4UIDdNcbdY5oJHnkUJx
CQf20hVtHibVn6EwMqt8AayYAC98MdY71M2pSf+6RTzaalxozbe4dB6XoN8EpFEi/xlISPudEBi0
TvnSpAXagfzqsK4QXpa1/VBG6Zczpfx6D0t7gqRgz1z3Qi5dMq3lHAHL5WPmX32Avb4Y9pTyUJTl
PDeIYibuhV5bvzO0lZMTtL11TDRWj4xWi89O7vvKk+e/j+c4gclBBjohd+9NUMYWtr8weSy1dxL2
HKkpTwMcbKKc/NUDlQASTmDL9z9r+MYR4ChBctQRFMupMwPGUDJdoOnEBrs4ZWSd+TfGwv9qbq04
u3MiLNQaM71I9e6ZLThKnrSaVXCD4hulB3Yd4y+tde/7x0a6r2TXHdKBbe7BdMw3DHIEA6HRlBw8
y3qZQyTEbfbaKyxGYzHJzsDs8v7sSeTPwVYNL1fKKZVHtx2m/QA1mvqLFCQmTOCdFt5FEkYA8aCQ
VzIHi9Vs9iL/sjLkxjBtAL7nDyOU645w3zPXhLc3fXl9No2UXZv9kzB26duHtUTYmWz/5cBmcVbV
h1mT1VnA1XGxZy7mQ3wNe/35TNeFanouiOYnPAR5b+ShIkpTGg2kBEiPtWcCHwdjfeNis0XsnCdA
zfbdFomYaz+/HdLGX4j0Jr8vV9FxdhIXio5BG4LohMARJYkUGPOUGs3p1V5ov7cI1u7ek2WFQGNM
rCLHaEZlWCB8tr9e3jllLAFmiYW26M5gETaANYtvUKRUoE7YOS4ICClKFd1GpGUq1bgiGKqlKqFc
jSL7Wn8PD3RhgSi9OmoRICQqD5J43UTr7vWAy1Zbo0zgHSOw+vTDEgM68LtFZEqOyI3KtyqaRXg7
K/OZtqpqJzOX/YTgKQxoBhkxkx09irkSg9AcYjxsX5OASH+eYKuGe3b9SxF0Gvpd2LqQan+KwbEU
HEfjze+/PFIY0Jf8JDxp6MpwvQpy/JLRHFXFlRQBU5+xk7f7X6mWg86ixVEqCuzYd0Mf/6EDrz5N
rpcYjicCW9UPA8jaQWUkmbmCdiOXf+m1UVFsODibVxEjZdUxzmlVd59itrH0MvmCG0Qn4lzb8SnD
NQD+QFWaiZ2TBp5W0E68r0cIVmqnWIEqlgZ30HLajg48O0JICIdwuO2GyXN7KNyrL3os59baTJPL
Rmot8b7Xa8jeCOSrKRcX+TXkRjSmeQoJsmYgl2pfXE6tkvLHmlkA6Auooy6DSFNXoGbMNJIx7vqF
jGzWa6Qo5nyHt7XV3Iu+5P9yGzQcOTmDrPYdk84du+coKQM4zf76iWRt5e0ljVHap4BAfUPjq/QL
7aVOUvMY8FjbfCyAGM73OheF/qm+3H3QFyqwRp84CpWRCCYxiwzys8JCOpH1Wjo+gXZ9x9GpuTwE
pQw2dX0/fU6tSRkgQAXJuzDfRnMDxxo1NJowm/EjCZQWRZxGUGTEpW3U9792gYMNbQEsOq8GqFmE
FtU5s74yqaMIpVyEJQbgFzMPUfdfzXGVSvuKWhUfhwfLA2mTGykFhGLHMe7ZZnj4+wmVFiprCmnQ
2u1WrR4L3hh7NlLeiMZ52xF5Jm/pkzipbi0JhP+yUMG8qlbECJKhOmZslyaHNIT5BzB1cqjDOai+
NYdbj/JYHAVF8xvUs7Tgsltgr6ahb68BJeemBBEYsN3istQ4572mEJ37MYXRbdisCBtFntKZOXu3
v/t6DegvhL4deSYR8gJTyj8Aqck5G2GWh/vSbTpaB5OTqcqFcNqrpmsAWokRRmK1gPlQ/5ZZ6pFA
e9os2YMF4ahSfwVZKylrj37kwOkeO4/5OKzX8I9M60YH+c+hAnMnL1/WkLAIotIeoP7dB2nZUq9V
nzDjY//jxr+A8mPU1Yh0zO+tH8WdoaSVlcCVN0wR35g+QGKJibHDD/sb7j0PrugvJZpyxJGL/IKt
rs5XU7x1r00U3vSIaLy0TnAFoQ6Da0nk/Lo9i7Qc1AsH8UQmEcduiflgaBolgkIahi7851/9BK7U
5lrmM0G4o7ZoCa5XKP4VwjsAYiUgaJ9CH8Nyl8gEtciArqFnJ4ljqOB42Ndz+r7ZuZFBvPZUPzGT
Mqy5XfvJnGRYVF78HBgB1k7rqi1RWLNMIgxJvJeQz7jc/3RlQL2ZOCno7KaXQT/ZYYq3jRf/TnYR
NO8PfqUWZKwayeuHCEXfxNdp/1VSExfwuo8PiRBOLYTvlX6oQSnVRGXdiAe0o1weqC04RUmYTkBu
rD7flQxJwN1q/PTiK9bGtJ0Mtf4xB78PD1ICvTAyDoXE/2LP29NfusrvxXZUZCqwuIPFyh4H/THJ
pTRhEWrnsbUL96Rrdl6w7KleQVu6xrwh5WdUJ58kY9avvdpoObp+ljF9eMzUz7E+4BXllnuDYSpp
Rqio7xMpI9reymOKRU+C9jvQRWWZIx5vhe1+jEO2T3OGWN3a7Xyxkk05RdIwzpvz3E4WbFi9cCoZ
x/nGgGfFE7WkT9315vWiOkjP3nD50eAoyZQbknQwT2D0Sep7bEiqqrlVc/bMAjkv+UTTBnUx3E/4
HXUzAAkmA4qA5lhCUR0Fz5KeWcWwZRB2Y0OAGL1NzCWfpfRhrCEF8MDXbVH0NEEtDWwssE84SWse
wI3AWWNrMs6jPxv1/2ssGp+st35cZq0nxjSHDnwJsC0CZI9g4xzG4EOVyRWbWDSk0UgpnzrhPZYz
9yUjC4Y4sKHn6Jg8D7fxXXK8xb5HJF6hGS4O/eVpiWcnwo61P68v6v/e1455LE1WLfSaFUmbi14r
JYeIND7XaLXyukMfaaUAIbcDMIQCrJb7zjj0lc0AikSUMf97SUCX95WyhG0V/IVPAd7eVW+qsT3/
ADA58Bc2ZpoorIF+WXgLgssK785OOZjLSINeoNcoVbv8j+5IwBvbI/7F0d9UbpzGEoLPvDdhgG6T
HTvSenxF8GfR6hWe+huZT+xgmUQkQpaTXxxbpNyBbOQ6F/snzqMIIgw8UZNH4UxzfOgQdPv2CHp1
sEYKrxQxlYJVJWvXFVx4+iW70iazCgioMMzicbBiEQKaMebGbTBiy7a7Jxz8Ix+7RQv1b6GssMC7
eDoVsuyO1n23zSW7urW81hcYua1m33GkbMQbhXWD/0eyjGdCndPBlxl1pfr5dLVPllST/QNsPAyP
PNhiwZRv10MJE7TUup3foghw5+B5tYybvOYV6b4WYIcHOk5IRPal/FtJAmYblRENX1FjGUi0wGJt
gr1R9imrM950L+8il/utTUhJwZ0FLtEPUWOEwfvyuQixyWZUGvEIpN88taMspgcKEvbHOGvH8umz
x99NyAA11aEGRMWGZKU7lEHTMkQpiu2I7AiV3VCL9RQ1FYFqVP/tczeK9HJiS1WyYQjBmuemtCS3
zEpnJkpTLAF+ltDBn0i27SFoKr0vwJJyU7R0q2+RQ/90Gw4FIHvakpz/7ylCVam558fyqF2042+T
Jf95DJQ9Qw3PbdH2ABuPg1lyfxrOsk3Ph7y4mqlD0acMW4VfXD/aw0mmZYkGdYnj7TIHUiByyygq
xPbkJ6xmnBCRf5BdGBxa7AXUTZZJEK7yiNNskvYjXRuJsUY9zY1eXVQC5OEuiGzDd63dbYS08Qax
zgSAeT/Esx6/E8TWMPsYgDf2VB62V0F+NNKRCa956ZGW6XmZVNKtRteeJbeZKKrzX/gCb+cE1jsI
lJe3JphLQPtPDFPbQ2c688TpOK2u2NEASyrmNZIZzt2U2qk+4Iu0BGj3Qu/pfQV7azVSOTkuYUwh
m0dK7KTk8c/OQxfJHYqrtqJ4K/5Z8N65GcWYd+IEl1YqNvy7nTbdyJTeBsHYQG2IgWZJ984BVwKF
6G3tw92T+IAcxOvb9EIzolbpU7y7pEszmuPbT9aISW+1Q0xGajfsZc6Qi0Sfm3Nn6sVLpXbcYZvf
vNxLvSpXzikXB+PATvlCL2Wj9yapcyyu/6BXcsZyHLlWvz2DoXvUCLEbF9rS5kubIkMEBtVCYo60
pwJwUJAI5qZkhhWhcKYGsV978X1qwA+yxEZdIsWdqRoIcHDaV2upV2xWu+A6iE+siS1JdtK5ssbY
eRGv+uESG/WbYqOhPP59DpOQ/j45iJkL/966eUM/iQPsRPccPQnI+Z1kRnCDLluX1RF4mJ7c6wGb
G0RYs995l6sD1A5DMeKNGmIYfpNm18UA3+USpTcJTxj76ioCakQM4+FguuadWYBGRW8spCMWUKmq
VJHIsZ91FjmcmJREWxa741o0RLwm90G5AWbuISiVSwNeo+dVvwQq3YoE2rOZ2mgwpKxKSo/T7rHR
JEcBAjTMHRgES2zp37SwK/z8hyQzE8dGxCq7cGAYaPjlMoFsyXSN9ZXnTfTPiQ854k+++ZZHkhbj
hQ2O0waRG1YJ52ah2KprUZIIyUM9vh1GVZyOWQwNpac4HxOlLWDjqhHMU/Ah7cpjfC8lJE2dUCbI
T6hWUZd52PiyqHkMcpBEHtDgLgkEuv3Zwm+DCDKLLzZX8G27P98urpeiw0up9aRPH5oLif219IyS
f3GKiRMEiI2GjerdMkREjErI9JqvyOn/fddtcy/w3jA/fQc00vZuPTrTTIn8bEvoml70SVRD6RUR
8dh+O3ZZ7d+xO7rl66n0l+s1Rzc19cvkAYhf4paVGRuVVHGvbVA8gmL+L4BMRUul4dExrPzTIonp
qryfhBK+aWND2jr3/vUyxInWc4CMEFJN/G9SXHB2dsZzIb3REGuRslr+WU7L44XOd8NkzXERClNh
/bZjmFuCKiwzPCiz9f42cm83vxSItPUneHF30C3MGTu5n45svUFpsNyjFvAzUEBhKYqxp67rzzbv
uYa63KfkT9tkQeu3v8m80Ce2DmD0IT3t5SZun2v1yaZ/Rif1vO/hM0HSR3mJtlopL2lec23pgxtv
dZKxpSwwPJIFzfCdH4an6oiaf4F6Wx8g2XBQZTO7sP8/ZrVZ6O3uqCtq7+Bism+07Ry5pylw3FZ0
csYjA4tKa9CdQEDXaHr/jOjMKDXtNJwVkaD4UZb1z/7UWGlrdACFeYaDlXo5vSzPE6r9A0Uh7If4
66QIeJ8Dq/cb9bg84HACJ+D2BgNIfkK4oRAe6LOKt+5xBxTE+1puSslatxhKz/VPPNncfiBu3fCv
puKRxKcPU6w3qY+CjDMsuKJ0Kpa34BQJD0xriTl61P7e69tXt3HnQ7KGmqgCu0mzLmltoIF571s7
sD9HGKWy4fAqQnyqdLwYyJmIoY5NU5RXuExITHA6er7VHJa/0Jwaobol1DDOELpxjZg1PFZdnzM3
FYisSpkZ4f+ywrcGc+hI7t65ou+mapPQ+os0nfSM9xg/NRn0KqRXEetX/1E2YHzpLfP7s5K962l5
UsHX2RurNyAoVmWRVSZFFgQuZ+rwfjeGo69RPbgKDftvsgkp80tD7V+3N0oJpT4JZKox6IAx1cS1
i7DueXy1b2IF7XqGztoj9S66cpqYURz048PDwnrnD11DUQSJjYcTw1yNdaHjBXt3Tv723ArtVVAq
aSfkDfL1F4oE1zN/1Y1xpbESU2mbx25BvB9IStTcpDhanERh4naFdX1m8qxeGoFAqpnpElAYL1vx
IzKBrYBtlqpYmzEiFXSAxY3YXZQlZC4Lbk1HtxBPBhcUCwTSk0Elem/x4Nwx8KgIY6g+Zsuy69n2
RqY8YBYx/tKHI5aSZB+/exdUyToXSBfCj705RYPxWAoKdL8T6wsKWpAwizntJ6BWNEs5izj91URZ
dBaL776iNanDeoFTnM0txMlscCO7nzvOTZgdUrv2fP5+cO77By81HcHrTLeHrdbMl5yTQYLyR11u
tpRjuHTwmQeYkYj61pIC+OCbsTmnfO1gv5/buzlJMuuX/HfJpem2CT//n2S4pc/NyP0YqJgbHls2
KBTXUvLjntsiM8LDGPtxF+Xc2j6rkwU0rLDWHwvD93b7UvGFe05hKPs5Yl88PUzQLklA9tMaihA/
ZJGrNl/BtM947mj7UaIAzuMySAgeCQOX9Uqwjx7g3MzZhwgcWU8MYZtadFTSPuau0bFUFYg1IbE5
QHrBxowEusKmDycjhBdWQ6uTieNcnXAztYD8U8MY2TAu+ggvdpfVIPsweUTdZFmazPPvxnzHy+Dq
80wnGO9LCvSk0AkDJ7K0XvDVIe4Q1rmEwXBodHJFFN7gkzpWuHZiYRZI9ZAnS3gSlcPk3PJ5PJHt
XqDbFHPbDpDbPgjB62tUr+BYBXlemvQpwQ4Cm2y4y3+hHLF2RDOKxlqNMEo1H5wGSHmkuyEZK2ec
hx5ot+HXH3DeZV4OytBBlXu3YBaYb1FbkOUHtS7wn7tBuifBGAzYmLA2gx/qCUD/b0+kyEcOZDH8
eM7rgrcxe7mWLyLJIBkx+/s0PpyA08cClgIjONmNpmGmRIDJCzf2HF6gEsQbpT9Ot+hcXcDzJgp3
10MAMQN7jxE9GUasZ4EXpGdFXtsWmfOt1+o9kKMJanh/hc0S1s1q4rS61Xqt/9SvRARGqiGOfbwL
qhPCv2YdqrqBmMLRGD3Qz0TX0VATW7uYtDYKZ7bgP4kdXJBGfup7q720NS6zlkWXI+vMc5EL31ry
ceuci6OsnThSmUllUy2UX3x3jj4OENVvTdHPenaW2ymB9O5QX01FNMDIT1K71c0Gfc13zWkyRcbw
teeRCtZFG7hqyGaDM79tE/kqgRauTfwDZs+i8+z5NPZckvNOSHTg3O8p5WUAwr6Sy2LCThVlTwYj
mcDk3rvnfi7rdtaXfvl2A/KLLe+5WmfIPINZZwYefz2XCTHY/DbDQlTvEpeU0wi2aVnzaOOu4VeM
ECoOtFGhn75Q7Jhk3UZ/zweWrEfPZKywzwcMDIECe/BXctCb6JPAPxTW1PD6bg9BeSljmVSgVbKO
k1tyBqx0uyTDO/u0pKap1Rf6jnqsN6JO0I0RWN3BZD8OixJEeaBJwPsPq8rQyfI+xh9x2s9TXjsD
TN5IgREWk1vBMN6cNSfaQTMpphY8nC7GOsUZ9iOz5xaeskoXQ4bt6gmMjE1ywwwYVf8nplpVR+nD
6naa6xfovbGXBWssc7sf3XB+c8WtOXHehNaDZut69lIv8NbTRw7ueucD/WwqVi8MKx0F2t1d8xhs
7Ed7dj2AF96oBLkNW/T0nozADJYNfu9/kqBgaSSiJf2hg3GA0yUiGWbpVMf4SkOHH/BLTNKlfrVj
ZvbDlAv9NC+tffog8jahvzRq96KGVc6yYor0YhaE5UGAF0v0bJhqmwGjP/geSSJkFNKPzkhTAp9l
N8y4GpS3WKB7ilsn7IoQ1JrRjCiXqwcCXTrk+Q1uC5S6ULXON+HxnAWM34+Fr+ThYRniP/1urq5l
xC9JSh/JMN07lc1FhsDRWLYucP10OvjLrJY3C/RnRk3dSlAKAbAe3esP/8U13LCW1apst98YNT+w
heCBFlrZ1puQkQQ2qllaOF1q6YhUnAdlnAPSBuX8eWdqcYCRO8n9heN7csFd+/UqC7c589l/KABB
n8cKd1CjwrD7PakbFObtJE9C5rL5MUOjVfwzSHG797E2aXrGA5ZRgSq+e5zwg1nblepH8exZ/fFA
O9XY7uiWpXV6zMDpinZ22JDMPCb5k2GWYGdifPo/5l9esyO7WRdNlrn+lyJDGIUWq1UweP6NosvE
pL6Q6DlU4xc1YHiN6N1MX6ffbV+T4Dw65e5S+QkzZtLOvJwWcF5k42bfQnBubuWZ7mUPoA9+DhFB
PVXeUIWIlL19TRnUzo82cBYUjL0croDiEzej6umwtKLsIlwHaH78r/EwFvzaUltzDl1dYCR1EAFF
q6Ljpm10g7DReyICF0T7SLHvpQl3v7/DzDcZ/5WIK8DNA0BcIMHW4+mhmqJTGtTSaTiC1sUW9Q8N
fkpGZIZSSmzCJl0fAG1CuXkwRRLfMaWtX0mfDmMWeV1entSJ+aC/r3PIo3ZrnB0rdvzxpY8UUURR
lqmix2/AfAXzXfT52n4dASDKhSZTRnKB2RIIxfLlU7TDd+klDvuSKGUlkHy0KzL2h/DyQNJTRHeI
dzl2ACZqlVP1BM3O0YIi1QUl6izz0f44DpxsivTT1DctnVeUjF7cBYJ8egiumZTy+FL/XjoH+FB1
lWbzZPb8t7HHQREvKntvE+nsYmjURVUYy9nwtEj9gvK+Mukmi6RruwaFzCQuVOuc70h6UCziEde0
/5HyAK3RYvSljZGmwZqWJaFyYSs/mwqQGcnRhkrSeJPvJntJntxqGeYeXaVmg63A0ZHMd3UgmMGz
A1lNVCBQm8O/N0Lqd64g1tI6miFY26nqIxCleJ3SEfwCHssjUv0cNYdyMjMNAFqtMO1aHAzgdqiM
+JOfoxjn62mSDBlNKlrPWbNIiUzZQI/ba1UZojJBTfsEa9rnml+0V+JCXvWd3Cg7A0CCoIyWBZoc
QGgzYxfmpdvuT7uHQed3r1IM8yx50tqQL5QVV2DYokSD2mx1BKALkicJq7SB+BchZQY6v8CyAwlw
Tb+WqSsJ/YxPfOkdghCvasRkQzaVYCwtJFxCkarFhVjNn8MuyPcm+0qNRsJeKnrQ7AmhL8f26m05
jlX2QnhyZAv8zZEPwV3hxwUIOevSTjIs7tm7TkKZ6wRK3e2QAB1kPKOoYxNkxfnpGY8jBiK3xx/3
nZwY01x3m1kZQOYVnsVPC0kmS6oAHNQAuvwsT8t/FF7sYoPvV723sr67AZToEtGE7k0VqEvCKQez
9UNKeyqH482FUQvF5rQgUni07lp2zHE95nsFj5utgT+Gll+JCgu9rOLVoKVm5b4OaqVQ/7jqRvkN
dY2rlSXbVP2YzMVFXWo3J/GdlPaJne4nuTZRWpsd/CFA9gFSXHnVW6+xPYLK170ir2qt06R2inbI
bF+5m0JdZsl41AQrh5Lw51BDu/a4+jgKEZHbFuSlI0CiYvLOQDW34c//KvCkQaYrQVT84lDcjmHt
EwMTTn7jtW8YEKIYuI5pk5UzRgpUPyHHBp6Y7u4vkSDV+rTUdNlIDfg3ZYWcdURnhHFzKgSwYL0M
SlvyIOlusimaqerfkoYZ13FL1p0dIWIRiUikAbc4nFQyMs+VMR2rHUqyuY63jZks1PlnLYd5REko
TLbke4atQMj/y1QnuybmkdoXICbK9arnrwBIhKZZeagZxUSU64Eaq1KbR9zHIqMO6SNS25Byyazl
AOcMQAsNudrIhupEnSAtf6EQeDD1qOBnjFUfcRVoFvkawVVAFB+9M3mmKVp1GLj0nP+/lUsvS7Lp
G289CKpMB176w5JSVbY9EDye5zGnIHtYo8aXx/fjV2kgtCKiMqYWd3zGIvLDiXefPWbVEJiH4TS5
STiitSAXvNFxsmOup+eGBqZTQWFr/gx3kLU4/rBYBqXS2prmpx0GnJvON8CwUhy4KLPikVLG6YPy
Nzz2aH8lELZ3pcL3ddLdQba1qy1HNl+MK8JiU3mvGIJBkIvbroOkPXktO5LDsiacNIlMaa8bPHyX
0XK62KnZGdKNR+Q2hd3oaYBhCtYIS5fz42cpSRqNMsRCVsmQstKYzROpshhgpuFNSB5N8UpZTPMM
rrsWrVYLYz9DpOgU7/8tYO9PnQujVdl3Jla2cBJWqtxwsN1lF7ISTiEKTOFaZk6BoJa2uMKNTHE8
BdCe/HR7rLoN6vxqqO3b/5yvSJk8ZlBrOx5PTLNj/R1CPyzqCa7iIUhijEgnvvbu3GA+gbLDntlO
2AeI12Wld1CHg7a5k7Zo6BJvvkX2v+expRceY98WraS3vmhQ0iZ+K6og01xHYjF69tZGijaasXfe
+q7L8wQFZzYtQUu+ZdiZQXMHbEp32yxro6cd1i0dQpHFMh8ZP5ociTmLjrcOsmZbCnNDhvTdzbBZ
D1D5JQX+DOsUfoJXL+gmYH8WgKvgWuNfE27+ADvnVpnnfW6/uEnPq4BesQAQjCy9FXzpDt51KsNF
pcOqQbOUyF5LVq/hKuaNU4v9SaBmspVVget1rrqLDAG5zRXlylKlj5h3pjDy//K/huSSc6WZamUw
Y1K7D2YtZCCCG60t/3dY08vhe8qOujN/SHkuttja8mRI/3Quq8WXqoxJveGGXWni2EESwdsRrvr6
XiJVMygtuGg6hhR0CwnE538l5DtaMKKppro8yXW8q+uBcnJZdVoHK9Nr1Oy7rPdzOoFrTW+SxaZ7
unMkGkRa/DQihhHfJIbvJPvQg9ir8OAe4cGnXaMz2nrkhoj3UbyTuGtXm8jEzNs47eMybugcprNm
JW4QsV53G7DY5BAu/w0MGYREwWH4Y+czlrT6w0+tTWlBmmYDe70dcmoH2n8AhCMI2v6kdtvzHYi9
pwF1LCi+aN1YDsvQTIzPaGRaw77BGRro0qOpAmdV/HX+8VL3NRtRvLPeiU/vX1AhXpI889ztiC0N
mQ+fzAlEPSPiIflDSJYZGGMtpOUDVAZ2DvCNVNUPZkKlp/NaaGluDX/lLsHTue4mgm6xP/YehHB4
wjNXSMKIGG0XFIf/s8TiCgCqeJWBrmWyzNu2j3pPWj+3xJDCmDbceXg/7cBXcOlseiEs+qCppIK5
XDKP4r8kJwrVeQlZoBeBxYiZj6gBMKp0u+jQ+nfu0uDUNAaezbKVPCZyLxHvOfYT0KFOZwXSnl7/
/vXObEbJnGLvpTR6YZmtOszkGrLWX+Lh2PI1OHoc7fOsyLrUJwgkg1ztH/cc9mWrLHQCwUvKfyLL
DAXWq66AQ1sEZN3zIH+J04NYJdAP0nJ2pJpZjLetfLLlbvUlt3sLIZVV3WG9CtYJ/nRfz4g3FNew
dSNhQT9hlGuem+Wl7FAkbh4+R6Z8NK9NdlPsytnBCVsy3oZWefFrOXCYYeKEcgz/zZEZIMv8DRJ9
0Duz5QOhjv0mKB1CT/pkKym9UiRG16KyTY1Bx96+/izFf+MNb+zE15adjwlDT6nehKoDjSLeyfur
BFbzEMpnjEXKhh5stjm9kGP4i1gk9WHeu2PCZgK1GPhgG69pYqeZKOOaQ6zTNncr/5M+rF12gcno
BouWOZ9Cr/gCock38KXNGFThNJbbZ9DSQMeecbZN8aa42iofKVwKQZ3eiU62hXLHwAp8H4u3cHfV
ScwZMop/zrnccvL5gaRAM4uI+SPf1H8K8Gkd+rfewZACS94Wfxohx0HDkpvfUoiWQzrO6wXkoN1D
F6oX31WUaC/WknznHmx/QPvjgJgii4iC6woTC9RtITEO37HQ/zfQIwkB0bo/DU/PXpewDBH3kLuj
dZhrz6yIKo1CL8nYcqmcR8uivI1axiuw3MVwWG4UmvWplLH4vudm8HQfl4lAQT16jNOUAOOtfy+w
a15jDCIhoAtFuT8b4elNfAf5wtSGrbCzHB1bsBj0rx9rzCi1SdVMhoALxKxPqluinqAIJK0iPumT
aU8zdGCEoW6uWnxpd1V0kXGTEQo0lnm/PwyvnhhGCd4ZEelVYO7z9EFILLSGwlddl0/Z+nluusrZ
oX01hKyNkLjZWiECLdSNZ7U7Zz0ZIUUbDsvQhrDA3DP4uQXk9yhIXNUN7Jk3YHv38RjstOxghtmQ
rrimDbO4kcx7cXcjZ57mzLQItpOrJL8YsTQ2qUXq1oUosr11FpGzcOvYQfCHQuyodVOA+EXE1mRR
GoDwOd4xEWWNagPh4fnE9s0tDXfAMZ88v0Jt3ZMB8SFFR3OaB6xetlmDpEm4FgfO3Aa3x6fOUBDC
rXqwyUGqrNsDzqhI0g/ZvheMC+yh1MtzfTLH0J2ocz8+q6b3QaGkmDixXSrGgR+NLNFkYlKg1JH1
9Yz2MI6EWB+gWnE/8mz/AZaIsaAPHgSwVRqWevakpeQ31QYeGoACgMhx/S8cbQ+C4vXXXAkQ0fWJ
lVWP8j3532JyyrC+4YkUO2ssELjUgAejL3rHR2DP6EaduwBQUdz1BGMqxE1D1BC94ZYwJTzKdymc
7jloXqzoXoud4EUtZR5CxUdVD+XZbYMk3xLUjICcZrV33ux7zZjFBqUQ5xzFklNKqeE/wgHLGvBz
PLGGbRs3HiwBAEbSzWUV60v7bypdTNYx3BXcGC6TnSYSTQ9kjKANEExuAuEyyUEerG6R0xazNsSn
/0bzcn3hEIMIW95RvpVYKvjuZcazvrP99SM3+XGtkbF4LAqA3b6h2jR/7RrStvhphFzMbtxRVCst
QUOJYFe5swugyKY65Hk+nFQBv+5ycQyoy0hFWxuY7ZCGELaEjmLUTm5R+Hy/E0GXm4Psgwta2Ew8
2AgkY3/M+ogAvY1+u9HWCh2I8eGqgFT3gRzjkvZcXrMIoDOhhsLFy3UmZau0Akptgn3iv9fqCZdq
92zV2DRQYCiXDxySiuFcciuHnUGm69RJX/jG52Hk/gdj6hEyYow6J33GgpqXBxiIQvSouhUsWQGB
36t7yURHgS3UOxql4QMKb6FNLIm62Lf/s1G4xid8V7/p8XcnDxoRbXEe0igTMoZgH/LTnvQzEroW
dweHG+Nwd62RvIpU3FUAdVDrabMlUp28xzFEasRCPfIJHzzjuh/E9LAmE394h5tZohg7eMUQlZrd
icY1uKeZskSNvWE9XRk8rTI6/ex+IRshAeOrG65qPmjTP0V283CAPw3+RcSAUMw31mzB/mxlKm9F
FbswDhxyrjY5qsWZa14BXpFKGneb8dwZ8uXkyoQ6F4q1cRHXbjobLcwuL1Gq2TpI9kUuphKRFk2n
wQnIzebXLR6Fwc0NMbkvA005s2kSSPuNOJwZpQhi76h1ZnfgjjWfTRUSXkUSKcDH/J3tbBmF3HYL
DGgJtV2RdyFCe1GAATi/wv4xVdtlrFshlWl0CoidT8C2NXR05SJUosAtK32uJiK4PusWqJCCWyTf
GuDDvUyRpi3GJ1R6XPHtcUHt03R/3yWLN2LPL8XLYfwqUVEwfhKHgeJb+pjQy3EdlvCQ/e0DFTPt
23feaYM32Lv4W/JRWLeI6mZFWhBV7gKqsxt9c75KqFeGad526utLYl0bWBB1ApFVrvttsfz7KgJI
TgJu8vHxHc3UWp8zk7pz1abveciIRjIHxSVy85sSSzIcfjWjal6eouDP1NO+Ffbn+f7OHxkyEurH
cZLhdrruU5tI70TK+566LkeCASVgVh9b8lkdmYQMk7kmsM9kdhoKfzI9p8BNm6ue3rtT+nzdOQbI
C9FNpsZAaqGB71u23VATcSYhBGu8+VwzOiIWPRnagsIzU2hib4ow7IDfmuhDBnQlEd2H/CvTH4Bs
8QN5wdDaToszS8mF0zXyZ+hicg9a0kRHczl7JkORntWVTjI6gdWRgCgUnmmnJm+6+PAAZ8gpsFHv
DYa8ufgEYi2bs9KCVLltosTeb0iXXPuAPpogLVDzv82wYX48OkaNHZgukcPYG5HF0od1jaCLO+88
ZCDd+aseToKEwC5cYGE43QBOlgi0NK1AEZy2NvcUoNudBC1X/3bOQgGUDk/dGkDKCxwNbF1qBoY0
s/HWRbPqiLDU/r4hXGAOxgzaem0gJtBpyR184IbvgcIecTSOQ76+DVl63DLVadhWpvQyQG+Zhk6v
3jLcWlZwziurK6YtlZiUlldioYTHrpG5egBSMgndiGVV+nuJhJhaoI/K8edAwveXtIshaAhFSSB/
9Ha9rqoM6KIUa4TGKEDwtdO0tOcV27/T/qQ1Eqt9BR2i7POfQaz3iT2VVwxAdSMCAV5ct6BJfCuC
k5n5UIOw8PhEcC01tPgM9wjkKsW1G1+j0Aca7Kgq3OWUKOv00IVRtYOKMRswjxvMXQOmQ6ILaatN
oTMYSoEeTyzB37fwa+uIoooDior3cFjfNT1NwhDuTrNpBYgoXL9afshRSbvXHRYlMJRdTOeyBN2P
gCnMvdwwheiidwUeuK3ekplDkeJYza4WtAW9VLHW/dRRk1rlKGMogsoJWMbl2Nzu/9WmPZNGHhma
LbjfzDl4EMi1/vRwNNuykStzTzZRGElpFp7Vy8WvRxdx6DJqPVo+PKwhQ9sB8tsnoI6Z4/iapC92
LPqGG8Cwf6s2jC/9E0DVZWuWT10yTNnNeMPSdj1A27R/I1u8StH07niwcFRU4ZTcQ+8nEXiBJ0mS
wFNRZk2fuNdZN1CJV4RvBMmUiekGK9JX/lQ4v6eIAitXF3plv3hHJLkjT9TkF4/Hgld7lZAzeR7U
y/SuQe5MZAt1sRubbmYPL8dcibba+WEVxg7Nee2AvkgPOy7o4/0vKgzWnZXvWXoEboJQaxAmAUo1
Bk/BuH+JlvjgWZa1PC5E3IiZTva1r9MydUu+CU/uCvz8nA7mNa+P/zQQSatAsBTSHgBaUMf9UnfN
2tRRHWM+EHwXPI8zo4JsFCCeCKvp5JQvC1SGiPqOZxFXi3okS5YcJGD/4RV2I9TDiBfMeYQRxA/X
PF7kkdUSe+hlBofOWIRLYO2MkowJg97HE339naq1yr4jqO0yf6gGYG24sqO+eLdAdKBLMifmOX3e
RGBNZmcbXgdAauvPZVNlW+vw9BAA86UCsaLdoLOaQKhIOBfUhULIiLLWE5KXYJvd9c+DahDB6dcF
Nzp7cVdRrq6rYypDJK9KmJbfVv4AHWDbw7JocoWHAgtv1dLqxnU2juv7RZbEQGDX3IE4d8LCP9j9
q7pN1FpNQSVwZ1uKQKDTnvr6nAjxgG/qCh7iSd78TVdpbDY2GOpmYjQw6VunTZZPWbMTuWFTp3Ev
S2iOxRfkmdTGiUfrYjRY5zjIyCwnZ0vJmyDBrFPJMPCj0ZPDFj1p01NyY+6YaJdhNA4wGqvo4f7g
jxCuwsos+MUtdjHaEaIw7cQ8lyKsI6WUgHT0Uo5TSxPcnwlNpmJ2ZrBFgIYHBHmhuR8uMCl4cQ6v
PWttwlKg+LljiAGhmLZgfQ2qehUDFk+xUKQg7vNik7tobuU0y+Og1gUqPu1cWMCjfqmhhHGQ22Rn
BRvpMlcy0v7wpj8YEAoZ/j+3ZAMYa2hXiY+AP1q8WVRB1KnCUynCAG57Cg4YZacUcV1ufrekwJxH
qhDbBZrls/EN7w1qUuRk7Lo7y4zy2rvh0bS9k4MqgzdbUg9KQ7i5K7JIZ/L6yWRNPDxaawQv3eBd
nxlZxl/k+R1027QklGLtQ0GPLYKBYMwev5oCLAEbsJO1LDZXyEHHTEFtr02EMMnlEKzYwhQUUBzX
GiS4HnMSGBkKrPbgs9UM1WKUluw7bzLjUZBFuxRq8EZCAowejw2/oN3gdQicbnwg7jErDWRgXcYg
b47RsR1oQ6QjJOpF4s7S49SzPgVP7W3HfS9xkOXQXnKJa6eTXGkdhD4VWI9m4xXs4hSI6/DkwVB8
7G6XXhdYjGmAe2VczfUHl5v3I1/8qLqk9OZrKiVqwbdpn3EHsHK7nS8MAKz3EndtSgMgKWBmyOZM
Oc0/VNnbcEzrE+CKmNOblyGB3TKh1+Xq4XD5rO7gSm0BvWRs17S2dHF4HO99Tot8cHIgM2TgL/6O
YYGih9PaYog5A7zRu46MAyz9dTRADfXe0tQ9z8YWqecrTDafzMW8B7cPwo3pkKhrju5cjpAzsq/S
AntEWoSw6xJbw4jgQGDjAY7FTWv2YA9SQ77EXw6WSBcUr4/6hBfDOiuH0yG963ihHkcf6bd5xYOP
UbxeFMFMHdw6lU+c4qQA3BPEcIs/e8R2DH4aDeWou902Do+tswtQT6paa21PqqkvbS3t8cMtJAc5
wWsl30z7SVtBgqA3Ypv2Lyp7QMcgTJaZ5F3DviZBLOergAjId9c7/x4IaBv9lFLt8gc08+VJTVmH
+81W1IW0CKiJHNIyt0uKpJBxUKL+U39HiSZuldvDYvGn8ZoRpVxJkdas9M5SbjoGO9vH++AkRAFV
ZhAykpRUZRl4ZFlyBwsES2k+AsllnQooe+6aBCzo0bfMCj8DoLH8O0Aw/2CS8UPR0/djnaAh72Iw
kGQo16FO2pdFYRLPnzag6wUWhfcuHZlGNHKzkXYBSy7pyyfQQStgXbSkxYaX3nK1KojSupiLcHxg
9dSlvkoYaSuee2IllpJZHXGBpB4eKx2sdscspFeg24WZDu+Rv9TKKqYsau3wGpR8/TP51h04pYHg
Rp5yLrliwyl1qnth4tH0pXXOwb5kF5UqQ6H06EwykuWCtCQy7z/GvAp6RZIKaokk7K4GoCReeHIW
Uo5Sytsc7ry2+agcoEeFiHXIQ3wi4Qmw2zbv1GlCOuzdURL+plXV6udNIJ4cHKR0dsJU+Mz+l0bd
NPAA4++pOEeouih5N6+J38mhwfNNTm4LXV31TiqNmplQ2mw/WCQ3yUNC9GZGN+ps9UHEfPrXiR9V
+UvRGRaMDhiKnAYFkBy+sM4CzzHuvD1SENGqHowvtoBQFd2f4eVNQd+opSqgT7L5PVV2lvhP7s7h
iQi+hkw1TuVOqrIrQuawXcFW/IHAIlRuAX0T5k2SmV4E9t7+LHrfU2Kxu3DKJbOqeUTBoXhaUC4/
mZWzEJd+xdO0glZASXZpC/BCGOPp+newNO2iH+mrKSTeM/qHr8OKh0o6QwZg0caxSP9YJfvdTgJ1
t5nvWyrKByCWtAcZ4vvBMzKPIwivQ0rtUvTRfCzO4y0zXJEXDUY2fChPdUL8pAYztTq3YWFYxsVs
KBimn5JN0GTUS+rYKD5SOWyuyRad4N7OB8NWt8+Hy5xDcjDxqBCVZPewLpqCBJPH1XQr8kvYCdaW
K5Jhzjj/wFkor77RhI564HZTOoXNKeOctam7cy/Ty8BeBNIbIrrb5FtcxAE1JTAQ9UsWPClMczPd
WNMvsoi/1Ee4G459BAGbHBQdY4yrETK+OJhJ+JQSfWsKtfR2bG2jyT1Nn1hR/3W3hfB+4qHWhufU
lUarWUmb+hvVSSpjaQb2EBXIqXYJfXSfcoF4QFcWBCuHJCf9B6JPVl2md4Xu/fZp11UsJAX9A8W+
hY5kBnLOJJhTGY8Dt9lt/zETGjwbj9MON/7W8a4cxLzt8UsEfIvUKKMPEPPFV2UVpH+g2XUhA9wT
85nZxYXd1EHpNvUMKaJVMENkgqxN2yTSNwPPB5BeWwo1Z02XCJ05JUPNZBAE++xFxwWqoSiYFpuJ
ph63zCCNqCIrmb0L8Rcd3sszaKOVbT+xdhZ7g2oXwlHQxzw+Nx3JEKoAHP+Ax2U7kc4T/AvrGAOd
Ew2ZlwMqgWGVgHOgc9D7QupBQ1V8x14l649K2q8My3KcCah4meaUtqARFmA1SFL2USJkczdIOOpy
iyQtXvXXAO9mLz9O8LgMZceoZMsZ5+Cl/SSrCQEykyaKlpKbAPWIYzzD3lfWZ5HDbbbMUbDGxNyZ
nzdZZWu0qtxfvtHO+naO4sS1htWSIEVs7gMxv1mOXPXoAIHTgaC6g/H+VecPEyY3uiA8M7Ezxklp
Q1pBOAl9SGTAFc4KKez6osRa2wU0NG8Tf97VgmsF6hZfGvZ1naCIGXYgStheFy40OO99Yy7UhGSr
n2uJz+lH2eS/CArxhv/C/A+khsvNKjw/WVPgc3MdQRiinHfz2nxcMsRaC0uYQmYQ1Nu+7CzSaYxC
rtoQXBb8ZpGgI/YIGfXy1BA5VBakOl5bOdSHbIB8B/kwhAvqaxhFkucNJYrzZeY7wLKXkS5u5u+Z
wp+1bpwRdVRnmpJZI1t8a8R7xtIuoECE5FWEA31uiGPDR36ZJG0Ltr5IlzhHhfaXArDkxGeH5p9X
HfjCO4Lbb8pFTy3LtqEQ+fOK6oO2KytgnadMXg8YWjdjlqprvk0OCWM4lNOr/lmSw6uVfmb4HuQb
fl8l22gT2sEtKIpVeUSI+ytjdToprnkF4QO9Km9cWnxFP2eDwhoIczj0WawxGBvrDr7jI6DKHS9w
eeGG2E2b4TwnIE89KU3CJDH90HwVwC6awrV1qrWPUclHUjrPndeSIiVv1GthkwFbg0VSlUVuFcAg
a+3hjecVG0hb53tAv+9MQYLLIcLVkOemK6sHdtCO7FN0HMVgycisllQipe01AnmCKSsRyaOUWmvq
kkKy/u8/5UYxqYZ0PLwg0c56hLnedG0JB1gHgpVxKVG3/iSDwUhNyhWrBRAr87hIkEsrdXRbmYUK
JyoEUwXCFb8jCFZBQmUwm5VOSYL7w19BwobZF7J4yxXVeFEvpoMyDJmVtLv53X1S4HP2Tf+hv7D3
AYAnS819mnAd4t6fgv3pkscsQ8XemkFU+bSaW9oRa/n6y7WFwGYC/vSISsgf5tNIb6UScASNUtiZ
mSXSBDe7yp00bq91Pv2V3ZOaZ1B+PpkHO3SpufgULAZPxUmTTmI6iWDjby6wj5cyk7lSZctw71tN
O0nhFtgm14RT/HGoTy6tMQEQWBhQbCxTruMtj5FsPmeJi6uFnq+9ubUeyoxzZnH2eRC6p0maoEmv
WByCwWvpgUq7IBWypSRLUSyXPHiA2scL01cqByW2oLX9T3aMJosM8g1YMzbD4mUMGMTo3Sq93jUl
eG6vLtIETVXrkC5FJaNpL2QcV76ZHdXb05sZRs5N2rOfcwy3QDDkZ0JzDQHRPL95nSTQ5DjhyOZM
0hrhcSuZpWNDOaE9GVHMsIEeLgZq0+BvpF6ign08PxG955yxk/WV86RxaCpDtCmm77J4iufAl3/l
g73za41bhRCu33PnB05vJ8Q2+VFFHQ59xGy5EFf/rkRfokxK+xCl98b4Ys18epC/dleG8wUTsPma
BUuFHoadmtTPhAM5rgwbFJFWA7EAjIiX/yNXj4ffFykcsrQVHi3lNBP4rUnwtmHRVoV9Jdtdeqmh
mI0yvvelsfN7NOfO8bkswEqYBmEXvD8oZbPGe84/nbMu1tj95NkoOkMyCWdwTiw7xNrhmxNOWqYl
m35+zPAMeo1OpeXZHXmo6dPyJvU9RqVrqVt1464MOq7XlSLmowgJwzedASBLtDRlL7Ohi0WEiqEN
q4XYSgq0YD7626mdZfm1oXWCx0DQqJvlH+hh22TucRtmp/Ib5NFW8uV6t01ziCcayqN2vmGVXbAY
kIHCJA+GsCLJIHZhdxUpEpLd1jKyLk6e5ISsN1CBxihYv+n+Xu/76SlmZ3jFfZTDo2jKYIMQftq4
32SWAycRIMUDmIKxa6eTXJ+gH8DEaGh2x+94q7gIfojF7Vct5okqTPMMk+6sqJiY2L3dHsav7nS8
q4dDeAy29iRqYeU4L0+PY8ojoLAHUqNAzyZpWy7AUx57hcRinSTDMRQ5ysNfH+M0zTT3wD80Qvwo
WBhx6KeP7rxnOsf4AUatlnD9qNZJe+tpWCB5u4VgVvXOn5+VefIDHGQi4w52KpoKNzoUadoQuRdM
RwLOq+UzweNHg/7IdHS8s/OPqGAEA1QRxr7v8F/R6qvjRK6UhSQo0BvpV7TgH/JL3HZGmS5m5Mog
skxXaA3ckqkfXa67iMd0HEJYbf0iqrCdNrcL1KPOl//Jlx/RFfzQOFbCuJjH7B2dk8Qium2e5+hv
oDSBMaQZnkJp2VITSAGKXR2ZPm+KocD5ED4DtErH257MGdP469KNH9yvhg/j532OMprcBY61Lsi8
1MY3ALYx8P8718rW4WGrSvjmrdwZ4ACQYuiiRo0mXEL8yBdO+dy8XPl3DORxqz8oII0tw2WmrTB8
/KZMwrzhei737oV8TgdnVGCWJPqei1bOnV7LHLRZk1G7wOE9NJSM+xJoegobi1jR7QwSN7BBF3by
Rt0xBgAHOA20WbB5VH2tQJNZsljDTF9+KaZojR6fyB0STLj7yD8qYhHVhf7h8m27PDyHAQDORC9I
6GNEenQ22hMlWRQ4QTe/iU03RHa2lhIlNfTbgDuXxdt0FX84oBlXnZj9Uf+B/6gVKNzlB7IL1CDg
js+t6TY2q4QCVfZvzpY4E55R6FLIf5viU7INpZsml9egeLeYf+YOFzJIyYO1V5E4ozHjTNGamLWI
buglu4dS2rVKwsRZ45CBaJnlFvHCDghO9qxKiQHxhXFGU/2FLIom/chMAacjpqoAM5ie4glzJkHy
/Yh+c2d4SDzFMgEE3WgZ1MgkSRxHi/0wpnXydiqdkF9n29wV5hW6gKFGNw4YtSg0FK5A0/qWOzLM
dr2RKc25mihyzVBAryeZlD0Xf30Ww1MEGsp9dIs0MhVssF1VrLgfK/6PMizShF9a6KIbENLG4y/j
hxfeI29ukOyFfId/6DZAz8VXC2+lAdTW/DY42q7lktNG1+62DrfraR+65lFdElVL6n58JJWVyBJw
RrREBuiTrP5AwIQ5vH8uJm93nvcOB2FqjHUEz9OonTXxNBnpmZQd7IXAprX4UOItCViN58bgMWld
8maU1bLRJUHMXuEjcJIkJZGTUaSmWHohGo2N+HptK6XlThRP1fD1PplKQZKZIGn8PuDYccmgcmod
lyNFgel/MD5fFeGuEgQdaPTTXMxYyJE48l9tp5DdwHnDOD34cVHLXsDGYoubzCKIE6Xd7HRmT0Xh
oHqaRhgGemiB3PxsCbI2rb8564qNu4U48kmHdIbG3dZOqUhSSlNJZ51MBi0TdOZ9NXVWopnahY4v
Gq33UFBqoJazjPtLLxg0iL88tddlcK1ns6fYig66qkBpv1XdvT4ViIxTl4vfC2aGmZo28eOzNjLK
sd9XhQKI+/04V1LMo+DSG0rVBo0DMTf0OSAshnTtXULI5F13KdfBFAhupNmsKSnQSHwg0c/0AwXG
o+t5+QVEB3BiQdljb94DfKqYPSozU1Lp/5PhmsIvzhLQ+OEsmDzftpilL7Q4fWY/ShSKcKLTpZ6p
v5o04NEN5ShRFHtJS+duiQ1Mej2hLgNz2xiXRQT/yCxJkPeRzNHzBIvfbxs4BSZv4sgbqJypJbIw
V6i5wIw+fWfJQIL4PDJDptl2nLgef7KHf2PTtETET9AVbeNkAcM7tGIymlzx1O1G2Mmv5QzC3W4/
ERHOdJlYfsSmsVrTNTD93SVwFOWpzBfjYpR8S3Rqx0XNehvcj2R8v1a1MdSkkbjcGTMOOnmHp2AG
d4wJmnOSAnx8yCK8FTh00a6iacf8O+f5DlSqYtDyGGWV2GXM7DHvc8COxwNjb+PN4GNeakkt9yp0
Ls27XC6wFSk55NC7raPj9IBAw7RGv6lPbBynvudhl2ltMt10OdECN5dyVi0SgtrN/Fn8TQxRRg7f
Wi8V5tUbAjLDJXME4PEZmWbXG/C+6V0HhKA/QCSIc2KJi6gKM3LWUJ8EibZhQMe/CSVXSs4pZAeR
1UlR99JaumZIspR5E+LLA75k8RP8HG21wT8kQ6bASlg1UqEVQuhdcwopKZKs3DXjaodo3ipbg3ly
JNvFJix7CEvlQs0gjHBaQ+M7KXU5im32RSYp6otmynQ+t4K55x4mtXbSwQka+Z9BYlIdFcPt2CzC
Q2zp7tFEi/TLabPetQ3KYS08lb6Buij7qAM3nJxSGj+mfhWvqOG6zGOb1+ARTKKpYfKTLq4pRZ7a
DCLpwSj4zGbsBJKEd9xvwUD58s8l3HsVQELLjw8VhWrYg6qWdRnqN85tKip5lqJa7EvuVgcXgbSz
pFj7T/1alrkyAiqTrypvmyXBT/wo9JhaKxP70TISXizMdmcrgsooCSrZ5OT0HcWBsvFxBi+Jv7uO
WNxA8ey7lhWTf1oSi+0mDTvNoiR4EDv6Ru5qWtOLxF0Nx1UBO00nw0kE8FnXSoemza1TwVjdaUMh
1nARyu9Bhn1xm4oUOi/w1BjcZDRsAhrPjXRMRSTFDKoRGJgtjaP11XErP+iScksiJ9ZcCCreIWiA
yVx8VDol0FtNztbGX76UgUrA2Aq9X119KICKr/mlzajypC1ql9hgyGk/QRYf3UMWwYaYn0kIDs4N
yG+pkkRIbFAc1+uGrAmSjiQYA/Pq1Nee0dNw1ivVLGHdfYvfY7wkYfoJ6CIMgnElNCyYkeh6lap4
NdhwvSS/4mMNI48Y8oX5kH3sI7bUQC1pxRyFKwn+GJiDfTH/rCetP5QfL8a9Z+EdDREcGlUo8IPf
kXJg5F7ezYPdapx89rqUS/1vpoiMio8+watkAg8RJmXUJTBq7NuDPNWi65FrwOFM87QD7789EE5X
7Qe5PINSmIbryudihBMPcoB6Iwjnkdfcy1anqG38MLhxLJ+uTkeEbmMyYnJ8cNPLoaqKM5aGTLFT
SO7pOjoKra1W150vhwfXU/raYHShQqNe5YmIgypRcTR0turT3cUCZwdrjwukIAoTdyqlFHl/mXzh
CYjxhxu21inAP6NCZq9i5g6FJt8fK1fxNC1qB5A7vPuBK8cm167V+fYXO2TIWKOLP74XKNsXwyTb
RbIL1c6JO2d6YVr8GSyENNDv5OfEO+ZokfDiXmEa9q0fsMayzKvJ8HU703hb4LjUe7ueLRM8GF8f
hdnsZVo5SBp/ZIm0tagBcZGvJ10gswyxvqy3lLNE+HGXdkCqLs7xnKPTfA9K/wMJbZjz+9RNdjCu
bC1t3jP7O+SFptd1zXzONRBRdnF9ZXQ3Z5yupd8c7Qj81nApNSgYmKnvwjouttGBataMZRMG9Pgz
G80D50DuduwgwaxyUlMS5ZYDahC13kYd4g3snMxyRjZWEbGN6Dj8fDgSj2eKmAtjj3S7gMWBIVuh
+T8GOKyMTNNBjBLQ8A/IBqJvBPC20vqysfG3ZyfxeG+r1VWo8/i3vSrr/JJBw/zpPXqm+bNloaE+
mqF1cjJs9OP5/dgVJMEsmq3k4dMiynq3sKPJ3Gt5LR03Yi3Iolob61N7gAeaiddYJx9bM+LpLNDN
/nv5FvdKj9uA7E2pvNj6vBm69n4YJ7rpozYaOU9E5LGqJZwT6j3kbRRY0ZU4aSR79D3K/sWBkLoU
iu81XBRaKvN5JflGC9EFTwPGXM32CRtLwmHo5LlsUNw18YQS8AjXjOhQ1fbUX74E3+eb7nnW+odd
kgWfnClRlYfisVmH5QX2ps3xdrbul/avIrQXzZ4kzzq8cHNQi19lbjjKKR25/JPSF8pBPOW2Qd4r
3ImdFHhwpJSFnoSrnjOiCPM6FDX+5RAVYetO3U6j2Chs9nJKWINS6tGU/Y5GTfPwaOrZJr3gQ8uZ
11Yy3VzwU/jKmiiEI91fL4c3q6l2tPAqvJwHtuHgSWyAlYsBaU5hnJ2F4JjmdHgUFfeHUpjXo5i2
/ZqDXinVoyYdO1BlCOyZ/01XpXSTZCfWjV725aDiqkqu4xJXjUCsPffUc9GzH31mZBpjiaEHArDR
aTlcaqNvjIL1YdZ3ojHDFWoShc5EqDAcCCGTgZ8NCNObYZfF/fjn9JdEWA8o3dREZ2+VUAyXf5ce
qh5oRPY4cwpr+av3yoxZBNzwBTPnMsdsbrIWvTENdhTgfqUvKec218mCPpXEK9J9brnVnLv/obg0
rvdugn5WZ6HQSvSbritu8P2bEe9iK7gFMK/NQCIBNF9bHBv0ZtWCjQV/MSjgVPvJ7n8Edd+q3wGv
Ud0DBMDPxOenwJ9W7xniS2RKZWmk8zshCCMtDmpKDmeb3tay+T2XjfaPPKmbm+lwna1HEkPNWQsJ
zfNy+O+861ZErGKyQdNkg2sDhgoBkE1wS3QpPFLijkWUQAfwmEJZyMV0v6k87SzuwvXLZfInVNYd
l2dg6stH2DuRVGk8OTf+amrtW/CgDhgW6ZQidXF0c5Ed2YHFeGhEFhAutLGt3Up6afTiOOO1AwzZ
4jQP2/xKaCUcRDQP3/nYx3Ijg32BFymHFqnViof2u+Xoapq9WQaIQVXqW002CcqxIGA2JLKrdnUj
gze2CakU3UQVDwHWDF2TUskIkCy/PVpAKPbTh3B/WKKmXRlvijHdgnBVrmLQoD8ROKyVJmyUXKK6
Dl8XO3j5ro39QMmkab6CoY1jJAv1dJ9SkQ//MvC/JVipN/Sc0Tk/E4eWuaDPQxO2rdu16EQrM9Yb
03ovGPzyPXXL6PrtERuz8lzRwUVtW6MJxNKDmK6hRB8o3qVvB7EB5IBthGBdfar7RH+YyWDC5+R+
AjwoC6JnJoAANBIx2diZz7OiI79Bp2tqTYp+n6X6gG/GsOGUPWK2yStzJy0pKfJZ7M2HVzh07HCA
R0usGt19qhBXdfC/FDmdWdXxU4ykGBt2aI+6AxX3uatVSg0Zf2opEJhaPG63oBw4wBjRwbblhZXS
htUz0HdKbCEsnVddRMmTos9M1op2B/J9vabtOYEEpZNSqVymAYWN0HX/y5dJ1NEXFC5ov5bDVF6p
qxEU23CZ5oyuTQ6WmLWel2RCH1/ErHvK3qb2VDL2RKyMA4ZZKKNgLAygEhpWh+Q+/EjTgRiUH7un
VZ0cktIGjVMamie4nEpXxmljlK3U6rfTf4ubkB2mwNnCOIASVHpetFKBQNDowJaWMAdtERu05sCM
KqEsDn3750+4UEyn8hRdGirTEMEIosnEPWiBwze+8JY7a4ccsEUzrFT0mUtu86Uii9SQblgF5ycW
ixzW++ogAekO/nwgmlw8JhAHhHySGQqZyLKZUH5D7J6k+iCnNohdoNj9+k8WFDmfUDGz+Tr/Qcc8
7yUBkHTRyxbUwrnAgnI/dXN/VWLy2b1od5Tk30JEl+/KV4K12D22g+TAObwZtBWdMTqdxXPHoRqd
xeEWFULCjC98FMsn3eaKESycv2WkRbzLXaCRYhsuSQWxe3MI7zLxn4WD3Og213bwzoe7blIkg+HC
NxEO2vM+xvP1YzPNpbDqSuXleEMdcy5WMLaJdj2bfO9tDwwu32b/KwwX6Eo6pZMcC0ITCsVN8m8J
KqaFVtWW/PgXKLv8+qIEQl+zMm7ZF74yqdGnG/TWEo7yPHjzDUfxbHrZHuRm2E2ITQgpR0pTkBWs
0bueSOpDoE8OdHF/Ot/yHw5aDpZw/EiNQPkRvzu650asKb2rg/sJSjsdY6hnIXVpnb+RtZS8C3My
9dD5pVnMgjXh6yz1oyu4DMYVd+YuURubZ3ft18Ixym+QSIulqM1hIjTItqt6qTHeBoFMEOCf/G2A
sJ8eZ0zwgk0UOS3Vmh2HLI722HnqgYbVLeNapO6FLQZ/4seeE7GwPsDp3g8b0yLwa29hY47KOfne
rFQE+7XN8ZEoDaIBigL4G5fwQaHQroANKudFAk9SsaObuAe+/joY9mwn5EA3/uRaF6qoaY/r/tA5
O9SvYCWcbHBkqaoenLK3DZ2qwj3VhnNt/DG3U8KAe8TN3k8UAXMuUL/Y0ujCu9ArI9QLKGjLmDH4
csXivMzJ+lCXehc9KiSu1N4YDF9WqjczZ6Z4ZFytAX/eQ8BAu+ePIXUP6HDhfbdDA/6Tw0gAvL4W
uzP7O9b99H62l4xbUK9SKfllLlUoHO4Q3PaAvLFo+fElNAsu/JDCCvJ3X4DGlDHrles490EdVVNn
lys6hUCIsx/0HlVxeGTcMq/YZvKxhOnD9PnwJATJNH9TdM8FwPMuNvmy60zX/tFMXTOfrtmsjKb9
HOHMhUjFDRcLlV5RkPivJSowpxZMhQKXeTO9u8b08pVR/0/+Caxvzh6ySMH9NuYW+VzKq39OYzq2
yXTJgZtkTMlLmHZ7yuNtX3KaO26Wjkos/zTzjf49NxFImlOlnu14cUEjQ2a7inOxCXuHTpIJU+hD
9wLk0DbNR9JuyOMGYVFjV5jbP2bk5MjkcqdNxWeZKDyJf3Kvugte6GUF2CHvL1u2jFRauYK2gBCY
z6623pekFVaIMRzftVMkwt18eE+x5eyRUIvU9vBP7Eocw3i1iTDasyEZBkYlmANHWtqm+ViowL4u
/5CPtttn6W0PnLa7BxqP2zg9LP4dGIlLdftqkyOHE1EL21bGafvEFvK+7qrNaXLzwl3Ddm9iFO7H
b47vQqEpqOlxWQtxauIzvcR4Z1Rf/MvYsY4Wrdxv73qcZL5XsS+lA2P8FI0my5VU70YhNEfk8MQd
6YwGNR2ZUSXf2XnYIKNW2zS093PUBSHSYyKJaWQIUHidCJ+uhIebzLVxTe9FX0BXDerUFVMBaC8Q
cZkd/LJ42X28iYyTdFYzJqW6CMtMXMh1JlQuLhCg8Zmd83aW9YeoQ0vBSm0GW3c87592cq5hkdKl
DFBU+KdHKylOVy3IZTSN5jZUX4969Tbdupc3G9zciEwYbAKETXoVFTTTudLw8gIwSFYedfzHUbKE
0fNDQEDkj4SnCAfck4O+x8iH38BiWEBPYS7n7YhYVpmgoRW6xfIosQbIu48w4wTpcmkH1CE21P3z
H6U8VSPPgyOvNxPtlVtE6S7UZSuHV9IaM2+WF4+AM58OA81Y2DmOBwHmN6ZY5GvWCC8YKMGj2j5b
/Xzum2Tf7DGf7EVbyjbQM33byABrPHNFeU6rIvA5ZtLhhcRbYiCzOR6uevuSjkMmtK+Utty8Tdr9
HNLss5XAXTrCwOAIJYIdpzn7pcw9ZJBWIrZQbXMX94dh/HmLuV2vZIT9X03qUxnMF9LtSHZdzFDV
A9laxWKv2tKYleXfA8zzxG3IPPDtnVE6kjPgR4PkZoYbbu0ro6stU/oSXC9FZ4zPi6qSwckjjqa7
2ErvWJnr11O+48gtEltm2HxCLzktwFz7yQ8DvXbFCa+LIWSjmsIk6HFUEUicLfXmzqXvn2BRQSug
F33Gde5C0RYloLPfEtfGGvusYPNpgG0KI8oaSIwTrDNJ5VaX5p08w+U9ajRaTgbIuJE6oH/sPCgv
flBGcvOoU5if6Q0uR1jyoh4YSyk82qB+IP7cQ9QmjbacvPRSYDrcROkN0q56sz6s3XXfLHbSjHRx
d7ZvIXQG3o4BTGiEKehYq+BfSjjk0Q3MMv8GEKRsDUCbgtrJJRa8xwM6QCTI3lFPjvf/FIHUzVDh
1B/7LQZHTYr/FFg+Jp70Ff0Y9CWES0mhfYATVm3cOytAKY9zNZbfJkHg2ZlAnyPyNm6yG21EAsS3
jjuMaocdwdCJUSXmxCsN4ns6Du3W1Ky5lfIA6kCk33esN2gT37z/ixR9PMNL9cyw/GujnvGd1Z8t
l/ZYZmNmhW5ZLcRzIz13L+DU2wmTKx3K2My5TxexL4zNWzmdVynrLF5VASvM1eIyL1IImKxzPC3R
jAdZJuIE5y7PY43YCfPVBR6UqbHmakUaDzPyNEuZy+rt4mi+BMxqN/mxrM6XGvdKl6UabtfZwSIL
sxest7PbQ3Lzbbniqh1kIeFD4Czs8Amag1rFWq5MhEOriUBragRLJheS15bZ71I3SxAnvmNPBiC5
68N991vWhoEE6IGirdWLbgMeugmqaQy1aRqFYwcF4BUrJ/FzDJY2k8+BxSbUvox/6XB3V/YDiGLI
5l2CqFdypeXg6dEa8GPmKZQ1nQWy0e3s44L/MN+4BE6YSXDrw9B0pzbi2ak5BX7rR9RRWflN36MT
5Sm2EQcJACL5+4p+vt35dlNOIynCW1n6jvoWme8NwUtc8EG0h36TMjc8j0msk6gZBYyMkm+XRFgO
OgPNHljgupHyCd58PsLp4iHXgxdsbwcxUB/JVoM3YImoGNZsBLp9JRe3fQl1gSG9QCTFAG3vSczh
zor7vmRsnt4mLd7Hl7npBncy3AsO2Q2LC3nGS7wlr/+klVQD/HojR+eC730MMt8wDMKprXMllGto
lHzJuK/Vb72Ghs/FVk855eaH9zI4Q9bkXSvN6MOSj7s3Xx/penqJpM2IubztWKEzo5p4+2RR4r6q
qPmQk79ODvDk3MpGktoCLtlBau94/+LHxYg/5YfxVL3xHac8+IGQNDAJdpQzlwAwR8FrWhJqDlbB
6Zm0FD4NzxNc71/OYSaUaqk+yui6+iI13UjGpYcAKMwdjX54/n/WQ0IzxsVPbEbQMBUXuiKM+RRT
yzUuw2Hul6dEtsXx4t1+4Yor7SssTfThmv4G6026PmZu88OhrGS0gElTiap7JJ25ODAWFegq5vA4
4mA81blv2v48dR3UsM27L5Rpd9fLIVpAFHxQHt8Um3KaYmoMARF0sKkaePQYBuDZv1IGQ6cYeDl9
XCNq0yBYP1NspxDlQuBwaNRA3+PpOPmHooLb4uKtdW0NgyTWC+ZE+CHH2NGBUthotRSXO6rwC9NU
hWitBrCeNT1Pd96iOlZYOPjf4OBYEUO+b92ECb8E0iS8ux8+NaJTLA+PeU98m6ESzmIVt8wcxCwA
yV3iochsiyVHSTzY1l8Aw938pV9vMbiLdmCzV15Rda6vBe06mXLUQyw91rCdSjTEKYq0fXJpPpf3
HGGv5NdUat8yvn4mi4t39nZSWsI4KAW2OVrfcaE/6jpjlVrSMElAQAtC7HnS5cwZXbNok2NUcb4k
4DFwwOzl6ZPRjdehfKEq1VxDYeyumGUmfMjeBOL7pfdt5VlzgOjrmfKQj0oc5xigS+NJXLxxz7l7
DB9YfCC8jf3rqiJoOyiX3EZ6vF2gnw0QsDbYMkPVaAezFw6wdGHcgo321hcEUUzOJ3Oj8rBdZ4k9
d1CmtaZxBnYYi7BLHCtDqd6iVOqP6oU5ZKy02Paz8OlONmLz58sEGYb/xr1P04AH37SeOl3SyDD2
65RQbV7oKMJ5SuIw5r+gVjJJKcwRoHRGyH3aCoXtPPayi2VBZMz93vzi/ZPIhPrjLMedwvUaxmF/
RKQimrK7yxg6mn4QDj5LS+EFwGDg4Xb/SuP17GRQpBmP7ttSZQCg0+nk/WLNBE+/5Y3eYK9wuJPb
QkfgyjeFfLRtN0jR5NlApH1wxTJXeov45CzZZdA2V+sxAKSApT+HUlCjrsLsOZWWpl9HPlYDt3dd
soGLOPuMff1aTQw1vYNzEAPi+8MVYXcORE85B4T4uN3NVNMcJ1IQgEN/Z5j7VzdUsnK3Fssjd4sh
oFGWN3Y34psstdSglx7oEjvWrtQUO1utJA5rt04pQ/0O724eLeyYrxNLjJW/ssxDJDWhsuDkwoDV
9S8E1reEjHAJNQCOy1P2Dulh1HvEX1whO6kb1OdDYthS7XgOai6jXcXC69Mi6I6ox4fLNsx876dY
y45PlBeEcXvZdXhtcckxCqnDyafA3kQzgsBDMbmkkjy2s2dGIWO23W1MXgMvR8H9RoV7WR4msisI
tbCgw9kJKFX57zSryqP02pBNfXmKCkq6vaRxHZuPRowe/xpRw99Ivxy1bwVWw6RdQ7Dyc50xyvS/
bKjCkQgjcIwuSdC+DwR2X8USTRJ1zcBcq6TyYGHsYGoLjb+ga1rmU2WtU06fz2mtg3xiZ95bhhS0
gWNDKFRDXw0WDCnA56BYL96U2OwfL4UwWUbk1rdh39Io4RJSleUTE8egIsqjxvhGBS3Du3wOQYTC
Z2H/vkX547FcwnBsTLtU5/T6F7wuQpYq4StJFtlIsoCn24cu+7W1wqxUUiUbO+P2qocK89a6zH6P
+PfEZsalP8TwxGD0jwNyU9coK2Aw+ShIV058iFdwQVRjlVS87VIL6SrP9BxuB7mZq5KVm5Tkv9SM
j2UjeSYvquQ/yYH9zPHYxVMUTGZsJXs/hsKCOgS7FD86qKdT0vo0Bjz1Yr9VVZApg+Y95PxDWF+q
0HzJKzx7DpC0Rao+VhIYi6VGnU3QpANBkOiw+84ted79XMcL2q67xRBHt+Cmmn/dlKjfmW+GqwMp
bGPN9M1qGR20VxKwQRxPl7vxaZp/RKG2pnFtZXieQK/9QqJOl3hm5wP+E5Xq3CzO+LHc8xnB3Js9
2OAK1h2p4047diwAyX6/ilcyz9F/SFP8IAEcZhwE4ARqU/GSdY5UEuzDCkv2AOw86XuTdSMtSaNM
bx7bJtMPrkOPODYZPWLiGdBNWG+8xjIh9vO5rfzLtjFR2zB1ctRVzn9EWo2nhOuwqd5hdaUoSLvi
4e9fZlB1WPdhZApMlN2AztyvEt5KDIfSaY7DYufALp8ygnKjIc1hAb3mcaNTE+LdL6x/dGHeF9j2
zL3aVbUQjufiHxuDq99J/1qxmXVL1ucPKWDXW6UY/PZiVXmTrNxlwCWcSHJTcw/qQzlDAPe5ZD1Z
CRAsD+De90WrSYrnV5rXCUASC2WXSKtaj4GXzDIvX4icLo36jPorXSVGVRVv9qOYYO/VGJV8w0tM
3h89Z3sNf8zs35ML9TBN0tMmyPsLzBepJU6oDUKLA+QKuc/FVaeWnxE+5l7cKKhYEXYG2MM0qXIW
cc0oRNyDsed+td768FiRVkrNT/yAhWnDDGMZ1i6/H4jLrJdoQhEoLzaYG4xQ9shDZSaFCAzHpF05
xoZglMkvYsLF/dfCocQuk+PEKQxQhTJ8W6RYg3Kn7ikX3y6RTiHP6ZCflCGmTEkv9sVY9WqWhQ8W
u25wLMZqpmtvWHXk4S6wvyzwoLhne0ZJ8Gm6DRi+aSbsqT+sfsFgyaRNvT+r/yTFo3gsG8MTdaCd
sE2keBISEava2c8sgkqN+6nm7+99rU7CZwKPa2RJ5McnIuRPHAC7TUcf0S8F6M1CWjwPG6yoso/f
7BgW3mKi+tgKlAYOqZgNmzjJ8QSokjywRtTsyzaDLfw5OkliQGzB3l+KpVUmd96167WngZT5yCwX
UpJ7j0I0n/Qtcr6oDmfy6o4ZRIRWeuQFp5Hml89PgnU7qe9Onk4EwdlOdZ7EndOY/QClrMiIWDlW
hDL30nfT4jkce3GIWydA1GM5B8COCdJz8yCXd8IuOWLwB0Mr53urEYrayiSt+SizT/4unbyE6cKN
eqmZh3NxY6iSQjHusOrluANCov8AxF/AGMrXA//jx1kBgJWAB8EQEKMUD7xNNgGI3BxIpnKLvwKD
5o5iJVXzz3sdsq/OGS3c6jXx8VMI0Cizm5xzFu+MhWkt/ARZM9NgpcYyi8csrJPgaCfTHSqfaCwQ
rQl2qSB4xTTuI1U4TWB4afvmCMPO7Rt/T143V5YYA7NlRpJriEeOI0LW8ehx/pbtRLxTIjtZJmst
xwS1DfixOW2BK1Oz2kOu0sDVTm9BZXAShWmrPIXXvGi4Kz4xZAsce3azEX6cOY7C1hdnHjUZ8GBH
mXCSsmIpMAa6GejwazeBScFfX40i8alb/1lNt+gHCjJblFhEK5wSx8eLz7TkwDatRzIfKwWgj45m
3++9iTmjODE/cmUzNziqaNQh5jRLg1NeT8GbMqJC8ST7AQ0ushLVCLTlO79yPD37Z/9opWua43wM
uevKtT0PU2GfdrkPsDw0DN20n7Ysbb1Qlq+tYSvodBDin1zp9wr9Ri88CaF2vnkZZ95vfr+m4dAw
0pWtZup90aTZgchg/Iw/+NrH1FAvhWV8W2bD9S8Oy2aOVR8StFgnSshwa/3XDVTcnV3qw2vqpFmw
UP6bwBIRUBREowGtIdpO4Nq8qReU81iQ+2UoQ+yz+nwVyZcompgTOZFiKWgSkDzcRqib0YqVADJv
pmHD4VlL/SVxTh3QXhiNUNAR9IZrj6yjPgUknyjHDdnHj1shAgXpUrmQA6BYRzlGAUjL15DaAJXp
wxFFR3m0BWmIC/Afj6z4dNODteATGDzKpceUEZKNDHVsL45PE2OrfL55PnVpHO79inCX1dq7xRbO
ogrJkMiBarPeihgJoicygtkqTaO27B6D/LVjvsyXWA/IrPnSy0IbVBz/7nEmKCYI5B2nVLPCdhFX
I4bH1oZZ4INLFIx/tGqikZsGBcbOmlTXq+boKRyukFsHLM2a0Lf2K6znnXGpuHUu/3VK3ehwNTw5
TSO/bNh4QioNviHXp+l5VjgyfhK41bOhZb30ZfBZGjafrVrvxOOKXllF2jb2APRglZmWwOIWIZdi
qQmbtmIKOOFvRzIt2NhrZE09oHe4Ry00P3ewLA16F70hA2B/GSid9aLL51HUUQyF0M1I4A0UASIw
apckckL61T5hIAw4xZe0pWvxalCQg+ZOWkOvxv/FJSl+M/UnwsEH23AxvlV1GTLW+cVaa9auB4Yd
ad3XKZ9m/XE90ZhlQ99n6K0WZDtUcU/fUZp1HEPc+aft5JxNnSWyA0DGi4b9xdhf54aIn8fZjsQJ
wCo+G8ZId6xjUVPx3fRb1Ic2kv41xEFcO2Oc/piQaYXBRQVJCh1D7nS+GkWHd60kDLwInieBjYpW
vhjM55J3gOx2eneDXs8g1hiWVdNEiQNX4/sfZwn8gawVbTnUeJ2Cg5x/kgWBwf8sjdx1xrNlGLy+
/5fjMcKI2HQmBqYp49yLKVMqz09KZJYampY6GNCuRn9QKs5YrW+MnB6eYJYpvw38iUOkv6Kiv/U5
WJ4Y+2hPlK2ZircUWSqJI6hJm8GuFOiwZfRtO6PhAH8t2k7yqh6Huwtb24zJ5dNfUMtNimQ5tw6Y
yHew/kU65LAeizDhxnT/xsyH0LlnCo9+BD8/srB+YgHQGFXuStdfsBLGd3r6IAKrYMnCARBG8bJR
LCpUek1ZyWHXqM1qo35Dpxg2FUehouUKZ4P3C0GT5HfB4KaiG5dxPQjxYaAxFFdYDlDr+D/BVM+a
TcYifWFIgYHf6E9D7KvJ81K+LMGtuYDK31zLEZvzeBxSoDD6C41E9hv98LUzronBLON3xALwVLpA
TN3qQEUXB8jbcbFlMphQSHNc6FlHXHv1NhNePdgJWC0rc4sEBuHS7IbCEG/EdCmOtuxQhJ18NW8Z
pNEOBmh3wI0sTaixqACWi8LmrafbJdnsVJz1l0s5m3LNQ1cLQReMtIjY70GEDXbkMghN3Fmf4B2Q
CvJ6sFW9v0fc4pw1DKkraSF1zOJSolJe3UDQlXAISfSEnrlftiKxV1n850SoOJyZ2gsQlzOO60OW
sWLZZgmlwbuULhJqLP3Rtd+6j+/cOCb0COGiCS14ddBNRGC9QynETlXm7OiJ7mqDiCEM/YmUBHwb
ptdEHY6B+Qr0rBqyXDLnrDx48avz4cRg9UBALYytzGJw8wuJz3d8tCpn/VOOvNydv15yk4MU7Q3+
saCqQ+Fz9xgjYaIoNwsRAPjFZK/XCa6jHsW2McG2OcUS/O496tIDq0fCm836PatcQwvXHKqFzXAS
kPnAruFhtTMLw2xIAY7BvgWJf8I59qtL0RI2qZd9Bhoa6ZEtTrHjbhOLnkm6ijaTVmyJTZzNjvA5
loA2KPxJn7r5bbB+Q3U8WmS169ErgqqT+azKkxmJ0HHYGSreFp032M/7tq8BKmCvg/dMzvMM5nYS
4ZHKocXonwIxVoST/rZi4cn6Hj8najQHwcPX+YIsB4lGtgSc5p/y5Rg9Gx8q9AeHGoGZHnbcWI+X
oZfhQLWwwE2C7HzUZXI9K+frIkqAi/JljoTGwn7pNevy+fQgpQ9ZI8LnJp/j7dAeuERdH4Kpzpcv
oA9wAiivIHay8GcKQaDy5qCGjbQCXGSvwOobrnzywECxqAGuUwNEvoyl8Tf3H4iJwAPBiC2Kkwud
qARE1SspGlPEanvVqIL51wD9uNe1EeYoxXhPy+M1wgkF+nWIFy8jBHawGw12KTvcBng6lFvHhEhf
/HG6u2ixAZGuCljPawU9i8hyUvWcO7rkNNZCij0l4N1TWZIT5cHhIc2e631dE7ozjdU0JzpuBgSt
47eF/jEEa7Nc/WPbc1d+/qQwosuBOG19ki00MObQ+bUsvPfCgqC2CyXUlQlD36jkuhfihPFNYnD0
i3jgo1FJ/Mw83L51j/rD50X+P3Sx/PfvqJNaRQBoDc6YoRZ5M92Fc0InWgOXihLOhqPcrPV/zJ2W
UifdLlEITFrJynkd2adLkwy1Mb4yYgr0e4tBYu0EcVUhjaazI6OV+z4sRr5Zlns9Y/p8NIOjJODA
dQcCqaq7EfjcTs1j3/UU2qvYS74CokmGr2DgdqzskWMMS1cYmDjxSeqeEny+JOa2bXCqnDb5y97+
aXEjAWeYZHK6+HiDjN+tgPODO8FRETiOy+lU2zqQ+0EIjgZ89feo6He3KCa22RvVXxZWhf43QRty
9yTOOz6lCLK9hddFShcRvFQQk5Mlr+Acn/DU1AVcxjZuXIkEJOTB1FtxPdDLT6sq+tEeXYsqwx4Z
2UES2IRAzsCdnPhEDaNGZX4idgOmrxrqkAyKjcR2F/5BSOlDlJa8pRLYeW1qjS3wv0CnwUoXMFsC
zlSSl1HHCOaM7HFMdDMd+XcRpTlsqVsyZRRIbJpnroR9iix014VoQwFwcqzzZviWCiV+QjPqW/0J
mRX4DOdlQiBEy1Ifo/M5OQ2O/MVMFLmzuXYSvWf822EV3yEG6305Quyv2vc2NvCpnIrQuzlp6zgD
lz76RmGCLPtCKLW9hkHeTkr9qgc4NvxDXiHvUvVUeJ2pW8AOij1jFrmonOYHgyQdhozwWIiezAwn
SR911pzpftpV0Zp5GnB7/6GlitzpXZK7vMuox185L2JczRgescGW1u3Ykfc7/IJgOZhcN3INYPQr
sOdkVkScJJFVl5dxGN6hOqR0IxuckdE9a8Ic0JAF87sqStT8FzuRejh5vJNTkCu9YluPo0sYZU6j
xVti2B/NvT3GncV1w7605RI2NXrbZUiN/sO/cj6okcxrdj6BlIP6TRjAMv2eTAOM+e75JXhLbIm4
orIfBQ9U8YHDWhC7P4JLAlOdnX5Qu2SSOgYwYB62vcw3yek7TlVn6sEZ+fiE+/f/bilQFAnFmw6u
bX1p9cvxAHqsmK1fh7YISVMg5T83YdgBkLhHeDyeu+KHsur6qzK+cB1iMQbPVidN/y0N771qhF4V
1lbGJEnetd0WUE72VCx5pMOlEgKoI0gMQTHTJ5t/GDJgDMvOn6Yxs7RIZw63t2k+U4HPb8meKGs8
qT+UV0wJSN+Y+l53eIOw7UILvYBtStZJydcX173wvdyQXMQFoA4DJcSYLq32OhOM+YWoM96SR3/Z
x364RGUuMgKqAxZwkB56wjEIh1Kx4yqggTO3CAz09vfIEn2qtFvAkhiPIko9zEmgtNUDw3IBn+NC
R+HIPhrmrcUiOQEdQ7umpitzY4V37ZdNoDQq+S7k6JtctOu9rP2g+gEUDOznl6chGogo9lRZju9K
pIlrzGv8bGUQ5w2DGrFFogSmvS2jB2NWBnPDHq1DmToBjkNOzHVWWIvrsua+t6GaLtMfHmgnfFH2
EMlBd07YiftvO3iDs5RvwAocmqZRIfsGz/R2FD96Me4hRZ+JVI4MJ3JseJUyr/YwqnOOZReQgmg8
uBQVIMQ0T51i784R9SISTXitJYfaT56MXgaMKvshYE/MWqTeDtZ9+IuDQuPr7JVe05lSPX2H5XmU
Bc8m4C7xW22y+CuHRDV9y91h52nr5LzyCBnoJr2PK+sJECpTDPZtKQ914xj2pK+WF2oMmyPQiK47
Wyp36kzzWBkaC+Qzf+Jv3If+MsJs9N0xJyJfQv0TGXuL9TOFDeiG8pj/H1oPq2RQGBtJK2Ju/qYU
ITUrWTINPXQLwzSagA8xAYJyhjXSUuxVlZqSrV59wMACLJna3IcEn/256ITDJIhmfv8v+vZQ3ZvO
uqp7Gjh2crLBOCLb4bgmguqReO1cbHVKenoG3tQtxjWvbu9p9KUFOL55IowLxeu1QEX6kl1KkxV+
m43yUyWLzSwO2Z1RPVvm9dzNmI6CUckcFJ93eGpXLBQuSJiL2SIT8Q2tSz7DtJcihnDbnJz+HLkH
24REzGPT0fV5Rj65Bkk/Z2gy9mpwZ/pj7dFR5tY6j+U1vgxuprrXG+wc2LXD2ZimNAoIhKjB5mGE
JtweqWbo7AMYATl6lmCw8KdmzMJUFNE3msE4/IdgbO7sQde000E0/auZM3vF+LeI9eZmvnO8PTym
dwjXbGhMsA/gClAjyIA4QF2msZZQFmOab0sK7ECZPac9LyZOuIM5ObCDg4R50KqlGxW0S/TV5u56
YWCzmIegmCay53vSyQbhx1cxz/HASDV2z0mVKNcgas5JaqItZskKvYjGb5JRiXwHzp0tlPVbfHlu
kV8Ks+Lz4db//DQoZnvZUJ0JN4aH6iIck2ydjozoL79vPQWVazwDDXfK/sEQOyA52K2DLZJpLPtT
epVOtPmxAU0XRipEJHT0PgIlR+EGWpXNAmAFiTgo9c6HTNyzEoh0/sZQycwHAd9yeMews6++8rwq
QZdXA0E5p813b3iRwz5R1+8x/0QUitQTLN+/nlIsQ8U0hSkA146ST2FxiCkr1tvlRheXf7zUF6ke
5NwuRYgI+4NPJW0mLPIO6beEYIWGIkLaqjrStkQIvsuxsVxdGotSE6Sns1B8hjILUSSK9dKM/2N7
IS/uoEDGlayjZsDC6sOx2griPQXu0ps0+RXG+PpyF5kxodW6epGkrQDmPS0NmWkNqIdyuTcyTxCy
itUl2ADXUyjb7NFzvSc7SnzMiDDVeLM0WgWxsHev92JYQq++g4C6KRscJxvEqZ2iOAczIZ/wDZ9n
8rZka8SROWpYvhuqCXb/uEoQAwF7fEe9i5XkW4DPhoEjrP92IyCgkBXlD/iX8yxQIrOA5xNiI2M8
rKdZdR6sPIVqCB3Z5tdfEgtjjSSBgYgLpC6MCU7zYsNsTTazXjuOBPDyUgpdp4D7Q5uWfYewdOie
yXhMYxbKiMdqwELMChlC3NsJUrxLR8uwAcaldBlAx8EjlQXZ4cYPPZKH2k9f6HXLJlTNuO4yPUSl
PR5AuxDxaEN6cZ5ILvvuf1fvBzazIMst/bpv++2pjDGtDm5J8SvdIMs++8hPueo7PUlaTNoFHlp8
nnytWZenLTkM4urG/Td9rPhTco9+gqtom9RUecG3FVHV7pE7GuLJ7iD9pK2u/c0/VSuToN/DWWsu
W6/ZeKcyJ/IkqlRFQEepN79OK0yS/BjKZNVxO46TX6g0/FujIQfjcDvCmCDuvdUhFgrrEvPLCK9c
r5WgqjFwBMkEgn1HtI3ZlR0NKIg7jlqseACOPReIY6yu8VttSdrd8GobOynjz0i1RSjjntx/Z+yL
O5WJ2nHxoaHjawgN9g8aWgfUMoRA20730JnuFYZ3TmKV6Jrya5t3WFIoZLE9V5a828Wkl7VBtML4
uVR5CQh2SftoFSNm6s5hLYlh7jMjH5GyI/rGt8sR6ya0pKQVQtpGQ/BVhG9n+TCuRJ8Dm8R48GKm
8kvFn+BkLb373EXMWz1hnSLAhUfcNhx56dpUc0UylzfGZ0nUxFMDJ2A/HE+YYowMp0HJIStIxEwz
CWeBNXWvADMo/Xp8/2l9zjW3NdR68uGn9meALoLKnSP8cIpH136kmLZgPDk/8wEWPPrEwNxYBFmc
dxAvaOwQjztDDhHff/f+4+K/GxvV2LfyRCo8QRSXZU5WeFzHbk3y+DhA9iDrBIndnjJWrds6L0Hf
p2k0fY1ieyRJl/qJQRoAeI+CSZyXoC3giseKvOLPlPTLTBl8vQrq1qXsonPVIe4Q1T7C3e4IlC9E
c8I+R3U5FS9ZGVDEpVPKg74WwbVMN8F+hT/Wor+3pnTIcmgurbq+kaTZWp9wA8FmF41XRs3wFcH9
GgtJaqm1zftBRf6RSl09irVyS1EyDJSpV/eK1HzbIE1Nd2ExZITm5JhoD6rhNOWo8XmA90Rrk5MK
09uwEKkYvzebL9HRMd+e6qVsGFwfWf5rBlUOX5Li7P6q0kHO2LtndnoFzMEDvTKQwpneVR7d8vjx
g185NkSmTpRs+w1VOiXgFUg2W+zp3yZCuYoEjIKnax9psGgnfchp0J8RawJvIkr1CPGZNlkPcRHs
qYavOqiFNg9Gs0+Fu5/Z5xbyy8sbuywOHpRPlZmesjhIj4IWfIiUzZo88f4kJFJBV+iro2MKOnE/
te0VX32bnLvQ8102XJe3I1b8c10Jmc0IP9ctfQxsHY/+F0dD5Pr16BRabJmpqh4NYY8bfOVPzH9Q
JwLYHBAZF9k0PSLyhmHdhp3dedqKVSVpBcm7bg7OdV0l6aAkSQs5YWGnffyEu7QxJ5u5FqpDiagm
es/1EJ0urX89oLlDO0raQ9nPjcWS3cEJmtXbD/6/FxGcea7WxjhIL1LVFMCULSeoxNakeu4+sHES
gu2RhkzmLIGFcKHuB+zFIOqm0ZtV8B+ijRjGUtxCFY+vagm8F5msk6GGxdJti+FKzfdqSjR2FzHD
oXckjIJGtj+GQ4W1g6JC3e3+KWJ9BIADPTDm3Oe7sZGs3qdUjFr1X1bz6Uq00o5zz59edV/O5UGJ
qeK+N3gtT7xeYVNHcgNgOFq+tqsoguz931MnNMt+yeBOys8IAPTt8RtGDgwKvR6Y5ZfxIG9m5OUu
QtqELSCAnjgMfDchSa5kRsYVc8DWC523ZNNEznUBADxLAiHZ5DmkDg6tNCeflYE1OR+Y7mNEXnvz
GkWcHcuL/ll6+qFp+YKjfF7yrsphjD+OrB4kZTJZfHsTCeOhZp9jeazEppr2GxveTUD7lCdji14F
VvEWM+oJV+Zy8tmR5FacgK7Gwyr1v8CEC0E0c+0bvnE65B3yOA1YyUVof8zkkHM1WESqDRuN+9A0
3v63E47Vxw4LN8odGGjp4X1aNqAH94YFBSrs5TCeM57GHs3bokSzyZyv6kkbLHN5zOg+onrtYag9
Rj13J8u/qy20XZvB69509o9dc/Pu3M8PfYs9A+spyy6NgHrkk4bz+49AvCgU53ya4Wes2jYUkQAT
nhsdP+zjg/dKc+8y3oGdvJEe1oHkOVLaSl18R+7NE5fK7yPy7Sfdp6hp4NlYIAnvHHT5EiHmX+Yk
UzZewv+XZQYcyRiEzs7ONrujuYesoi65Z+/tlZhS2q7c7wbX+rdWFwMSZdyBIQ7p9CkTzOHCYKCU
/C55fY5F6p4sZDDFMFAvG+GCxK/Esj8g4vGUoGsajKlaIOJMFVJd4TCmbw7/c+44KJ1kf1cMiLo4
shyM4WFwcr70O8jIvcvwHbes06faBdUe8WV7927h6lFBrOYTkCvXlqR/KeW8E+WUkO/ruWgSZprN
3n1E5RAZ5FdsetNNnUpTRCfFDP8Vq0JMN17QJaU46culOF3818xHzPo7vj98RQUAY9E8tC+dxqDx
O+FFz/+9NjN49riYHkKPl4K2aWTSag8y+4PecAxJCqXaHxE79aGA6W505qXWuqQi0A0sgHOHxWzv
0CouPxWeGL4uluwLjhf3P7psHA9AJ+wL59ZjQx9LEp7YUNnNffbIc0O6hpsWy810j5t2SLcxxSp5
ORmgvILvkiAyYoQ3uSzXLFdZ2/+Lb7JhxUGefSXL6ptI3j2M56Vp6gZgi9PPs/JOKD2lJ/JkuPQH
SslBqjEKQ2ykQkElJDwzWqvOO5Pj6+eEBPRt6XWw9j/kbPr7w97LUM5S+/7sYE+azCa+hAzbFZ67
XgZXBCDP+uScMGwAEDjhXI3eiOhqLcc/lda060ZwRnF+U8I3kVJNupGuZv/endZQYRiBv8nPHzP/
3TQSxxzdBlS9dLq1R3OuquryzaN+gNkfuihviDHR2IPpc3FgCoJKYOO7ctg4hN7pRozr5AiXJ9+u
eX9IQ0fD0k61l/vqW8/DEWg8dHiLhS2hebJ4fYUx00A9l4FdxFtXnNGi8yKJF7FFRpinREb0ByuG
Y9ObZexUVmOoVRwOEoFFd2/MYprhiXvvvXJcajd6wWiH1q2qXJbHVETw+Bpkf0IHDP85SbqfjTsw
YZfBCUIR1QEttrcnLEKQltDKUYmQZE54Ltp+XEYVQ7JXFyyB3+CTgmvFqwES+rCvH/N+zmvB5ldN
1QH/CGZlNSewfNbA9M/Iprziw5t79+n7N5/7n0xd4yg5wh9hnSgQGVBzZpHs2yUVGF+1NMSeIiAW
2HiVZ145IKFT14yH49fT2aN3Tbv51WT1/LgMFRr0Os19KJV8nhd/iWNqx1v1ik3EvvgEqg5+NV9h
oOlv3WPqNfN5SQD9eQR4+EaeNOxjkqNPKSgZjUG6n0d12878pFoAs+ojX8zcLroQTc4aLejV8zyb
QWa/NmXLAx53j26LaV5BwWc5CJeVB8eFrT5v1YVIwy8t8Ao+ppSXCnmTjWGJDC1nvYyB83AD/NQq
eiCwRtfzJJ/35hmeIYMM7enYIO8AfFVINOhvsffzyEl3z1T5sXoT/9qf0I+B16c4eEa9SbYOdq7L
/mq6wSYshWoR+JJ6srEalh6FhkMvf4bdMgSMoIniYbRW8r8Qr34jfVwoZ3wVAPNiy7JVzt1N/BBb
jlhArs+4N8qzKuQe7D48dUfYvrqG3RJtNNX+ygX1i3f7Z2nGoLR5pJ++HE4d08MyhLXQ6gac0dIk
fxUMhCRCo9X0JE8QjeF3zpgpipjc3llL0uNdEvwcobbwPJQ1qmUPkqY4AsyJlgGiA/RRhrm8WuFh
vlOIgL81mxtt4map2a7Sul3wtF9wPSaUvH6VrkjxqBjT7zhMdC9sUv+0dyoypRqQA2t8KrLGDxsp
8Jld8twropQYiQOnfCA2uedrDXS3zVIjg2SODlaCXdONe/zo/N4QahfhFhtHOzsV6v8aO30JXgna
d/yV+hJc+rAjnfXgk+DWm1Gte9MKPtN7jPX7+/c3fwn3Jn36fxr37pKAkYfJd16PC5Rnmct550os
tUSEs/pmkhxwJyHMqub76G3TrLyfibD8mYLgzND5/7k4df9O7K1kDg53NK15hd9ttkZZfw7o7LzD
3tXL/gfJpz6mr+nb+r7uC6KjU7TW7H0qzlj5c6Pab3WX74Xkbp1vrCRAqL+iNG/s0F2Lr9OhenKH
IVDnSYpmXs3ehF1xK9PvX9WMNFS60WcTnrpyEudUIeJI43+X4nYYWc6DnTMgBpAKeo++5KyFqzCT
TUijFZCZzEJoVhqExaahhNF4/y22W/Z4mf0it4IbqIeLM6jKnM4s9wI5jqou0J1hB25Mweul/6AT
QaZF2oHVsDhZRVfIxDfvU7yjfHVIf4WIvO3j/C++ap3h6JiwvBzARGoKsrUrCAP9FHCuaIVYiWMR
bS9c5asbuDY9uydmMUNqpImqHwRS+YXuSBgwr5tu1cecps+CdhxgEnysrbVumRafZVwmgbGZDZaD
3hq8ML5kz/eHJMqTP7/A1w5X4MYkpAmeJZhN94iBGNl/LyCJypp0y/m0UJUeixDYVPzx8nj+bmF4
aw2e8Sg/pxJsRZTXeB2vHaqL5BTLq0d6nUVfbRJ0+tp3xhhn/AAUzq0vUP59lgJaULzRMCCKWkFN
CwvBTBuUkBtYfjXRZlJyfgjCWHwEv91WbnJGBh+0EoMkw21sUCvWZmTnEMmOuTO6WezE/Wt8HMSu
AAXcPX/y1k68Wx+SpqUyqCrW9QEQWXdyTDv7qF0dsVcRrcuC/3cBmIW1Jt4UCyRk05/LJhlsCFPB
xjnzy6Zldb8qomAH3huAw6d7/X1V78tA1ffgtbF7EKcA/aBfTX0flGmmsL1RrQx6J2HztZ5KGhAw
ELRTbieoBIliyBN46D6nM0vg22pOWqUHc4814Osx6q06GkWjOVN3IVOjV1GsOZgusEtmRIYgz48l
zKepcuf4+F/t7vz/p6SN9vvZGbJyV+cilR4cvlB4NDdAwY5i8P3gw4nnIzTKoW7y3OQk0ycXuKRS
kZI46KDsxqFpRcKV/RpZn2AvnPRzDXkp7PkJ63+cMlVJMWXPRVTMFuuKTHAtLUWsphO+YuXMCbwc
1rgGjVWBET6LsU9uAI6VJy6U2zfKy2cnv5sWSJGcxcnSgApBP6WFD5C23X32Kysh6SYPLHGWbY/9
W9zWeO+JWoak5pZ+K4aX9MVQXbvAiCPvFjQ8Z2gsjm5fk1Dapm28EY0esC+JzF9RNTlaYf5vJugd
ryhIt7CGnrlGJ0zFuxa5BhbveCIPZWE+j1Kaa9OrEYSaqFoNKNfr26/X7koYlme9v69SbUDRPJ7J
JFqVjE5K4zs71hDsrhHqhZdfoH9MXc1am+HbdUT5whU5pcBAv4Ty1Inc1j9+B9/3HMlePwHIW5PZ
OJLgiKXsaAIrU4h6//pMuqnztTUGz2f15MZOPAOqq3cH0d9f2afgMABFmPGoCXD3E5xSaJ142lFc
F8wDEej2JpNhgtTRoCablKvDriqy19enu0mKpiN9Ho7RhtVegN438j/dGDgx0RU615jegINYJLou
15wf7Jl6GzeqsLs97NncoTgglJeXd3Bx3cRpgD38HwdU4qcWtD/p5BCdqW8nlJenFKPaO/mL01OC
YfCOwAzHBMAQZBJzOEbBtsrtETkBwdOlXybU7U0oHFgj0mWsfxCa1Tm0cCPXGiJ9p9xQHqiYlr5B
7/mZTospCGogrcvlO3rjWSvLWEpDE3jk0soerIqHYQ6hCST9rdMFKu0WqTFMW2k3QE6zpRF/X6NC
R6kOiUb9YhR33HN62Z7yUEDbbZXhtOZnxo0UCL+698FBjWjYN3kLfN5UFAoEoO1sLsa/aPeWlUX9
FOK8QfqJ9hwMhDDkwb2xU2TPJfhxcC6mDoo8EYGpiUnzwMSMf0WKppKCzU6ABtINNrv9VQMDKSdk
WecaNn8oTIvby1LMLmzux+rk7GAdpngg+ohbdA4M+TeFbRhE05amZjsLC4P5+w+qdl5x6HtaERw6
bRvKSyiFIx9pfhm7FvNXY8hSaDG+kn2AUkTJcgT/jjWVOlAQvNI7CqVUIGslxmyB8sYN/VudlNqW
cDhKaJ7TP+xksQmOKPzRtqcaPzkz+noyoZMVR61tmnuazWVpQ/zezCiMTeQEYFU88Lj53KU1UtY0
EOgbaRgW7IY4JlEEzF7F3y7vg5fdE/55k2mBhvyKtlb/3KSxYjiyE6D5ujdmnmbfelUbkVVlq0Tv
VDvqjEnpd0B7rPWNRjRzxkV0c42E9TIrGdEiHBapkCBpp6wrfbJkJSV2+z/+JJwkrxZeU7EMnwI+
haV4Z767cJFPLZKcjL/AxsUIicsMarVCiil0sOcyL9o3n2ma6n4o5hax5S2lVEyKJM4N1EA7g7cw
EL9/UHE9Sts3diZ4WFhN3rHfd/DVeBR7iK5b2+P4jo3cnEZ23kB50rOtYAzTb5mKfwvtcc8tDZdz
BiTr/T+5P1o9QZyxMRznwBiQUvUeoYo6UCr130rzYVg1MI95BRMqA0BjY/glIUPKG/Uefsfo3vBQ
069wRFaokGzthNaUEGnsjEz1M5blzpmywv6FaFSReI8EYpK3NPyCDhSLjM3Yp8bkJQJBo37Ou+dQ
nn0CqUdVi/xQFE0pVUid+MKf3xVJjFEqYyDBkpkzUsplaoss5hcvwnyz3HaucHFePJKnI+GRNjM9
719YpZdmNSlViWcMs3yuq9gZFBBIsyAayl8T3l6ifhGKagJjiRHICmMT9oV+iU0ALjPrsv+rDJAX
Hqm0iBQW1KShpNa138gAN8zL1TTUMTYejZ5YNxoDIWKUYLMyzn7CFONRO993GvWxk/4hFZB+WIwY
SL5IaN4VKXxd74BKoumfK97W5aKAkP0vfEMLFUtmDB4DaVzYRol8TVPPBi9QL74oMIKsGAVNQNF2
HYF2xJy71/+pP54sTBS+3Tw6FeJH5ao91cB4I+N0G7uyw1LCbDTMkSfSAI0jh/Ka1QKoT8OW1G90
OPLcMZbwa1uJdZBd+bYglf5M9GAt6Gg2PjtZUIHH5gnpmi9NHTILQxmffA/HQZOO1TfvJkVLRKzB
QvPaFzjqnqBgy6SRTPyZlH1ABuhanzbQTFpAQlTB1U7IUE33xQorTKp66xrTaYeiPtcuhNpeEt6m
5evPdVYdRufoGpwNhUn1zOuduupZjrQDtD5Emcp6O5LylP/xGyR0mJ+kOCKZRwWeC2/+WCgq9nd0
bmyPqB45ow/3qQY0lRU1f3cRC3oGB46TPgmk3KjJyrBllKLSF3aneK0g1ol+PUzcd6GF8r3prOPN
6L+JcS6TwWGVf3tvW4qjITwsTwETpImEEFzGbK830E9irisebqclq7Ca0CUS9qroy4acLWT0C7gr
0/J9nypPgNahPj0KZEPtvbiZAo4DmOsnC/KlE66+7DErMsxbACiYS4AhTZnRSlo/T4pYtjBW6Uyo
oA6cRu1VC4093pIMf9tMq9qMuKyZlyiCbN8vvfSx7UMezsQBODGiVgkk3skOZJXifmcttq/M5FlU
dMTlRTfJZJAUkV7hx5eAp+tPaONEhOgP7AWXCkgZnJIb9PasMeJEWnBUhmH06i412Az41ve0dIbA
RKzUBkVSIFv+AvAWxX47bmcUHKLBA5LLTR8zFU0ynFjfYv0rRktfMSpXM+mjJYNQki33vxZrBcaK
DCAusJqSFHBR346w/BcS7MTR8x+JI0UT9BcL3d51fRKM6PpKOug4qSiS4DQSpK/BY4d759emZCBP
TcoLqlZK0Sn/OxphHaFEz0LxQkzzttAaQp+HvLhGvUyEUHP5okEYw3dP0Mm29/OYl7H8/nXWJgKK
V6CbC+GGUMrSYl+jrLUiFqO6pMpNbtFisgg2LuBIbRzQCSAIoaqge12zJgZvVm31s/6BUgtl1Mjc
QUtgsmjgO9nIsbU06A76r7owGfpGzuXTLs8gOUZMZvULTbpGr9gxSdpb+wA4BezqEdOoyLwDJoxz
ZBdyCgUPYFMwWhuu5/Nr5Ct6M/cZqfeFPxeKZ0MxBkvOUOyZjkvpIzYjL1HO2Hjvgm3GMQ4E/8L7
Vm9C/0jHyzBRhQd2jro0Jj+9ylF7/nSAJXQu3PU3Yh60Ox0j6mhSSAb7HenPue+/GcH985iF3PBN
Pf3XvldsUsdz/t73HJOK2+jc+EOG+u6eMsLQX8Q7ECtwCu2Ogp5XWi9hdaliBDrqH3oczu9Ex/GE
ypV/7KmHn0PoymEWj3oA4hSAmFrgYNTHldbbbkP27GD3YczOIQB/rHE/vgGSKBRKXqGeXKAYAcrl
2dZygVd9AbD+eHQ71GMSLmKah28/8ryMYdOk1PkD2uzwT79xja6au46LnA1uYG3RD0HzJ6RO14Eq
MGuJXTMtP61LetEUD9vJJzaRrZjEHRWfVePmWSzClZlIORRobvXUwEsGYel3YqjqTjixDN9dcEMT
FF2hhhk4YdMJ+iXCnNFmpydNbswSGlivi57BhkQpZ7nP+HjZH+DFW0nOETfxpmLj5UNzzjmBar9/
cKOQP1mm+SJ+TkTmzT+K9YH7C2W1WzVUL2wboRDGD9jr999vWrDGthcHRr+SgeCWxHBho+S2daZl
cpK5lb10RwWJE8uoM1NyMt8Mg7CVzEyFRE3SFdY+PhckQ4zaNmUvbT5+F/+WNkGjX45+5NFWFFgA
v6DY5t1wRPecYVWov7kYTl+IZrJXlpzO11OrmECYeY0VWw2XfueN2nPXf17uLnuz7SQaAEZYMcm1
vA/zHSIx/yfqTzD3yF2wZgLS7R3Zy0Qi3dbc4QbTElbND8yesIeVxTDC7LEDenY32M+OIuDtq7MJ
kOgzeKMOwa9m5e3SHdl3TZQ8zNdwBvwnPe0ygf2geQdnLq6bKvm48jO6ugirWiSECLfvZtmwaUKo
ya6Mh07x/Nb4FkVQUkisS7IWct7K5wlCHMFVq+I5a3TkwPcZ0ai2chhB+eRIF2x6J4EFa40S91/9
pL395bTOt3D4FHiYiMWc1QjJ5F2HTg98bWrIwChoQztHYepFxbpqPIQ56R1gUThfp6IWc1mO1MX+
ZSCYvbx7C8g0PIuYk3OUQXExIfQTOUg7yQfchGyDZADTLSif9SH6T+Lh57zM8C+y7DeF5jCz4dWH
/29Oy5kyntrIkBsh3f3BBmJPoNgN1FVFCNv7V5wDS25deDQCkcHA9yPTScdGRJULCGscwBRBCRz2
0k98Zv6RqNUp4+ulP57N/9cV6C2f2Dh3YfMNZV1jh7KaIDHu1K9QjFbPu87XA55V8g13dihOkuX1
Ui3zQ47pEN52fqZsXVV6e7IEVZ5VdJ5zA16cXZp6cdGIyJkQhpzk2Zp0n0FdA2Pa6lf+DBB1lkkc
FDu6sHGiNjDutj8oMsEBEBJ2FmF5/NZfeHQf+qhNjOeYwSzEhbexZE5aPbr4S+4GizoVvw7Ypnhn
jkuTjeUCid01H9YFs5ec9fDNsr9e30Lwti3JV5Ys5zk653gKW+pF49K35zVX+XAiKwXXEK2/D3Ck
SGHJFQ82gwBOJzQIB2jn4FNU8KqvsjvbpvUBKHzaQbdxp9pVV+4Rl2AX8ryJb9JNPsLXQ40J/OPQ
o6wakkv8M0qZ05I2kek70G9C6CNizGvErupFDbQ3Zq8x+Bv9/zpsqAWQbY05yokji7ejt48UUD+y
U0UuMhsZfLmvaTtHQmEcZnGeeSel2SaMd6En4NXT2ePjyzonLuCOJgpsqyQGE1IPGeV7pq/aC81c
jw/lClwSzXcSOqNCnOEEVN4uLEsX/jFHJ5AK3WIZpk5PnXHnwlMJ10depXkKCXHtcmgQiFI0Cogf
yuoT1CSpgnueBpvgWMCmNQ4q0k/xbobRDI0iiMp0P93NyED3W5cE8s5PURYLSsow7LWyRx5S2zRf
u3qMqSbCuTDSuV4TyMtHpGUnLZo+CVO558llVGBUDgBmcYhvzCDj6kJfAItDcQXJuwIks8g8PWcv
oNjNMXeYtg0xt33RvsPlOC7lz7QIC1wQyVuHyy5FnrJ2V9jhr7oOcnobykNMLJHrXn40GqSo4lu0
/ruFbwave+9TM5ukWO5I167ZzKF8Q9YsO+YVvnjE+sjLlVr+htEI/S2wW40arroFtSYKBDIhs+Cs
/QWaO5Nmv5CXK1kE/tCnfcvdvOZaiZp9x7zC0xANrg8WkKbOzyvuOy3iavXWx3Un9Qd0EnGlNCcD
M0IDfWvmVabJgC18KsIBi87gnSJe8Czaer6hQbvFn3ByDPW7nESSSQwJ1cTfq7y2TctZq0a6cfWT
CFv2n8s1ojkNWgoR1413kLJWoAEkdbvZsB2tRUZ7H53kX6pkzH3Zwz8e+q/YbBjz2r71pJyztxT7
Jf/aQ2MhQ/U3x21pRQH29iNmIVyEotHQZQYbCv1fD75d6vt73PzX8jRXLos7wPcDHZZL8aILuo9S
hkzBcUbnqok6EELeJsj3bFSq1d34TXlSJq8uftYbtT5MYXFp8kEdy++j37F3ugiN0+evgqf0g+SI
CSv+BkgXE2Gl0TgI4MJf2E4bH6f728KKuBIPLtovG34oPYcL2uylt67dGveaeGjDuWNmvKSIRaLM
dln/xuwnKANJAT1Y6AJVqNY+xrprIXxE+Rk+zEiaTLdFHazhP/PMQJhGsnWSYMV0oDXS0/A4Srnj
mmvPqg1UG2q0xd7ooY+039CJpLQhnlybTOfCvhgHfJt5l53j28BG0PhkPIUZVgBxfsutCo7lW6qs
M7TTsqd1vEaZEeaaLNVtjlgvSuH0O2y2fTjkkEMbIuTcD2pRRgOwx1JxmbPIozYFwgBnXXq3ljIu
2qi+OZzM3N6O9wLPTn347nKoGQDRvXo7iMx8XB8dbMKrXt/95Dc0pUzyyuAN48vAR7H1sGHthT+U
W4pi1abTTL/RQtu00z4eYATa509iJyYWtQvTeayeoUIU3Al3QVX4md1YvVtSoZDpVHdmd5dqszbp
vGeeqL3ixnO1FOZU/53/vNMppDT4DlSOSh9vvCZiD9dV2XXDXoP6W7b7IV0wmT/Rz+OkW7qHmTcU
PFOpHybhBiJjwjbXUcxEJ+UT4HguH3neX4eg1kC9vJ1EHv+HW5QPH0ZBMoKQzWn58YlozVYD9tZN
Y+PSZ1Soj8wI3fq4PX7S0uPJPo8fvfxmc5FhHXB8+NBtibzmQJDXKy1On3hasPjkJdfDqdR3SfqV
znuIMBXMyAkgjLgXCZ/Rc/Sk92eALcVJtNR0C7p+sQ/RjwKc4geU9iK11w/DUuFJifI+nkjpBwZw
kHrN7W9oXwUwj+XYUELFGJC+6YIfWC6r4tbGex5B4ZSRmtgTAOjCtlMt3hy1icAY9G2VAFSZWLcQ
jJ75lxePpKik7IzqhZxjSay9TidtOovquQTp83IYzrD4Hjs3TmLYdcC+3I2YFJ6SAdxXIh9vRNB6
L9bHLcUyqGLIw5yV+AGfTTMihsDgNZn1iXJjI5e8ZfnbYCFEI4FeH948/Pj+Ut0rDjwY3aT9Gn9v
ONGU004uQotzur8Hppsf4UxhsDPq/ugAZ56LKLTY5DLGM1YGYxgu7WcKRjYhtfRSc2c6T9oQg6rH
JaX/F9P66Sfem+zXJ50mhc+Wq4OPUUOUF6B8b3yrovyQfSGbdR6U/bO1BcLbxi1N1ej2SkOQD3a8
fa849mzen6AFISBsrTekDq3yXCJvxruy5d7JZ0G9L5NiFCSP6xhXgkb3ZPpus42ycD4t8IKcAbj1
LqRRa5vLZf9b/PzdK4HNalbfProX77dv81cHkCD50BAAxigv3P4h6lWp6F7Ge0JQC3xG0UhevMpO
ksOS2FRMUMd9bkkq/eJjGRloCPlYd/px71Ej8UEJMhY0EGvJ9KH/Kfnt51kwoagdo0KmjjI802i6
FvJZlNtVEd7CY8Ju7fy6N15XbKJOTBdSwN2yLf7fXRnoYyju/XDYnoSr6zJ3wKEJsucsx3hI02nJ
KeC9cnNO84EXSQE7HQBHGW4dxRCFobYl4xt0dtM6wWJIle996Y5z5PTTtdMEFGmSMXrbfGHvcNvH
GsIkMiHFES5K94DUM0G7+4TGqjXnZtcGCfySwdHf1O3bhNez6t98EtekRj9tsd86VR7JlXI4r5Cl
VRk5/bom0D3Tvw8zWky22ut90FwH8OTca2CcoTTkbEyJQ0erJtKnEOpR2BiAGFgXQxLju/OEnM+Q
hdYj/mbPrFrQ/LlL+yHcyurwEAKSDGMVbfbto0I2fxNHPyxvIHNK42X5kFF1ckHddhJe5ZVz3r0I
HEjlwWR/DckRcHEbNfbkkg81tULPLe9iEDql7tcJ/xTFJ0q+Y/xXX8wnhVVxwCxj35mnq9F6WfqE
fo7//boLfbXHrB22zLIQTdjU65GBmwLW9/0cL3u6E5zdJbT5+RLTnhcNoP50qwj2wX4x1drBbLvW
zoLpfeNIGJYsXmbyU39SQ9ZlHZsWj00oapQvKZxNRiCzIEV248wNJEVYPgSc6lNlX8bArEV8YxAA
d5DtbsQzSRuzUKUeyN3C1Rmh6g29jTFxCf+aS8uopxpVtFPz7vKc8aExA1uG7NXD2DGBEElWN3oS
qlC0bLTwMlJeEjWpOpl1wcqhErituse/h25jG2v1UZ0ln6LeaGvVYOUXxfK7kv2AIWjrQDUvmrQu
qxDhW2F7WTGlcdliq3LsVxlVpfU+qrtG9ZCMZk6E+/wtv9jJjFiaN+TsD2Pk5M1KQ+60qDuxgJMK
gWbZ5LcSwg0w9NddTC/Cwsj8BExeqDZW/UBVC/Eykpdcs+xByArxf//TLHoMnnLDtDUXou2exTFk
NcKtU3enuq68AJWzY0fZjVcwifJFNEp2kd9/KAdoo2kIRTFAExQDtF0FuIh9QQuNCSMyNcBQZv/5
gSpnjk/g3yWSRrq0d7zNjo29O/C9sZwAtUyqkbd/AKwJubuX+kMVL51zM5iYXgbJTyBMjRLNsks9
R/+vLO9/86sUpZHKggPXPcZhOGceXNwE3lSRlJPvDFa5KAtRgBftgQqpQf/3L3M2k6iziGvPoF/4
wo/Fs8DIWjhkrCTeCjGFR72IrLDnwpGR2eDO2F6b3tpQyTgsNVxqSvqrC44NTD6GrlyyZuhRMZL5
ydr9bKNwLthYZKZ2KRy0kbKYoKpXeqNYweWwoUnrWAGPRC5ZsEhxO2Fr8lyCUGy08KMmc1DS2Aw2
X4+7VhPuDoT7srfQfSG8PIeoL/bYGroLn6p8ea04ghR52fcn8gQWi26cJfeYrt0aVxhCIZ2LeBIC
v8kj9oJ2arABJEdPECkQfqszDnIIZz8Gd3W29QsCFaPaHlzVMNHP8V3PGsNzQesL7+hsboJNKyLg
1rlfl7GxorPg2iqDKu4aKORiAtmB8sAxEfQHD+csUdQriaARriIufhzooEW6lkIOEW+JxUhfa0Qb
s6O/VOsCizgP9mjLZ1YbsIpHYkhDjyRj7A5hg68mZg6/1BcJfl7/36XDKCoUqZTZxtdCcvcDQTWe
/h7OX5PGMwLfwth91mrW+tBxEnJabZTV3Y//s4rgs/lEmZRW0XX5IwdG6KJt2a4U+tlNipxAu3oe
GRxmXc+8dwyVmHt2f9+kOrVEGQie3unhBf1piu9HIsBeVGp9PTxY5FQhn9mLXtaeW+tWg/MTCveZ
sc93GR/ALb3ojPytsFknsf8UNKH3BS5muylDUJOwwVCmJGZOK6loPC09QYM9DBCqTTqAxgUkyIj0
A5Ers2PH4fLiMUWj0ZVaZZpkP3M4oVuJFskCpiEy6bljWgkLJQBqwXM7czuqBDM0G2EzS4KwC818
M31kPqhrnSZpWFl7hgQdPqusFhjf7vXsVFKkB/834a4blmqWtLUWy6lEg0S4YRTm5Y/u6kTilt4J
Ed0zY5PZMY77MDQOUKfkPJn/7c7L+CW4qnDNeWjqBvboUZNESp8G9gdQ8/GJv2bnnrvYfkMNfYpQ
aM1+RSUZfDueypNsSgodNWqj+/NrPbmYHeQFexYQFWA0xJVgAZppGAH+bkKqs378BhKUUvRIWiS8
tj+m139qMGEmUebeXWrLfho+SoKHWGqPh4eZVzGVdL1qqM6CXnjBeJ8TjB6SSO8uqXfe0LBQ700E
u8cHA7lT16iuWFYnd3oUSnWZx0ij9h3zQEAlAPDwmIEhSwwTO0aFuJqa/kIpHIosujws95vTbpwX
TrxVuN6Ng1SlHHnKSYBmGbCFGMxtSQLt4wE6LH+MXSs0OewaFy82mMnS4Q5dAJvhY3yFtlRKV3Aa
aM1bw3yqPhJmfBNlOzGrOhJKWy8uu32cyPIPng1EMNBknCN1g8fMu/L5qm46ozKW9sT1JMIlRE2Z
fCJYdzDBGicQd8lenVn9NiuSQDUZtXlgvnrouJm/dO7tIzk4wCOEtg28t0RPLKRmTnzkntdyiAzS
8G/LvYciGRa1HcLaQPNVmVPKGR9weCAukTrrzp/fgRpAI7rrziOPdAGBPO5k0Vie3ApGUDArF8Pi
PjJshBf/xdU2iUXbVt5lZA2fly6a67OCaHLbuKMNFkAyMa3mLMNE3xp4UkcEl/8h9pSDY0aVzHE/
nlvhNRAs9DKDqiEKAMLDG08vZH83zBt98QwCtzbsB7Yygx7mEVJ5w39QufK8ba2EvxIvnDo7FLGg
osMCPmRQ+QubE0ezbCphc5wcz9hybRvyeCRIgnfPvRf4TNtHPjFA2UtMFHOqoKFxo/pa5W4snBge
hsLNzW1nMlFD4ww3ecvDpG5bSEPQHHe7UpLT9+68e/Z7Hc9ezH4A1YVOGmjvBBEop0nd3vPm7eh7
AsP52+gYejstr/HfT1vJd0SORI+ynuomayzJFeS+YL5Luh07ln/wuCM4MfslaNfp0i9jmGnMY0uV
KG5EuE5uWCfUKeB6Dql8ykrdMiXQHV+vymF/adJ6Lwid3Q2ezF3VqypaDMhWI+AeK+HqFzUxN36J
cE6LWDjON8aLFcIAK+YxZzpBqWGmmOYOmhgaur6FGJ+xAeoRvrRljodLGnCgentSVrCa3uV7o/1/
lSSQFolJCQwMtivIi5e5mBqCgMYKVqM7A7UFcTcWjnd2Ven3tyKvHjko3fJxeC/bgd1v8CxdJFWf
6mwvEAZTe5MYsK/2Fteii5UsYnjLIifTCrekjRb82SS3WNpz7vnishe7/EpjvBeAv/QFdRi9PNfh
t0wX0yTl+S3LBmeF5xr3y5EtXPJb/3so820yIGq2zR5TjzkFZGrUJyCkVKhMWA5JkvmjzrkUauoO
BE7l323SKHnfqfGlNZ1kg0t5m9gNzn+J/rWb5HJsfoRfAA7dyQPMeX2xjhO9IP5pRy+NDH67+PTC
+xN6R6lVjMkDkZ0pwb7lbHQK3vMAsM+FpDN6gCBFxGgO4SxEUZEZ8UGqSjW/ZPEL7TIxeM+ubSUh
3QFWlXhLuiG8kWNaH5RtZ90pHMmIjD7V1/F1RT6D385/APajCdNPvqfwfrRyyYogRQAljm4kO+sL
p4IE3t51uQo1a8DHlOAJlRgr0e5iHMfmTRcIG6+8vTjFD+I0XaDi+EyZnk9OLBBZDZq6mPirQAOh
krSMNXolsizph3mJ5dUnLH15XRz0mDmg0tngofGQknR66rAVBoIyB4jg8RP7DMTEr70zJO+EWemd
CfKQTLXx7cHJWOmbTnr9+CsWtR0YGk+3p8M+HaClKBl3xReSqeRTXdJgVPJLz2zBUpi55kReWjoL
x4TAYcST+9sVQf7OLRijFDAB56I3JkrnROPnQt5MdeKoT5EAt5q9ZMFaRgD8jXLMQDRhqrbaZb3O
F9H2sMvffIXgfv28rrugnK270kMKcuvHuY+74N6mxSEQ8cJtEqa/oLz/wq/yKN4e6lr/3Tn7jjfP
YfiWwvhDeQUejbl/B1hrdMC1cYYcWLZ+/RlvGS2bFOW+Ddc6ULl7aQY6sHLPZUUVPl7k3fDweaLR
BNP85Mf6COQxeS4Ybw4minj72d9Cn6GeKG4Evz5fbUXpLB6fnaQMaDr9tme4WEJMgpS3zEteY8Hf
0XX9Rhara031kZW9wo25uV1F0rGF2DaYhD+b+8SlmZ1/GLEiB6yY3gaowcl0jcpTMNuJIxt1XLAR
MreACy+dXly8mcXPaQkAbfxOs6UngJjuaee9mdgkBGsbWFaoFsFn09DN58p9tMJsl0QBqdpUbOr7
91mKj1Q4ZNcaGhk2qcbghQqpNU4zWnypxo/PUhIPc7pKetqnOV9ujte2dUGRWT5GfS/YE4Ix+B+K
UU+tTrcLGmZ5Up1rILFFckDi/GbXYdWAXBtOx+tin4c/DNzXcpZQGjK0GH6BEjyEZh2HhbT3sHWc
J5xbwkG/pkwa1/3owSd0iN6g77L53Cn10YFsTKnm2M/90NLEUy9qOeulfRLp+IE/jsQDfO+4QHHy
rbHkUaVQH1x7QwWNIn6YKCbkPKLRX5zho7DeHx0gIM2W/MdZ4chJnrGU14w/TZ/w3sLCkMnv3Gby
ERhcGFqblljDetWJ4TphDvsOrB8M6C7RRJhpPwn6MkjH/Bv7D5G6HrsvkaGFX8+J5yw/gRUoSfW9
dS8AfWkGddv2nVtaD5ICqRxQM5QjkhaT6sIXJ7I3/9fx9wqPs/LBkbMFBz32/4JQ/IPG1VmMWwtJ
jtsWr5YGF9olZkfps8ZFRBmrGKrtr5wlJeNFzcoJfJ+pBzy536D+vBZl16jP5mNHrYwdI9YK8IKz
hkTdPOf2pTH8jB1JOq2ESL4qzqw/dPJx39wxpPJA/9mIIr21HPBQ8WpMr0vG2hmSb+2U9x3N5ov3
Hdp/TzdYE/FiHc/bJg+YD6VlFb1Bijegf8YDd0heqt4N34UstK3aGeV2+IdEI7P503ovzHqvR+e2
Xg8LRx0BdRsT/ld0r74S1TQ+Fl6onsCRHYeBcCqxAwF9OXpx9b3fbvrZEozfebxSvbcb12+p2nRj
vHfBdmz8id4sRTC1JhK8jhBU2jSXqQhkc7cbQq3ekjnAMhidMoFdxquWODFRHASVd1yb/98Hnz4a
gOH1zlcWMBIZRkmG9I/BDjO11AmCrmSsq4Kga4dT7QmGW7Dw990RgRYYPKeBT6JsaLbuv9eN+Ayw
/Z3QGZRMXKA3JOQT8F5GV+ERzEsJ+RAT+QjIPFFsttYFblozM7BuQ0RvYm+5BYxVsPXNRMdtf7Kr
ZD0YFUjTrlwoTwYdctrWxy46rm5hPsIsT5xkZ4xOB6nE/sStyA3FH/33BBsKm+txBj3dymuXNa4f
29h80X5HcWCztPUfUYG/P6TpKaVucA5yJv8MSAUQ1wueDSFez1NEvWdgixBIvZcog0SzFJk147WO
H+XAkQktdXenPyrBm25z05uM8gEkQeMiozrg0Iy8GS0GkKHyoitukJ3TW9vvrPdgRDsInd6PAqdh
o3/l6+x5ov6+XZPmkI/N7WfnM0i0zbwxzMJwcPaM0BwYKsvblaijYVi2GGGfS0J8bQ0qHfgWT+QP
SdujSdoQ4EpzILue7GN1JVoMvu7oJ5RDz10ygfZxlaYLI7ORyvVoJvl2Wu8bcsvkNC/k44ZMaKMW
+WI1oBXCY8LFHIHcbfG5/qDw3v03e/L7JWWgUXXBbZXJTVB8bw9gWbt+1h9GS0IHSnsdTOi0DdCY
VICR6Ij+CGSAXP2th0ZRQN9fbeoyqb6H5nj6COdqw/aq7Zq/a4BBdz9Gk7K6rXdES75SVGTEaTu/
Iy/Fod5Fw9FU7gcnOrqX9tujkGF70O+4mXBT8O1praiQtXW4Pkf17Tehc1+hZ6jNW0rUQrwC84kZ
XGryOGZ/azY0chKrpT6idRV6Bn3XLx+KEW0+9/U9Z3QpjZD5Uf7wJgdeypOlRlCj1zBmlOXS3EBo
OorrQC7hOeOlhnttD+8N8n2gyy/gE30JU9zAddSYOaZkiOq2VDxaPVJO8A/yJddvOabRkrniIhoN
cNSdg5Rr8lqX9HTmW1hEyWFMUo6EDtpD9mTqL1lcUINIKs6Xb5ygzZ1K10L6N7Z7dZkm4z8uMovX
7x5YeZ8SK0qeJsEy/u07gl6Ne+dcd1Vk88zTf6YD+xvVPu6xC9SY6vMO2Oy9GlWS6MbcaYdb8Cnv
0YnmGGvXgVFbxfWRDdk7vvJqLdFqZod4OcCuF1vr+JUr0WYRa93WiyAlKOzwfMqlm10/Vy+2JPgu
AJE3SjMOjYShj4k1tdCqTp/OoyCk0QmjuAipNLKlzUNn+Oxrkq0lwAQNtrbCp8NdQux2cxB6MO0S
potDhV+NWs9p28naTjs1koo2vJCmbziRhwaS9lnqEwCZZwxZIl9BSjxWfPDiVcBB+qG/iGb1gUA5
4XuiO7IExGs9diBs6nTLuUxa46f00EruoW11lSCscfR/FhAGJmL7DKNK+gRrODAEGx5FODjGow9F
B02GgpowXH9KGDGlCnPfrTMwUYXp97hqHX54GasCfPWNUfkqxNcLR7gN3Jio2EU2WonF7YsKLOI4
iemuBSoktCinRHGa1thygIN8WHDBGpWqr2/8U/VEdoVEUMkvoaVsYBW93m2uiAX67z6X9tW5CbId
c7DEsCy4FHjgnZYgOmZbZhDGTK6XbEmtVFtTSYA/uQQ1tIXoT3rErUeoZKgg6CxBfysEp/UruyvS
N6P60ZWHQNkpkW2WsV5OBEn6oELSLONGk6uIMkKpHKK3PXg4ABj4fdgOnOCAmfy139cUqrz80Y8m
N+UbzJEuO1L+koJT8yB4taKeo7ZaacYQP9wptix80ZA+erEz/3Ltkvq7RvM4Cq+NEGJ1VQtGy6T+
gLFEzQ50yAwQKkKjTSoEltX5MQGFtniInsTCZv9Ay1NWoMgjsbUnPFTZkpdg9Vm5WiG1dSHNZj/j
clR/N3kokZM2VYKTFoOPUoZEmSgTqg3Nxv3T7I4jCuZitpbZZg8CgLviQu6BZo5eVw+/PV9vnmJb
V6AfqvcL8WjFTclINmQBnzOsGem4Fypx7OzdjNnnWS8aN2J/mRdcqijqUZc6V3llqiy5w81yqGf1
548L6/0vR4nXw04Jua6vPEFELVUFgiZfhRxXvXqjyIp56cLUH2ymjQcwJYn0SGlnyyZhzCACbvqC
QM8Q0MJF4aKbFxrWN1+QQE8qvQDrNALjvEMnKZn5cYA271kQY94H5cyRvMd5vVMRGSkZ02jW1Jlf
quWto7FlMCmaV3sHAEbhJMSFCLDU1sMwLbeNYH8KaqQbu4mn7UQlHGJPSOk9vbzH7YAHDi77gNET
BxNqUmbpnR9QpU2UHdVybn4OtitBWo4bVF765f9rbPpyg+l0eXS/BPBJchdm+tD1cnTOSzIwSl+d
IbhM+SiVEnT9apWQU83eCsey7DeojuspLCz/67vrNRDLCYBznLnOQfFke0LZAvcXgjnDomEOdrgN
Rj1RRjDdbFRNjbdRtQWypjR+Yf7RsN2wxw0/LnEl9kBCAdl/2AXa8nMsF3/VH4ecQJJyrVS0RMdw
FrE2jz8OR6bH5Y5yq0Wa/Wl+g+K8fAssOmMV+fhemZ/x8pbpsb4ckArtGIbIvaoK0yyOnopU/dxI
R6wIhcWZRreqXi+/NrcjzEOMi5qNoZFJprJa7PVztiYpoopMUmKZbWatwNOY8qU1KmwshRKeF4Of
fIZAu1GBumA9ErbZdrmDWhMpEXGCnqfMyKhQjHy/N5v0o9dtNAD5+A57afhBLg2pZnbLnmg5Hyp1
TMjwvduC19a7T9GoRDRZlDqz/rUFmDAq1484FZoVw5xTzZ8DJUbw4RMSZAIyrm1HoqysjFEUn0Im
La2pCSjpJlrG+FyUhu94GngEzafKylmuyJB2snZv8PjWzmG+8pjsCuSwOr8geFyZWBRAUableurK
Xnti7Noms38U9cFl40Yd/PQlHAu/usk9/54XY9Q3TqsFW0EEzlulcSWt7ZJPnNwfwnmEgtOn8WHw
nTSd5IAWhTta0U57j+x72MHzVzBgLDMAPC7Wa5nV3bQD/WpuUDe42UVqMLfzlSPjW1KUDf6NX7eW
FBucmX88H+nXu1Oz99riqIKLr3a1Bhje7e/b0/xHEdjFamwgUrsizfQ4FS9iXu077ToXyAJL5P+v
705l/fNKcwbZDH/3paJFq/X9NUmb++M9uT83YVa8fOStYRbTdXSrqnY6i+NYbHhRukApERxWiMep
CR7lR7b3XCY4xctRkXtWLwQqktegDQvtPnY4DDwJ3P5iWu6K/bArsR5xbEmOx5p3voYAVpIuF8fv
nAB1Ub5DWadmN30OMbnHTyYOPdoaa41NdMCBe/TgHwZ31lNw9bOp2QZ1doMmBFWB7Q5CrTtJDzLR
Blin7D0N6zZg1spBSRMQvCqxZ1nSVKmxt56IBfX3uKHVG7zA7capniO2VouTkLIOukNctirmsYLv
fTEj1nLQUhdATx1/S/yqrUH627l7HkF5mpGhrpnN0/DvhiEFYgmFhFCBFuis+VQdjrbgT8U9l9LE
z78VF+hXfAnRBHaffV6ilzuwORNDnEZhwDKgddC2fNUveT8WF0GfhTsW25OXG3GaE32W3ZjZU7rF
pAVdl3TSOPvDr8rb2wx2pvB1/PWBKdCsIxC7HtNcvh54pLeb7wwEzM4P+9QKPWFAYc+ROy7kSX3v
dPjLJXIEUO5q6Z6wyJR7e2hvFE+MWJzR0A6jVxeMM2MC0FFikUKYBwpF8eHd3cYYl+jfvPgBQf0x
mUF1GXf3EAa9XWnepqmimG8yzowmqvsLRld8Y9GAbMpAxW2tyQOYaFTyCyv3GlBe741TuUE3ih7T
LEqCgMJ7D1FDI1FQFYbiZqodicuBdAkPMy3C6x/MPbO69kKM75HbgmjLwmJp0kbcyP7DkalvdtW5
04a4pvOaGwNafASari0HWNU4mfFc+G5yKTDZre82NigEFrKxQBfHiFp0p6RA4IikxNZW2B78SWJk
Rt+RslwxhAOMdV0XYjfV0jCxoB6ijJWO/RAOEFa3KZj4I5AmkaC/YNtUf/Nu+QYjlCX4LWOwCDhE
gp95pTEFQ4XquqeEM8b9A9dfG4lo+XnbXKGpA+4aPGRMRalucPMumIpZHCb0lycDzv+UL9mP74JQ
LUnNRX8AQ95ll7GRj4BH3KjsPjnvpiSygsWzJSPKm48Blw9kXM9M8YU2XjzJ7GIXYbgqbrZu77BR
2fyOPisGYAeKdr9wP9Yu4+xoSA6jdL8uRH+VKAbLn5oG+U1uG023gJ5GqiI99Y0SRfrg/7B8ZPZo
+fkoq9hZEJAFsl4d2rK7O/hFQMRRSFsu98U7RtNrIK8p1/c8IXYiQkP7mcgSAUBv6FrQzbmFG5T5
z5N3sHCjB8eZeQwZNs6QWiJVKbNdUOdXFA8eI05snAykzs3NalbH0LgeGJ7kJHOsYLiXoHnVeYOq
S9h0TuWRWyXXqgnn2Ehjs/HfIw98j4T6Qg9Q4h2bb+DeGji8kahbvtBrnQQarHOFiGf1nC0IL4D+
dmo/+VJkeRYSsMMJZmMqBpmFKoWsFoZnqcHrhh7/qh5p9p+L8PI7kHo90QDAJQAwtjGVhC7XLJz9
D5XkCDN59J6c5ETb8SQpiwrdEhbel02DwpXxG4pVD2pupQUx8oDSkR7ZjEUTzJunMRxDn1N9OnBP
zeTo6mG/+3z7qxGLl8llARLYIT2K8Yi2DBDb6i1E/5JyOME3p60hYD4KEjhjvb6K+gaLh0Ug+dRE
zoJEXkNFiwT9IAH1bJU36iKuWDetSQ4LDTY0zeKGCYZQdWwlM2J/Ec5lKiiPZa/Xr4aWykxPGqZh
inefzmSFosPo+AhSTz6krmxFtlQyUHWOXCmt1s5jOvRnj6FbQqcTOiu43XyYjAfeggi2/zcnWD/h
SfcOq7MRCTVQkREsNn++mhCLK4feHllnxqFSKeMvxxH0EpCGv8iJju2ZqHgYHi6ucgd/Pgg2ZMZ9
mqbgv2RygYDKpF26335fbXMh/CpUy09T6aIjkcdJK16izsWuOnFbIxXJ9WVc+K99E0kzhEqqGetI
XuxnvmtxnrDJkwP47SzENeyNItxolznre/hP0PRocfkDhQqtbW84UBE8otvTlT5bJA2DOUl3GPEd
wz6oWldt8XeFZcJgNBiBhlGp0JqO/htxG8zAuw4JNuy5Wd2FSZgasxjWxUc/mIN/M/1js4ekewLH
OwCFM1e5YDX0xWthB+d4zgF+uoKUWLYSQDNi6Ifp098vfl8TSo8JeoKhEgzB+GaySEeE4UbdoXmm
CeHjGDFtqiSi62tQlykR6mzEt9YQ6YaYyCYWu1TZ9Utlws1EcQrH1MloNjHFlVTJaf4qIaRTgxLj
9AZC1NEww2PBuH0UZmPhxRwu6mDebQH7KcM4QPgyXS76M/t55QNfP4oRnuWToYW8YmXqTUiPZbID
jEDmVYgbwioRhnU2WzzqLEQp9tbsCHBAxUANO4cCUia8abKBmNnWteYSgd2IQoPUAzjpZjxhljEi
FEwuRWfAEEsMtVflQUy/P3R6kJq/kpkrgzihLDAmqdBt3Ekc6Q1Tqxebq8yzWUdLsTbhl1NUGq+k
Kxe7hKim49lW9SoggWBIlb190oYGwrJqOsmslfKS5dUQxJONNK5m/ppsX7NW9mkNtL9SbkkneuZD
FxpE1aFfdAB5t2T1NUztKx49RtRuZ1bAIFBPcgSo7cgs0new92cWTkgSUsPNjiYgMnfyZLbJmw5W
frzZpUiXcKiOIXSvmcXiMf9sAvAsu9rKU0vLu2clRXo1drxGoZsFUv4ID/o4v3sPBdZ1hgo9o4ev
ET6Z4oV0LlpEZ043iBwy6UNxlfzvYpzfqVywf8cEqdA/+csoJwbe5St26ZPYCKdGuhbUiobjt1zj
edvuUMtMTV3C313uULehqomtQwQ1oAQ2hYjh3DNR9PeXBURnZ847PwNa4cjW4UBuhiUF2mZxCaq/
2ziwTjwO/TR1Koh33brSDRUiJLxHSdgyx3IksryfgKxW12lMfIKtGO1ydDkPgj919wZ55FpvgRsu
Ggq/sAkICA0tE3lrwVbIHbJaA7nrBnlf04AAfEJC3lm/PBSq5iaefyy3dk2HKwbgWsf2ZlN/F+js
ALL2KDDdNmgPV8w8y0zuaJSt2m+DzmUx5KXGVPcdBLYFNl8tpjXmazAxAxkt+KAbV9OHHbUYp0V+
HBjKNPv/Y7Q3GuMqJcLuf+MeKd+yYZos8memKE90Js2yGU64fGPiWrgHzglBnCVHus0irJN+ajUx
x51xPQrpAPtXZmQGMpW9WCCI5KLbRy1+hx1CdLVC1l3W5VbTLNgUqJs/kJwG1sk+oP/akN877nNm
M6/i2yPD4792FSMDZZgQm/5xCEh3BcT6n+c3WJbcQicsKseOLmStkZi5WAD80ab9XSa4ZETcPNKk
8+fVmedA2JIRurRTbjhgTMKGSOtpqcUIqRAepzjs3V8lgA0Zw0jvdQpOXAcrsLxGy5SLdxSPGYty
vxFzuljNIxAJxfgRrZVCbXDsRfMO4bfshb1p5UhjoPzmtEYduxHWq6NE667F0YMfTlP0h9rPe66g
NInSAl+gsLaVMPCWr23pHckbaAEgYHCBScp571xx3bFhYBh0bB6sbRcvLYp9/bVwdF6PxgPzPx72
StzDwQNd9PzHfr64rJh1T9ojh8jEwNE8Z91dzmAGUTvbxU3g3XKUuRdw0jeFRDtirzhydBvla1OU
bqiEDSkDkWIx7t9Q4PgRfIIsAKj/4xFiThy/a4pHtvZ8v7RPINDd+446Himp5H+Kf0wVPrRdvDw/
KmIZhr+uFOM1i3XrYfrayyDogF6S2IZr7fTnuPdgR1ogCwvPjHoOeSdfDJrMxXl28diaw8Q+69ze
+cScQtD/8jideix9fq6cSMe71KvkfSHSVFeOII6cSU96mSV5+MmylE06RgXFPs9DRqP+Y4Zrtyyp
J+PyBwcRSTA179bNpZyBayThRMCefUmrbPCpJhkPjKpVCMkY9hzniAdipumCuV2bKOuCedRwKgCt
9lCeB8Bsrl+hOftlOb2kPjRLiW3k/wwRed+prkCpAQumYkUWDoq1S+lhG1xS7B4GC158bqYvZBSs
Z0AMg0Y2k7SgWai+QjkcAjxdmXGEWQIeHYb6elk+GCLwnOF2LAlsCfZY1SrphvqlTH5ANhEI0KY6
K40G0ei0RQ9yi2E/uNFy1fs1AGFwH5o6rSZW+9zqAbm7QZLg5SKSwVhz+2anSu2evHg683M6pLdM
DdRNoJITrnzHtBe+xKytlzln9eCuyvzMLdFZ1RWHKUkVgGoNuAgkkk9AQn2rTv8OaYLRHb+IlWTH
zp+6I9MOdsqMaoYjzbpu02MWgp6Lgk0ftzHSyiEgKDDreAjxpIQYFVmfOPISyBkqZZl3aCg8nMPd
Mi6svLPqh1RZnsZ1l2XH2SqsnEVeqbFdHs6sjkQXEiYbRYooaCjStUEKu+9L71oTmerhISSp/BjG
WY1iVTvwCN6BeabB+XgAXU/OU3kamfxQBEkf9R71Ra25KcHzio4ZD3PuQ3fXRSV2SJqCoQomT+8M
MuLSvDHqTuBlxjQEO4gHhJ83W8AiIfylVoFcZhkm2DVLq5TW9yQGzAsyo2WXjUyuwAOy3B8ehqxI
0FQlsFabk1IkHs2em5JwxeobxByPBJ6crS9NR1PubjEXNvPd1srh5l90M6ibCmPQkkPNdzUkG19w
DRtO1sySYAMUQ6aSmUjPrUeAb3GtvraP0Fd9743yUTc8tpjKYYdQvEOXPWnDdHHkHH6NNTpcYvil
50BcQYHzX1H3Lgd3WtSV7HHt+Ubqe23kFZDDZejuhmBsjAi4KIiGPRowKnoWT0Qf9KuIQnx/I0X8
26wVtrmqIjyLM5lNJinNb8fMbUK53lSWhcWGWP5WX/TbG0p+346r5J0j9gkeg88usF7wzw6Onxvi
FJyCBekh9JK268pbbrQX7TeTYiCrkgaasTduGzCkP7js6X2EdOSYLQGJyRnA8JnFI9L6OaRnpvKc
7gYGe+VW4z87IZuNYkYxj75G4Je3da9JoQ7PPucJZsHhUq/21SGmpa+wzL0AXpOF6eQ2wSzG9sfU
UbEIhRLGbv9aO7x04MeX86Xo93425BuiCrQkdOjQJVvn8JjNhQF9lPcHYwTY4EtAXOfTAR6U8TCM
QnEFFd621A+UJhtzPftzNwXeEwFGSVZmfzFaTMP2RrQ1HGNxqTLsTyhNvhh+DMJKZ968NmH9rRuO
4aZ6jWjiRCtPjVHBGbmh0qLD+Z2+iXWKFtV2MKsNSsEjHFGXCU/003mvF64JgqA9hiFfY0vKCb99
UZGe7oG7kQohUV4KwooT3/Gd3zVEeBjNQuhewRLG/O1Xz6GzLQR4VNxQdzF4KQ1Li84GMM5b1bxk
sXvP3aQeKIZvqkTjPq3OmP7JAwj9JKzTJb9+Q3mQPgODN6PQjHiGzUmivZwfJhv5lMo6XO4em30E
55BHL2byiC2vZlfasrKLrpZkCC3F3O8kXsqXJjP5qcN/Vj4UPvo2lY/lNFWoWRcFT1PCIeMZg1zh
R/QOgb2W8qHL9uJu8O1ihJXn3rR3MQR0jRApxh4Q9ecWJ/eMkHFwV7Fp2qbTzw3Vw3umyeap7b7U
YGHDqSXBytgU1X2pu/MvobLeIGvmOckQANoYpshFcbfCazw6537GrbeyDyUIfi1ka2rSeW9VTPp3
FoEd73/izIrl6JJnbrTB2hTcljpgUSWxf/xSe15U/bcqFwhfN5mtQrc6V/1KcEr1SBn2/zKWC3E9
Orr95A5NTQqYn+dU8o7dnM6yRzlxInc6ylLWqXOfxPvrJ7iuBijAnKtzPibyZztKfkqnHt2lRnX4
iNb2TJU9LFBbViiA4gvytxDIOYiYAms/vZixQ5BhvxwWheR0IYbF6jnIPpSye42ckwqDgiL3DYKj
zDxbU91miVO6sHFVC6qZSq/3AuLs5V6vQwZXiKz0aLKbn3vWFpvUoe1BMmucGuHBfMXuaQ+voWj5
duptrdVJitJcR3BuMZposMkhdklnfduyuS1H9rl6QxuONav2GlbMZjF0IXHHXu7ZrnwZOr7FdT7o
hiTwTn3UdYLY61aobAQqZgUTkcuaa5xUnPaEnEOsf3iBdUkJkUxGbSHyuXzTbJmLoxaYkH/Uad7U
vcIomNJw9Q7LhnUuS7iLCL9wpwUSVP5RYpU8G9dO0JNxmOUOIQ4OxYrfkqg1R7G5+KPp8EWUFdzu
grBo86zouWmo/6IfUiZjm0kH9AK98c2uFlhq4Ob8n43ftOIz9T3/Rq/TianNBt6Q6RB0FDvgE+S2
b8DoZWjJdrbScPNF7ElLPl8fEsRgrQzVDP+9jpRcIFXpy/z8ijMJSWVlkHplokxPmivwafEaMTw8
OAKPvM9l1MPd/B019aOMc7cpZtZc2FeDpfRZW6F5Yp0tACPlh8OI4N9CiqTIrMsd9cjmzPv7H5du
iPW8WWpzUJtlRVu2CbqViV11vL+upTd8kvnPkUpTuuXaU0B1NfRLYCCJqDtTPMeS03Te8HNuWhCG
YqJhVbBNIlTF0ZFeeVthY0YTOBL76HaRVaXOJLanLOYkUt39AhgW3u62ifbupuM4XYRoaGzGub6m
PN42ERuo+t/yetKwncjdXAkInAlUMEdkcDAlOS0fD+RfKU3jP7H7NBxuFSmk6qChQ8Dnk9dJTvlO
FS/4LpVy/5VnjSkD+7MJNeiWgY/Bfcf5dFNBdfxEyh+cI5nAZM3CFmSNePnVvECKa/BTmLLqpSkX
IUVdwtScHWyMBbCZw0Js8RiiPbqGA0dfJyOjP+DvJ+S36l2q/9kGeyzLPEv/Z4pdU/1biYtu6awy
8DW6BREfzwGMmmPxgi1q+bPb3g1jk682FyBfl9+lfD2gKuom5AfL0tTw8Q/Mg6Bemvfj+kLgzCax
jmuB13BD7i9OQlNQ/WayalDOfDDU6bF5XTyGyhjLx854VdcPciIfQ72f2bnW3WNmP0srHTQeWUTy
qXC340aUmwZovll3I12Gf3HurmnKrcnRNgISlWVMYGDSIHesPUnk/BL0qUXKWNtTpztv4+n+Uq17
m8u43PGvCX83IECusoXgOnR/m7f2WynsheopcTYo9j6kU0J5HcSoeMsXGsmOm7FMxqxWp/fluMlu
y2PF0elWgtaLYvBIgux+jN9ZjfrzvbhSQjoqH3DL1mfoXaTyIepdcZCXw2gESWrWOxpHfVSAEuYF
7rDBoa5ak23t1Ao/sdck0ySFc0B6yh3BVZvmn6VyzyJFScHlLTSWC3i2tldf3fUIPsRrS/f32yJM
62d9W/WsPgjwOdAe91gzxX/Ey2psS5Vo/f737o0/5lUJyUwjPHLPcdotSpJ7DfnT5TiTcNrcw2Mo
Z6Xa7J5CkteMdg38+5AybrW97G+i3kh9LuofFqrVHRl1NFm8Tv78xMOsReAHQR3zODyJjMmEW9Z7
OhoidEE1xiTN6hU5vptZ4RP9rFmcxFT7URQ6HIYYBMR2HDcL6G5gcACYbJNcCbpiSEUP35cm0SXl
7Z/OWIQN/e9/W1nKG7iDKMe1OqfFguRdYi+3Faj0wLh4WbB802o2Ezd2dTAY1n9uJsoyV5+7Nlsz
yKHtmUFvcWArdXxfQTBZRHBgSDM1BaT/i7Do0DLtTz7vW6T0qf94FDvqOkXgKnfhn6lPHczyk9pF
JUPy4Aq+PnexH39Iq5HJ1EemqS3fxEYl9EIU4nNWy2BiNzUKHEqW9MMyXzBVzv+hUr3j9wzu6CI7
5wmefoYFJ7L0UF/9cIfliPp4d0iwncLnrlhVaJLuQmoD8hsogUnob2ogcm7EAAU1ziAreYhJSfp7
t2+DsX6LnPBZ370lbG90KAP2g4USIMOyIPg+lT4KEgu1y68fV2gtA/MFp1IBfUwKv+Y/H6fWKcjP
lzSr6qYNlhzlZQtrt5V9hE2vkWhdAV6xZKhifrTO2+FO3q9rM8qyL+ak5NO7L1QXepCQTDr+6k4e
ytAv/ukG48hosLVlKlKWEsxh7pxOB3JerMdxK0WqnKZ4983MFRgz2hLu7G1U4X/kwmWehALC6XLE
Jkj8h+BK0lT1EpAbSXFSNGIm4K0hwY2Tz0fsN4queSMCrD4TOTYzfXpWkbkchmuLQV/39lWdXDZB
s0LNk9/qEut7AnJGIQ3+ZN5K2KcptNjMinU/4+vEHhnmVDmnBCqHyLqY5ZZt81UPnYGPHUfXKN6g
sSP+PTnGCjWb0iW7M0p/hEp/7/vnpAmisPLWcuwUtYjrT/+BvRKevR3qPTJ9nqYqqp3cIrY+UWn0
DqucPoO3vqoigzij/jDshQDn03VbPkSF80yxau+s/yiJ6ALsEbAkab9ptNh3cJze+ErGt8Pkq35V
8H0DtoBKxqCF7CzLmeYFA3XmClMP4s8wmltKgITJpdunnDBNdzkIcoISf8uI3hIHQRENVbRGlym4
aMSus5Bk5Eg0UODHaIHXbySSCeZFZ2ev7GGgT2fYjh0gMhIB0vuiZCbtRUaVCzqiu1tngCkf+sBT
2fLfiBLQP6w8VtjfJMf/lWSNfwISjco/l5B53j0kgZhQouS48cNyPLZMEM+E+r2T4C1T5EH2E2g+
E/RhMcu54ije+Ups5JaEaRxRT3sYosVkIBdpAiSLqto3m8d1FBlTwwY5/BwPeVW08NLy9l7Op3UT
tIcxU4gbj6i7gkG9Oeo66Zl+MUzjk38J6ulXed2KXDhLyFB3x9NfuT+9uYNxyLxn6vBA3RnH8b0R
dFgTn4vyYN94d1qHR/ICmlNfIcmjTdHt1pAURZQmz91Nr1Rsa17kWzBXwjWZRq6RgOvnu2rhI4GU
aMZctDcOjQECsQIVVLaKJj9m7YoO+aH6gwcjP+eSusNlSvoojV3oT40SmHr7rWFbWLPTxP0RWSez
hW43DJIzdHZoRDQCT+bBGBUartUkNRyenlFGpmorY1y5zID4rgO7DPDvk/o9ZQsxM20TtCac4NSW
CF/Q7NKwWujDNc0gHI7PAsQup0Z8sze4QiNbM9e2bNI9BKhiN64MR9TTwxQuj//X6zQcLwyHeMCt
L3owS/2YYr04mQHvV0/Hrdj3sPBNBgZ6+e1O5S2v6jPvvC1VKmXxzB5V83j7NHL0UFI9mDJpZy+3
KTjycFISiQvr6RNa1TxyT3jzzyLaGMJqR+B1HvVWFyoh5FGks7WpXG7WtoU8IWlbWcGEQOz+m9pf
Y9PadcbbojJD3oAZTPlHYtP4bzZz0IJ7NH/Z1eFt8tC3Au0E+6mz2HfHS1FKHkiilB1I5lBGi3mm
LKSzZOfxiVNK4IhYuQQdxn9FIM+zV0eVMJW2cAKGRqwPI0LswgX7HL+ZwefiBLr15OXTOtObgYbQ
J+ey1sOqQcgXcZjRKnvC3sVh30eE14XDcM5eQcBDVZDSojI04D3M0cpBkrag3ua9di4VFOlSrpue
h85YpdexpNflYBlhUUVCF/lNeCdCtQ3sK7dRf5EXwasdwDJamx9JKK9h64gK+jQEMkPP0XKKhB/8
d6X32IlKds0TuUtR9EEUOdO1BrUOE9vwoc+fLXcVlI4vfRgLKObxOpNgD0S+0mqCRjh/AGdqoaSj
7tuH5YP6ig5YOPeck0rY8rJlgeAowMix0nK8LpREoVAuFtvWD8EY8B9MALqGqjIkVYU+iYaOrgaK
PWuPZ9NpsZiyqzosdAsCeXrn97YjpzUUq0cTJK7RY3IWt5K0t0R0gFPotS/8yPxN3oddugiYbqf3
u3v/GI7885nAmcuxL9h5eFJxtuO2sZuVSwfB1fEP0SshDVKjxEwVaCZGcs6CLGjXH9J+qrhhnlML
ndk9M5x6lsGgJ5SvPO6/qXEDatW6oTBrXKFRZHtqxfLDQUun6/2HyoPTxkxMcNE043WGoCHzQXkR
d1pfcaApCSCAjqORv4LareKrLnXDndkix+TuXJBa/rhvWw8J2NJb35etbHb0CrSfF0kTupkiUuxL
K2SrHdR5RORkXvAx2mzI+2zjgptspbXk8qjYBP8O6YVc512j57TO4X0PsTd/zN71JW+Myb5h0vLQ
bXZcITgJhMluGfR0Q2JCnIMquLfWWBim9wFXLL2XKxHG550tkmEnDGSzBHHGlJXGw5ts2IcCoIrB
BeP8SN1WepSr8KzhfIyiL7XyjgfhjEDSxsU7FN+K6cx1dukdccbEbqR5Qt0HFeDK5Vk6DDzothgO
IFG5qpVbjSWkap066oQrevM+Fg87d/5pvQemyuBxfYQOwBWjbRSW1HUoAHBGB8i3l9Q6Lya9QBAd
CymAx++OtpgcMzLFdWQf2pYAoGwEVHpfNCqnho8ze4fUJhNMZSn95dVOsm2E8/VzDtpeQdagwP5L
SsAu/t3ehxsp7GtLMKnWj3q6C6hT8ycsbx7HznBdfP3KblmlrMCxqQbG4o4/smjT3GwuR/Y80YaF
7/al9E6s3+DY0XeR5HWQQcyXJ/ULFri55QfzT9yE5hvUjIezlmpn8sykEW0zyJJv5fmQoh7z2God
uUSjheT0R80C8bZcGj/0n25Y27gsCUDK1zRDah9ZPNX/o9ZHNcN70ff0rkwo0JLgBLssKCTWBE2v
SqTvk3g+rbKnmgGf/elhuHFV8MX/mwLqf3EeP8NUxALhDQML3I4dSIFmuO+/anq8uHbs72P2x21B
sLz0L+UgQThbHNVth2VpoiPWMjI5HHESbRQ+A6ByryDq5hgQzO/1u2N5RRq77tyUoh4f6zrBfycM
s19QBIrpoMPiqQxk8+BOmxU61kTrs1ym+M/e8kbxz1u4447L1/xWnwZdaO9YQLRNxJYXi1BlhUTh
oaeEUoa58swQbc2ezRvvQQWMw/Mu0s1LVVM/qIw9vREV7Ikt3KpNB0FJdvsK+iy+iTNmB9Q9VEHd
EgSfPPFjrGB0joetRRE5+XDrNax4A3rD8KEy1cWURxOrxOu5kWJ7anNOQJYZor6QLgPFgcjMKF1y
m8AyywwQb2AU0MGdKfUCzWQBfjrNCTzfM7Endp9ylT7D4p1szANXDOBBBdmmxZr1XZrK1XVWbZzj
QfpB6EB/VnPkCm7xsMN3y9ouhWZ0u4xkriSxX8dafRloVFfELG9vo7dCBTfSUBpITG37HQ0trBBL
x5recQ8YGhKwiYfZEWpYgmNVmwctzubKGgomGm8zcr+Dla8q9wnMeGjdBY3XFRpKxl8NRo4YohfA
K6rAimoF6R9HU/Qu28jGSkUodP/OncCEapyFUJSdxGdpyucCGCb81vwymWsZbpoNT6j+VRHKKd9t
CBbQjvieESFJh51ERSCJfFopz0MykePsdpDH0wK/YajtEap/ilm/A/e9FQzbnYsmaYXIMfCaYU5z
bz+y1BxYzUkEPZVzS+/nTido9YUqnGW+28UtP5vZKKnSR47AvLAvbKwkAhjsEgBP+8uEXrm9O3Kk
Ic3qZlbrhiwZiweZk2OW4UhotVsYOAGn3ObHO7Ove4fw3y3Ke6Y5WN/A2L75gKqomwgBQIqsSbM0
zI2boanpX88/kRKQHBiDpAGZHxcGB9O7rJs3VokRc8/GEl467QA/4kYllndOY3+IvCukc/jVzS+w
wyFrcbrjOYw+eENGbrv/qXSLqrVopIqUznXhJmMPxWtxGA7EzpN8f3RH5ZXOnTFglZpTm4vhX8uG
u1LmXEenqLqa6C+q1jYBYU6bXfThJKZYyD9CfodF409wrmUDImRGi2cJK+vD67hd11fK6sJz8hKD
iXsM4n0k2GMIk7NoSayaTdOQtSBlt2v8aTLp3FXnKLRB75RqUiKh5olmOxM1PwfHrwWnxkZMUsjU
24oGElKrh0B2EO6uycvq+rQY4P6cxBgioajPVo9uePiXm+8rGWY3f7wY2KUNFW9rXREk1DQWgrdw
AW06KXIPLtf5+7zn7q2/dbW05pJuApYZWz48hCfM78IJOgAdekm1VnnlWwBHbcnAdAqgmblfxHZ5
TubrAisVTNdXJLoU9HXNBZBAziPk/TUaudldJtHtaOktYwLGuD9abCDF2mewCaHEOb8ORIY6mPJa
Dvr6KawqR1dmu2Ojt2YJAq5VcRlNFXtRZSCCyuxxZSRKRFeKXVckPZKP56kmV9jO15GBCnOQPrZQ
TAu+R46laaHseq+F1FZCike9KSw72/AiIx9CkxgFOfguSS8EyLGPp1zLxWbnKlsspk0qCuri7RDB
uOCrTZuFz1ZxBKMXQRuKh0kzBAUL2UiKBr8gjvQLP001AEmgKBEEMDEGG/cYI0iX2mCXXeR/tjaL
xuAH/7dgC8uPoRV/cc0FeHRcneMqQb5/9tens7LSc/J15hj2aMBBRtqOrwj5JEcPI+26vZSFOOoO
IgxRCPq8j2921C59ECgsqINBX0UUdAIQQB91c9w553RSIdn+5hbA3ewtyREReGbiD5MjLQ5DCkfa
5FfprSsJd/TBWM2Ov7hbT5Adq2xPvUws/ajFqerZLSSTtAkiH/f3IB/av9sqNHajWodOIs170ByB
rvj1Dqtg7EP0m5Af06bsXawmQ9s1/IfLHt8XPj59+sC875DKxiSPyfjx/kcKVvU7cWVoNMyBP/KG
hretv4pWc5y//OOFD8PV1VXuolYr9bCDwtWMwNuSwR6mM3F+7Z4IwGT5Ze6nfeOy9rFMdAo+WU4q
FieA0i22mTT2eZ9Gkom+qbwj9SmPEfGnDaQAA1/U0o8GX5VoOEHU0YTljVyGrboHZ/ELJvor/O9/
Ri7H+wuigYj47Tijgx6ogKQVUiAB8N2ejkz5xv603+ca4QNQWmDN06fH/4L101BEXGolvJyZ2nfV
+VtUPDqaqibI4fRfM/uKK8JHUFaHoucF7s4eleFnB3Y5Mw6u9eDfXnMG0QVRK1AwCQbH43u3sQao
OovVxCSD0epxkjuAxWKJeJ+1i7zYAtALLexCMIx/LYve+wE5dmgZPEkIDZVpvjuJDwYyGdUWcJtb
Vv9NSzEUr2WvY7OfZhsCYpf7QfqDEuLXJfcnpFtMR6NkxLm8KboMP0M474RsR7Z4BPKrDIVLFiAz
M8QyNDQ9zeKVcqtwsUGdijNgizPIYLPohMwGymKlDcnUri2SMh14oYT/cmwtTIiW5AJwAFClGLut
vh8qnwP5FRaoYu7usXZJuL7/SM0/CIpLAm4kW6bDi9NorRRsuFN4fBsLJgfE9VKsGSEq8I4vSmGo
Kg3SAmVcj6Gz1btoFHapuRDDlHF+KXlQ8b1bKzTJo2RHhjjwkizbhbbgm4JVPgfWyQz4LgDqteoe
EkJPbzLEIZKJJhKkoVab+Zxyr9iPVK1tJQYySUbBulmGYhtAiQniMQ8JzVuNWiY5YVmz1fe9pOvf
HoMxLetE95WEeY9fF75Cb3V4I7pi6teE3sNBIZwW9ElVkPTL1QvmHixzsnaGfpe1lO8je7Kb6f2/
sFJA4M4nx9WMlANt288CKHyXtvNby166zagSzHWIImX52I9NuJJyOdVJIjdBl2vhpFVE5GBf2QDo
Bv+5dU5bgr6zLbSjhcCduEZzf0hPDoSyKlIvCVgdoZLMae2qVB6Tx9wCrTrdm0cv/fI8hWVU1V63
O+ulG7+UzUGpOQyEvnvHxeVn+axXrWL0odH514kJ/AI04qk/cY1eCykcbNa4wH7gKp3dj8+aeaHL
t2wtrs8o2HAq1OHepUQnPBGkFWtftUjc2I78pKMc2qWqO4+pMe+dBf7bOZiTiZzjIZ3AmabA90Rg
I+OTCtoWFG4XIOFBVGwjWrJo5AZkTupvWN2LM7wYcAWjDqK8qeT1mfSlnYlyAWq5dvM8dIXulaJ2
gQE4flw9Ze+rNPo76e6E5cmM+C0Ss6AzZhyCUIF+4vHYjhwQjDSE9cX4DxhTdJB9zg9m/P8JAbG/
oUUELjqbhRkON84fXCuV/Ie5AsrcdQDbISC+FSlbFgaQzRIHVg/hGsao/kiV1irC+QuR2JQV1Odo
oGS3rAFXMUDksneL7HHj10ZFWdNSSYFgrLI9ET8BZvbE6MhGy0BDmia5+e2AkepvT29sCMS6Mfdd
T1YV7bhFCwPr4MUGpeW/c1gXqKTfpZ0BODy6ELyd6JRlcs1aJb0cC//BPpJtkh4lamBsX7Es0l4v
D7D/z0ucHH9OPAkUakbg22wIkFXf6AnBFQq72eHzFf3UDg/RFJHpNNbfP80+Q42qzcHtl0Ujoazo
HfiLfHJ0F44JTYfZUFc3F575xqqmdMdqM9IE0tY4R7A9q+lPMaVq1zXrAgKp/jfQnYrc1rvVnlM2
44If8GokXlRS7S3hVwuYEBJm7DFEqZJYvuwttxuYRLsCBn9Z2+LyssO7coFA5LrKMsMd8sCd9nxP
vJGxZe7dWAaoWS8/FR94ZUOxYXhDBGf2Nun++dReUsV1OHWphMh45v8uQL8PLKeBmObnZptNbT9J
vw25lldoXyGTLfdzSlsAN6jJNQpYy6AlYHqNdHUIZNCAn+1hCJpZKOV8aoDlsp3bhZx0x2nf/PBf
tF3OyrY9VcT2nRlzSmdejLIeS0WA04KWPO7fLIOQBco0E0nQBV0SomljI9lAPFloW+vczAtRTV6j
C+XJrguKkMFi/KhJXPmiNBpILap6EBEFadIIClYuSCOe1is2F/W+IRzkSk5wUv4WuZoU6WFfoX1T
HMsDYFY0EPhRvBiSth7SnA0uA+8TMuLXRX8ZSKhW4Wdf1PCPVZ0wtNbuX7FuTZcwvDpxGflXSQ1K
LK2eDdRL+kCTRDrdb1wxzRLIC/rjcrclAlCjbaU0rUTP9PnFWDb6gM7PqradZ3g+RsZ/1CUXhspB
QaJfRencoUVxeuL2FHi9Fv8K6f59xsx3RjFvZjaCTonFo4pojsOfI4E+Gk2zWvOS4reiEGs0Cvl0
FCKq5i8DbZoC5MIJ5uOLD8ij2NaNcA0eltt7sbv7L0egPU/6252ft9xyauS/x4dio7r3OF1rdJHb
kpCckpMXGWDi29iM9Wyw3r+ybaPFAi33lXum6REcBAq/5pRD8iD0Ea9pna1s935MdwlVOxEwroa+
G/fIeKtZq66gE+4LjX1he4gH42JATq7Qt4KTO/jVdpxnk8PHm0w8zdGsaHxGx6Ric7XL2G8YfbYA
udkw79cA6kPh7QMkpsb0gYtABuv8jWSjU71mGN0yfhAxHxBh7j+n7hEnv8h4AxRSDhf2enwWTo8V
clwvHuOC30Ma610BSxCbZJAp5zvQL2kKr+abuDye1IenbhXGULFt/YoHzL2j5mIZWBmH2G9Y9GpM
INAlVbPnJd+ElISE3a2+Ixp2Q120nizuO9IOLpLl2z3nXyT9Z1j4teX6y/yA9v82hDOv+R96hLvv
kKGo9GH+UNSFvxcWPi5GkhGFxnzqcaEjKMVjwgy1fitjpo0YgSFLmOuC92LdCxJmMm7TWykRdgRy
YMX4LYcsI7ou7FxJas9orG0r0IMBQBg0+fEHqrLs77a+6poZWLBMH6OtMcB9EF8lYHeyxJCl5prL
i+H9JdYWH6pAyl8bAyj91xHbnI7h0KLf0HoToDMUuHVHPv1ru1+XRsnD7OFY2AIwWpY/6Mo4141N
cJV9pSHxbxlc7/cJssIAj/Rz7Zw06DpLbEY0CISktIrd5a1dMLNWFAnmMAW//KNIklY9KYih0Vtf
DJblRlZ8YCnllSw71X01tBDiTDVAHTN6l6ErDGZ2N0f0s8R8RKP4GNS9AP9HPNzzTcg+slkbWYSI
MDuElLAtCfKPgWpey+mSeB/p0mUYAcWMk+QjKjVLEJ2j21c/Cuytk1g7v0zuLYKamlSCRH1hcSAP
vFm69+6QlJDJAeV5r/xqBw7e4AhelRPaUS3cZvX1Jz6VmMB+Ls5NraNNxJbZxX06s3FS4tPZhSrp
S08a3tBX5dt//6h0eCnmyYURrr/tEXVTITsmFXN01+S0KL9+c0fFQ2JdlCYf0kyXU/NE+WCfTbLJ
ioj3wMgjVWAX2GfaqBmFwSJUdrJwRNYy9gYiH2+F5HHS9/7SO9w7bMb4gS0oLPjm1yE0FXhNHopi
hN7Btt7yHgeC+0Dt5DUBPg2EP/BkJSogwGDxPSGDl2F6Qgap61UBGMofh7m78KKPTU0OSLJ60bZ7
L1WgehyoL7UM1LzhQnGRZU7NmZSpqKxMc569G4QfbO6MnEZhsBmz96S0heiJ20DawoBICzdNkRBB
TZzyks99DvtKbWMohwFK8goqKTihe2KHz6BBW108kbDB2+FzCXTCnusTbduZVdc62PqlwULMUhTx
sD43/1nabYlRArV3GgJCKZLsOB02FW+o3m5B+tiS88NAJH9MwKrESHtFb63WQshaz+ODvd3cm2AD
UCWbWxr5z40X5GJxi0rJzaWN96K41S7LGb5gj1W+r+t1iSyAD0t28VlHk4PtTwzsbrTT929BvPKt
GqO91bH7nZEgB+U5V92P33xkTa9fvfzZllBqsY3ILqauEK0YudfcYhCGl6C+d/94p3a5vXixyQ6b
49J41SjXtA6L3mapu7oLK0EpZJ3ZtfRSxIFU3PBdGCOtag8ViNzIBgzPGOxMLPLV7XWMYIWojDA5
0LRSPY6KcBxFwlP2adTyPPbgFZlp1OfOoJh4tsNRYEW6IbA7Y8LsKInAs2RupAqAYOKmCnku7MHA
pQyXFvtSLGyi2Pc08d+KsUE5WpD0lyn/KUC6FrwHnxbC/vWglhtzzEt3ZEsjPyZotM3D7iFeBacy
mg1frDnx/jMTO/jio869nyllEYsRLkxMn+vKboWH7EpbzUfbq48MhNkxd3Iq5vAuQsmlqaoi6Q9A
JZrPjztA+PzbDMMf51QPzMX/7flCT5oSId9ug/qDTiqBUxPX6c19ROfGY97gbe44hJKdZDMjjGtL
LNlobvJv1/Oo6rLJUUCEJDOOyRGeAQl/6CyOepC6mAiMsLm+10+IdeaAOsGTn39xFmEsDN5TqR1I
x6T9dMCVyTPlTuGK+OW2yxXFhJFRL2qslUHJxvx6pWbxoL+MPGpubnGs+lGD2M7A2e15QVAShztF
pj+J5yUIwVTsJgVSmT0eV0ooMyW+X6PK/9Zu/rhP/9AoXoVtug317gzApzQ7Ban5ld1PHezH5wKU
9dnfNMzquUbppdlOdlSYE4vaad+4LrierdEX2VnHmYCWywTCbdfMQpa/3uhIF6UOIDM7Lj75gPmB
lPvzIASpTVnD+82DPndiiu+CFp5gNQm0g3TwUKghDRUoSR0groNTD/EHnYPT2qwri1TYMyueLpiJ
1GUhSCS6WpyCnXteyQRRqsyq7vj1Ouc6+ims/uebr6EplvpPNfrWiNgtrprAWKWKW/A1paIOjj49
mAIteGnQZB+btsQrdAzpiZFSqcgbhETarmz7hFFQbQDtt8jkSY2K2nUxVug+VPmTMKTqCaMM7ebk
ggNtiJ3ltdkfXyFrqTTLdXZj+NYnPn3rfnWIrgYgdy77EyoQH/aIxfpZHrr5koHns9eVuJYSZQrO
Oiws6t1XhFZCQz2pzLuX3Ez+cCEuvS/fUkaRKT8+spfKEW0Hla9uZ406S3NDAmpDwrQ9idJl9ypf
Ts6BlUmqKR2Ml3SxdrtMPew+MYg0BTHMJ7WQJAGa2GwROWON0m0OULSrjGo5khMbj3LxWeOiPydX
GqeLIfJ4eAoXWtQKbPJckbQ3YquBToGzM/+mOEtsOBTF7vyx0ShwmUOPJ4KbMj2x1oRzivQlDL1S
mHsQscPD0gGIrSQr2iIM19evU7uWJbXtOz9qOOfhFrVFtq92R0aq5y3MppJqu1UrTCT2BaZBIj3Y
oWUjr5mT7uIPxj5Vj9uBQGrcxHIY/d9STwjtg+9Bn2YvPMx/OQ2R6LbpcNTyFB+W0D1d2OIjj++3
NNwjb6Ei3oMhuMgWYm8z/F69MsN//ODC4eSGLINYgcyTR8Fum1hzG5+tY9o7iwO9kpqz1WXNKUEX
/GCxDESF36gb3Pr3lYM7avrEc1VRLpjwn1FAEydpLJ+3Dm1/LLGBPC3/NZxkYGyPuCtiRXAQLa6x
rlXMQbXMuNQxCD3bwC+sGCKMGClTz/GjRmZ4pozOCvU+nLBZNwQMAJ0Cm0LM/Pujdq8Iq6yzlz5W
cqwc/RWH8jlCaXKLzg/PZ31SEEcw+cERYQ7/NMlTo9Whi/+n91KGMABcNFcPGuVOH+R+ZkcsLmZb
eBb4MWhNvtxoJzRRTU8QgO5XpoEaVhuncqb6hfg9gsKYRaDeyG6o6y1WETjhaCImelbmYo+Bh5U4
J5HwOieAGfiDmq5Agl3YNbL0zZaun/oYiMnShiPscqFKTODzBMZDg9awBUMyf7BXXX3odHbAVASJ
UMpTLQzkFgsqgjNr+j+XCNKljwRsYwKsNxzL6MW9cxj3wLg6zWmK0msJ8Mqdt1er/A0S6usR3RVt
ku5QHRr9d/Ohgh/TvrBt65UOr7Rx0cU4joPKiCFIDJSzHHUqOaLInhHdv6z4api1Tl+oTYiRtfRX
MvFEDhhGl4KWVGoKMoMAhzHV79gGe9CyFl29EubDK3/x4V6WEErZrPHRMsdLTTcvu3LophhMWwrs
RiwTdyR6AOPiGyfkvzaB3YFXBGTZacrwJegW5oAE9lHPxzjzzo/uU7fosHYk/pHxM5ZF4jJRKSFL
sy9W+uhi51Cz28LMlE2d0uoWS9v80zz5kUPRYrAUuaw8GbctDVAqvsABBk1D3w6Sw77YbtFe5RiW
aqPz9YA1+Sa3wDDNTFHYFqrx2t/YUNJxzTJ1wKoCH2L0WsEI25Qu0BgjQyg7yTVFfcaMQHrotHXk
ADosIp0QSM+UfJjV7g7uXFxfMb8Dt0ks/XGmnqssHK3q1o8Sl30Z0nKwG+iS/mM2m/PDHYVl/Iuk
4Qv9NfqfehfGtw5qh18IQfK1/hoOv570dF+Wbw1UywiEOdj3fjoekf1GnMLJutHWY8imhAlG57W1
DL78yqLIqoBI/Q8Eb3VpKCrXxpTQLigaPhs3u0BzmKs3E/VgvdOM84zWDSEQvnzd9DY/fNzRHHjE
yzBhtCglCyLjDPEWDwAg45/4vwQeD3PCKPs2Zuf6pDmzGtqnUoqDIeYQHXA8FEV0qYa3JgqcTe//
1ZkJ7Brg1bBZ6O4DJ8LbqDmgJCnY49wjho9hhuRL+Dlv89jwD7fsViuB5D1KMu4QReyJISmO5D/c
84glE83kIMI0aFRQKlYLJgxXpoWcU0weZ9cDcV9EJn/wyIwum6J31CpkTVzv3yHjtyFxv/XJQTNb
zmOa/ROXERZz4LxV3jBxEC9U78oGGp52xpK5XsHpCYxfIgI7PlituBZ570NWL59adAhzvDoMS0YY
lhfYGnruf9+zqKeUG9gCmD1v5wh5dJwz7eKPykBQ4dx8STuMhGTR34m3QF321Zed+vLyySdEKfby
tRqrGxiO+WZNkZ068GfNque3UiTA3Y8eSx63gXC0yJQi2nfhsQAk69L1WcMqxmMiATSBvJ9P5+7D
YO8ml7QzwU92+fPyDLvXXm+YegNRQsra6lJAr3XQC11rgcZZZxKQlIbNRTaAGrfzfhJSgK0ijf55
pjsreGtPFGuQlBAclSgV7ZzuLCFaQEIS9wVDO7LH+dPQqmvNOzIPUVTnXUglNW25MojIbi7pMqZy
jiSjXEBtwXokwFo80qRQjZIoUaEBai4svvQiHgG2reXiBZzRNXS9r1p6jJybxr/9cixsEOoYkpbO
gDQaUnclGrEQ92HGKbBQ0KewaMjP/ZmMZXTbRE/DeUlThZ7TQFGCQBDUvZN4CTfufGr1DpN4FWlc
gGqlgjc4oF7E2wIbimwnt+irFvPWctTGH7KPjH0gZbjYjHxCt/849PQ0y2rqvlo04uxEGHtdybIx
pgyMu8STvwRnt1Qq+4sNc1UFKUa/+Ru6MC+Ddc3hB9Q2D7qxK96Q6htu2tPfgx9BX1pkK7i49BUQ
TVCYZ/ZMmJY80Bn3VwvMtvIAu+5fzR4mGa+yDCU6zW5wQuMpAD+61Ipr2q1qEpPzokDTHFBYkJzJ
9zuSmb7fayQwfavbZcCQlF+ovtxhiD2ChYH/qZHBndrgtKgovnGz/dNpu4GaKuPOWdTnVC5jMVAy
5/aOI5fDsJUp3D6H9vSZfM9C6lexakhanbYNN66ca8JmMS4LyAdRRXoQRIJYo2FU3IUH6iI0fCkh
L/agznmcLxsc+CepcUbgIMU4eWIo3zE+lEpq5i4TGgFwAG5vD6aQ1mEyAIul7E25gARP0jukY4rp
hP/AWM5ZgU8nIURkfavLcugaWksqJ88tDf70vmNpJtzqYgsAKYbBda3Faf6mef1obpAlyzlZdgaM
6ogpBvDBkr95ci2OSnjHa1e94zHzDiJJ2c5hJNgvLH/qeUqMrAPVnfgAWFMUGAbgLccR6NYSXDPH
PW/h52m0z/A3Tvj9F5q8GAzxjMXg0wba9N8wcIlklxRDtDjFC6rSVN+egu6csObI8DPlb2vbPbuZ
DoEgqK/K39QzM6VyqbycE4N58a5/ffle7Zn0BqZapsj2GLDDPApe2R9nIoD12Cw3X6AvK8kJVqeQ
kXFN5j8hZ+xTxO4D2VJ1ZvMFj3R6WXxLeewZZhCKKlENWwwn3IIUeYusEsEoCIwgdcSCK7LsDNGP
QQWxf3dK+aDPYFkJXJYamZ2MsgVFa5GDVszRgzaU2C+IbzccuiffEUdtbUOgqrYRemQsO5522BvU
uDs9TbRVVmNTat9jGRsfWhn2/iigQK7SqO939yhIDhV0WiHDSTARozNGz/fVdeO7CE43eA4Y1ywg
OtQ2OAIWd/IrPLKU9UwLYODA10dnWhB7Wz6oG3zTAGk26s5NLuQIBu/Tnaiiq7ZAg6jXU7q+neOs
fXDpGx3N5/KZ+icaLTGQ+abZkzzCXp+lBy9LN7oN1zpZTi3K7Z5o2XMoEW5ZgBA3/f8n4/bbGsHI
yfZeuK76xF/apcCY3eUZNXF1xswGplWV06aor+k3DRU86NyzTFFhOJ+wjWoxkaCKd2h6wND+hKEF
mlJPbiFAKXfNIsRjPNkSgO8cOEWaCpO7PEe0wDtI1XQzG+r6wN5aN5I8cM0lr9dH9J73DHiHUsNg
7l28qd5E8wwEWydmrAPJAqQg7EyL9CX9a8RG4muIGtvjAAfhT3qfehfsjc7LxFGuDsiJtJw43EIl
6J5wv+D1UruV/Td1FD/MKdk5XsuMW0zoa6ySnp25LzSXzXh5/AHmcUekAWffGy7DuNSoh391KB16
JrFs8QoW737BfvZe9xw/q+RNTpGZkhL+sTRSw52bJfLG38brAuRbFg+UkTdehMQ5sWHMIBVddtpn
oeEJvxJLbbjEo/MBUBsN2GsYEVC27flsD22GSCRT8r7A+aedLETDPcxaCyeSMoDTjOH07/AhCdIZ
X3RUfLClAZOBE0Q8Tb1w4Na1giyJB9vCJMOL00hzO0Qyszqoi/k0VpOEFTtpK8XABspS5DINNtb3
8DRYGTRC5ZqR1fVoUE+ugy7FJ0EfjdLhboLzg9Gv0dMZP6V07PbbXEQvtPW6Y+IwG8gs/UOO9klF
Y/fY5XWNR4RC3loRHcMSazb2jUb+VmjGp9Yl/gEbVh+Qg5O98fV1hv1tq6Pny/eJ1mfsWZcHT6fh
zwFPWcgOtQKxyqEkNaiXgGy0Z+lc4M0im4w0EbHWeOHMI2LvQG2rPUcjAJ8gJsX8t13WX6tZGkyB
8J/RCvyR9YbID0U1UHwBOe1z04gDv8hotU0xefD5T5K1FrXb/J1NVXpy3+90hZEfRmoaiV7/LjrH
FBvCMAre0bN7QEOeLW6Rq+/TjGtib8+qoCYDJEuk4VhCP1bsUlzrURb1o6y5S2PZi6EvexKyjk9Z
m9u5E1KOL0DoCYVW9LDcU44dJHsHIiC5QwhNmW3lOwDrvslQdCwY15Fs1TFZsJsNHUJ3dk96E4mH
VKi3xaILutyEFSEg8h7YcjMOSdWp+8ef855mQWo/e5ho6SKaEmL5hKyBECeKEs/U27mIZeBjdNCo
D+o5nn1Ke9XvdExv++tSQKp8ab2PpmzvYM+5OSP1DUV45gKPgCfWd29z3EU0XmBVzJ/CRhje9HKQ
KB4LEUTLdrdlC37joJ+O3jYqQy6xHf0XiBNIFKcP6x3IY/kUgRV5+HmHcPCCFzG5T8WmrzuGp2Ts
ZoaxkFTjmHK6xakqB4SOed4/gtmRGxRrWjQHMojn1NM8xnOyZSckdVyh0HY0OekXNfscZqgsaLAi
4l5Zxxx/ealm20BVVwe+1ETI8PlipeMhO9aCx/HCfiPM2ZPyPEjrpqwrAJdDXhxOWMmif99DwQmr
HTZhuZG36tcn9lFQ5oN22Hj9dc9ojrHkTHs9p6eyX0K/vLXsF2pUFWz8teUfEC1aO9EKD809WDbU
1fSH57EodtXif0yskeMhYROPiLRomAwLd8RgiDDk2SxtlI4QFt3hgqiK+Azrvxil2LwcZYabQ58y
CYHyiAbOpQ/PHjPgDuuZPpcaogmUog23PTyvjxRhPYJBPG5uaCNujW/CaqDg2CJY1WeQ9kPT1xpl
VYBhgS13eoeSDtKUvmQS8GVgFQOCb9OtX/hp0QNODs4NqVdUwLxUPahD2G9088hOk2VJlBbFc9Uf
VYF2NGwGTldGU56jX7Dw/DHBLWl/KnsZ59e5kwLS/4HBN+KQh/wN/I4BD/0mAT/abz9Fb4rI5m2B
Jb7mWxp4zkp0LDIupHRyH32Q8HgrVle1qe5hLXSg25FQf0fEF8UELJFG7Bnl6iams6luY1AQRyO9
VkL9cRey6pZpQadQIYZthqT+ADtCjuytggxV1BRleeNruvW4sCf3sKs8uA/NOV/U7B+QhtjQ5z5Q
wNU6pkth6UJ0P/jtqyRiVpBHcRD98//Wt0eH+fDK8tM8Bo4ZmKADWhbrKXlQXxY72Ud7j5/qAffK
cFb/9M50zosRw8Hd+SzKU1p1TbTet9+CLF6SEGfPVIr8SvMzKsADSKgj+eYlxXOzP41ZlCIawk4B
afeoF4iP7iDRAMjaAkwy/adVMqQRjvJm92kSeDjABix5mWYKrFMPb8Bf5heX5aDmupKOy787vluH
qc3IKoy2yZkmCSs2fEbSIjfSxmiMSldMcx1RZG7eXsUrmEh1MkPoQC6j8o5xydUPL6ko7f2pkX2P
7VjZAlcoRleO8DvjF5E0j9keluTzDr0DypVSn7NWSRvn+ddHigkZMaF9pyLc0l6aPsNmSK8BNpUC
eTmMenAhJmoJ8zSF7+RCb0fzlUWW58febWAkYMAU1MKAwgH7Bj0w4e3UUeVRI2ljimNow+X4MOis
uaL2a4MoN0vkORYfPiqySrw2UFGy3TEHUqZE/v1ur1yD8dy65BdkwhtXtxDlooGJ1LhLrBp6jysc
Gk7nX+m25PAz2ZVZ6IxIct4Ia9Z25lt/9WbKLmXm+uMPdUMOUAxWf7et/NNuddxDbEQOvb3oA/Mi
V6yFyB0xhiRX+1K/uuY1ZtAvohCcvgY/ardLwBbAhlREkcXd00VLahtiq3nFSfTuM6QjhLv1Pusf
vgd1y8s307uey2UBh0eFdRfIkrsB81MB5qVcC0Bn87YKlWAeVWtADEQKZl5M6VTzQGb/SLrNSuEB
4fTlTd7CM4YsLwNPfHUbm2ksvz3mvfnxIE6cW46C512+5Hu8pjs8TXp0GsuKpElNYg0J7WkKIK70
2Dt8RoLR9nb4v8dgNN9OZp2j+S+KpiRI497T1u/xS5Axv94RarhMF8Q/qVpbjqRFAdD4u/EcPvDQ
IVg/RUNYyriD919bdGZNqJo1NfJBKE6eRiaWRk6C3owDLu6bJjQG6RNA8uR0aBaFWE2/uZDRFKLI
IzW9abfPrM6VXeXRQPMZHUV0I5lQDGpr5sevDOOMGQUmVCfr0Z+JNxK/ESCIygTVp4r0Yc/dWjCA
zBamNMTVPimEaPVpCJK6LkCqYaEhgqVRy+hs7/kIZ3Enyj3tuWWsG/4t54whjY5A7AGo7FWgvnLc
Aqg7ytetJFCnx86uw0hDzJSnhE1nZKfsP+VoMhyInNOjNFN+GPriv2RZw/q/VGMqFKOceQZYI2ws
W2CW4HoJEjEhejDwys8VVNEtjR6Ws0bB7pMlLvaOUAh9D6FXbK+F6ZJ0fD+gG7PkxxnS46JHFNhE
yCeS4Hk/HVy1SSDkCsHpGXpy+4dxpg2XyserEWK6YM5wMQCHtKMRVh31d1mxtBbp6xhsR/glbCj+
M4S61lQZm/CkJmLjzB4WJOqqbr2Q16D8MSXL8h5bY+pgrAYZMVPvUbBRUKwhodeMX15y0rSHHCed
jUQX1SO1dVANrKPKR4f4qO0b5oTyGsQVD9meHGAgwHDAJttXgKPXNuWqwDz5RI8P7CDlcgLDrEom
uPmsJ26mnzrAWjnoMTsgVXq9A9T+u71lwDJm5kcWH9dEOo2O8Xche3JGkEkP+JZZNU0YFxbPRtSd
5CcKOqHiBBEP0Bdb1HUAraPC1yqExxOQnE8AvQVmM+TgJWP92jz1NJhBaW75T/x708/llH1eXsj9
Od9MbPL5bQ7sVRBrBgQjFNeGh9al8jNg8otr2PNlr2iB21hbhihENBoAAcy9/gdPgVUf3tX2UA+8
/xWjvrYKfGkPDHOd0IKNW7HP/+i+eAelrQt2T/hEfNb88m9DS1UaDFeg+eWE376ozWlUamMq+OYE
It2OHW492hhbUOlb+rsw5ihbfDJ77Cv+py4zejoewPYEVTQmKltziR7hcwYpJsYCsDpmNMYivi/R
ooYFO0imohEFPK4MMaszdoolen3nqu2NBknjWBTbFSUudgoO9i1n4Ekn0475MrAM6dP+mOCOBZU+
BnMmQvWj2dPYGmuYFJ2v38TeV/VMBJZlvkHdhDFDVI7KbOrG62W2X0bBuMKi0YXtfmnyv6NsCkBs
0oGOjggi+aMc4XILB+oc8MEXHnKQiIAVkTP4XJzn/2h713uX5yw0q9W+1yVyzPFX961II1vMBuOQ
QA5zXW2VRrFOk5suwH3coIHiJ/Y9muGVdNQf/nk3G9TB1uOwEsYm+ICHPmkWrYeip7IbuxeF8CXT
qf89qFL24kd5wsX6PbPK6hPPU5403yWxYvQ+haviNZGLEX2c04kAqgmYOxjTjXpePh4Xw2oZlFbd
pKdHZjkHOJ9tvUJ/154EKtrF+Lc8no7e9GZNT0pJfm5N53cGmoJz44kL9NGuaBRn1d97bT6Y5Nkz
Vnj5VRkXe3axP/tcaLrTmIfAcmMjhlYeQ6faKELp5gCSpyLxUCMKYKx67lNKPsfYaERxGHAMnkAG
KnugIPc6nDqOCnKm9z0QJvWOwppCzJI2+lmimmC+AK79LBAa2KMUHNHCnN8R3yiFjI57r0wyBdk3
TyYXzAPX84zXQfsrAjq2OjmJKzL7/wNt98HMB+QLxbKXr6O+JOSbFRQHVmmqVtgMdp/BSscEnvxV
+jGoJfMKvFGsCEHBh8VISt79Fafm4oEWeKFm7JHqQVSSOkOK+9ykuLEDoxmazKVNNEy1/PpueTVN
6/DlayrjFVymU6zEiq062k8ZsnthG+lGMPHUfcAiERhO7txl7IGI1aoHO08Tm/asz1hf+vsGcgDm
m5JswvI1z0DUojOzachvPkhEnsaarQraBF8B/9rYGfNpb7N6BYmZKYF9HyuCwGtDQEg4NjjEsoU3
2nFhKFOBM3PESihK5s/dzgVgTYWZVIcYiZcsxiAcI6xz13l+bcwVl6nqG8nJFtWEmGD+kdqOv68Z
mJSUKrUYl7C/uUWeRJMyj4loPX1sZ9FdQbhq38eu7KddkPtQaO7TEVoGsSGh1X5g5Lk9+GbYwxpD
iXFhOHXYkXIgHzZ88/V/dfqtVjhgceKMGiDt67yPrM9igUyYy/gMkFbCZfIR5pa8SsYolFPArwgk
8TAMFR6Aca9QUKs7j9oJEue70PJZNf4mWeI9aD2SBeo9xkEm1KxjDKEE+/4Kx5g9LfZeuOBdF1DN
Mb3ggF3bHfDwkKoMmxl7J+7jtYQyfOBOWN5ESLWF06z571zytVJnvJrE4XL0OAjd3VkEN2oeNm+2
mpk54o1+5+FkoQNXlVsuSkB2acIxbWSPzXL5cFRIpm4jrV54JTAO1zN7w0kikce12RtSRT44/1ln
5frJA3nyVAAqD+Vr6mxkW/FUMY8d3/76Wqi9hqgBPgUQB412s4ow07GPpBrsCrKYjkfKiApeWFK/
H/tp5eDKT3DcWld4qAJItY/a2FWHAqDnLr6/cJgunUw1I/MwVvHIGG0BvHVhTdVtSKLitZmUOlSz
rK3GWWO/UtQWvGUNbmScoBOFyi6Cc2aacU9B8uoGfUgqAQl47NXKFy5kIdgWxT4lvQcRdKqtZqBX
5jg9j+FG9wnbzXzMrIMlyebLaf/IurtT16XZX0HthZEc8Z57amtTtgyH7am0kGwM1apQ85yqdiSi
i7T/LM30c+i8+kkQHYgJeZHmIwWCLptR+HcRD5DQp+HKFSYJFqT6GH2Ky0IL7bRltuAL3lyr6czh
YoFFvZ9H8O56iFW5orDM9s1yTXlBXdJueHoHOJCRw17Grd0e4qvtsdluM+OnqjP2/HKWNa7NkbfE
TAEqVFPUaRCWQxAS1Xs4/THshvDezTTqdEQfi4IbOUmY/hozSrD9rCO6JGqTp/L9lNqmnDhCET+F
sEp133f5FsMdRdPtqt90n/6FIgReyvSbqUUeFg1dPsM8TCDTVZEpcFRN4B2uv9f8axrAxrsoFY97
+MsVTfcOGMAp4zJgnCxlHH9meqKfcZ0BaHCklLIYiDF87OkRXRRFFAoYFOkkdNSXs3NEaFj/ZtrN
tku/2I7qQjjl8dZ5XJzFudA4Lh4yFfvItMGR/bF8vM60fdm2EIPXemaSR+mzOgj5ghQy3mT9ch9V
yz++Cal4XOHEc7jeVcI8Xai877tlTFzzJRgj4e7Dzag9nUPEKW+K1r+cGmOSYPBYr5nfr3jGGbtQ
9+/0UvWwmZoQeMEaXcOGH6hoiqzkX69Otxzusx+aKLCPa08X4VvIsNX+aBcpOXz35R7kO/S1hmcv
RhSwosfXP0WkfDGgJEmeapFL6C4TaBk0jDamnKhiLHACIviw84SKNgqWBpxYCaSSBAva0ERX6PpA
OPzVFmKNK/u5PNxZ8V3gzPLXz3tFNCpK7XXFbmojaQYx8edOsXgSJQQSDvlr2ErfuzBK7wy60TQj
4GJiN0z7y+yFfTuPSHqOgqgUQZMjxLGdUcEP01a1Nu27lPsHBBton6IJOgUHFeiLVHgFNfbLUJ09
ZjRwmvWgSHq/MuE+tXxNOHtL4adOWL/JAZS7vaKU2ZTIvF4Oe7sZaLEWuNp9vuHO7fdhLGqI88Qg
zgsGHXP4Pz+TsCMnxveNjC5rXquUsZIrOecvQtiV2Mbx7RlUf5ZRy8z6mrEyTHAbDNzrtg9SEAAs
dojZ/Y5ixNgUxDihRZHfoQrGgb2m1OjTbCOaEvHAVy8hr4FDg7Ffu8oo1sFYWVWfkQVlfHi2o+to
kZu+u02tT+LfZmTPtHfBqXTF9NEN867l2WlruG9YztPKIUSz0ZZFz9W8ABQdmCM1AKvNFwHl8Yvn
ezl2LpT/JYLo4/ibnR+zjrJLR03TPQ0soL7tl5FqdwzKRtDHsYvVBFJgSLTaXNqgijYF25/CUgG4
2cobR9McqjXQrk7p1y0j6JSoA9WdPmvp8/6fyGWyCDyouLP5mzLbSJA6Eq6igoauMwZRYBmvIliu
hahVV+xgF34YWdxYxMm/Zhfk7zNquLWf/DSKHuMnAE31Bxa7ihhNA9Gx7jzGreU9Zdo7i0+tydqr
8dpfhy0ds+gcJspNExlEMx/kd4/fM3bUtVJ/1LRXPU2oEOoDhjA3q8kyepnD4dZ1IPIA3lt7ThAb
RqodDFDVwVaRi1VSS5hz57w0OKxRwKgNEOAgnHG+KTMxFOX4tJlBfqGeXpHfIZW2uONmXYWTjQWb
oLD5BiX0L5Oaaye5vLmM7kFOqAPmUVmk3R9Nc3e2EIm1DZ3WloNijdYV4sNoJu0MPLWAUbWVKoFF
ugP/qbqz55Ba6cm02AH025tYrNBdGF0hbqYVTcI1GROjnwVkhNETMnQTjSVVm7oVDgvN6QZdYNIa
ZTsGmQ79oeOjvgbhIVZveIus1y2PNkQ1930RIJajX1f1Knb5qCEz+cslD30fLzZfSAFRL949vrp9
6dFGLw2g+fIiJ9ljYDj1ty+n6BoKtjcmU6J94KOD/I/ERk3osu1eo7S1ICHi+zzI1r1xSOdg6ihV
YQRG9SCfXK9AqvULAWkwrwp45mTMNJDXmFRKVixKxoWYtckFX3cha5/pL8qf6NnStUQQS8qdlG4j
KjkfTdylvho190XjjGri5xRHHwoQFl3iD3T+fzGrO//tadiE+ft/MyMVQFnGu3nFo+Fv1zobV3y9
a8RVZcOWmmaE0gG6ljO39jeRoturD5Z0icghsKczsPr3Dh2BdFWZpm0W1+Zy8r+4CBBuTSSaQgGu
FAfhqGAkbilpXH5KNGJBJORG8fCD8ABAG7dyi0Byu54oJoHwIhPwpp2okA2LNawuTiOY3s0o23mh
qmMzLJ1FSGVCZXmKf7j+1uglNlbyrjqcPDXitNLeAzOG0Tl8XWXHXMS4pp9zA8Tah8/fkxr+UnF5
a7mCLxKOCL5eZqA7e6OoOzRjw8NmVmceRBvu1CzaZitfbPdCN61M0nOFx75tmUuhMyeawpXkybXB
WUzRuitT9krDSdxIdNhWxr5tcYluHbggUYbRQBxpU6fkLyiGwnCOk+XOnL7SXwxMEfSc9KVfCgVr
XXpDiQTid7FH+AzdoxxsoKhZA536sMimdi/gxW5eruX2RazbC6Ly13yDbmdFlESpK4bsTJjHmNJz
nzwoWnpxb3m2on7PsFPynjAgzWTuzze3cySg9WSSqTw+eMXt6OjjGfwAs6fJl2+RLLBRu0J0sp5b
amMk4hxkkfZ6wvQGzi/qNIWBReupnVkWsRgHhIpgVXV7PjZKLhNyZX3huAhur2caIug+QIlqABoE
8c+CBErF0v/ATWFW/YEeEs5MrW9gDdAyZ2f6WD+X9CrlklW7BddBbhh7P9vRUseK5FfGoJVNTVQ9
gfh2GW8V59TrijoI7pncSwrCBgn84gxEe8CxAjkhcFsRt8Ga1WST6pyswPORXHr/kG4oytMQpQaR
Nv538nH6LRFkOrhuYVGME4CKRHVRyxFJz6xxllLl62nHbZzZjfeuvv2rhxo6GaeX70zok29JTuA6
tT7Cc838KJZWU7tn5F9C02kw7QpVWYkv45h1q+1vbhTtrsndPKWKMiQCQAGbOfsnqw1Kuc8BsLPZ
CpfOb3IByon6cNcn3We8OGMh8kfsNWa6ZQSWQNNYy5N3EVJJI21XzOz6O6KLdLj9/1LxM0j4NexD
LwFozQXxHgzGSuqG4aDk6LvtvHhqm/JTxAgMc872g71+PRKDTUsxJu20qJKlACa7if8clEk2f+v7
jFPHR4zPSrGmjr7gmMPIENfu3AhGWnHhEKNfcq721YvzTql7h5p+YEV2wlXvkv4a0O8uqCG3jgee
AnriUA/u4VeCrOoh3i6PoplXb92nmfqn+SFYHVtBkDJEVqJ1PDGgAyA3ldmAkVlG6JdZ9XK5lZEg
6UVi1CDRupKlnuFCT4ck6NB7Gxa0tmKmXwqIn61CJQSVWygRNgQuXwgas9mDUzPwIqjcn20fB36z
6F1bg75aDhXEYh0Xi5SNs68EUPab1oF7rUmjL8Ls7ocstj+jxMxtry7n2QVwaExRuoIGUTk8lxw+
7FkN3ay2iwTGmlVAyRE5JWRMPwIog8OLn2NnWjDrJkquK4/koEghua4816xyN4l14nezcUxguAoy
g2dIMl6jfLn3PwPAeTzhY18KkIJC0QA9bzOWY3Q0QPAADwkuiJpARf0anfoL/snkuXOWla1u++e5
YtbLSWzSIQMv90zatpowfMm63bHny4foj2TF7QYjYjTnMoxWKRWLxhvhZ/k+OM4Yrb/sYWzVdsI0
f+7nsTrtUA+Wp0Qtbt2ypkc0HkjfknV3vRY18TUSo8kIGw5v0Tmit9XF7I6MUmiCTD8U6sKdBJCL
kDIeuviBv/QeU3VCM90RYnOrWin2vUi/lyTQK2AVNFm2JxLfszzd3fi7R7Ag8OHcMw64EfyhS1mh
9DNH8hES4Wmbf+bjxfQ/Zg9xDx5DySGJoJutWwyAclVN7Gz0dLUCD2yZj4qCLCPC8LUiYRM+8MNN
FnD+E5eLWyk6g+GkI+xivMij4YBTDQGOHkmr+GiUzaZ5uDaH3nPlBdzJFSoBFJb4V6hn1lPkumbG
KgBbgc2yP14JThpcCNL7+cVXDcmJewUES9cUpclUBcgJqdFOzUpqfBo8SIkic/Q/JqlGQoI/Sad0
n0zqLTV43gQrWd0Cy9sEkkAO4HzvvoRXWjI5My6f+VJKw5diB/kLdv//QBa9RUEjBgmVSvGhRJUb
eEscWmX2V/xAbgLfQJOQebtvzp8GJaE5FtPnmDC0gUH/90qDCUS79vKzMXXEnlbQqjTMPQ3tnRje
YLJEviUbVzfb1ujsk1oVM5+IlEsufq54LWcOsybSZJnFUfaOfPVfXEd/Gb2UvII+DrpfeEFdyh/F
Mz+SBE8J6FcFckjWVQZw4f1WylVXUoVvutvJBZ6S7SS2fTdCW6l5p/yRktejtZpzQiuDaLd6BmEN
RtgbWyA3q4Ls77jefcny/d3dzMGKNA9/GzCBRYjclz6cL3SWoGQNsVdQCHhlZblnk6+KeSr40gxQ
kc9UlSSr/IsV/I6AyAcEVK8FSHxaX5LChs9E6jYXZP1DiCwp2BlsZ14EyffI2i1xqT9EPJUERy7S
Ko/DOZiqoNXtE2NGkzoTUWumVL/tYiYL4ESQm5Qe83FbN/IGWeI0WXmhWgQX8q385O+8Wu/4OxC0
894/oBvqEXyZO8c1ZvFYlz++gOnX41UkE8GebO53vwGDAV3uDW5JKiQYcxGAtayuOCe0Ty5SO2J/
bNG+G/5LsgtE0mkmzva0B93VwUNCbfpO05+Q35i/mqBSm//KRbazTUmeNaZUs1PIArBNpM5S1F8Z
ejQ3q+ZqK5AOE/4iaLBl+sCSjoxK4x8ZxVGGU/+t2te+5JfRQcSZK2xXj4I5RAZmPIdyVMR3hQhx
jRR4QHGuuCYlYJKktT3fKl2YcNXzNl0G1GGtte26z+X11HdD9rV25GDH/Tb6dd/jZ0j32yxGHF7J
r3cdMexVhg/bRumhcTz0WJPkNYQYSZbmGojMRc4aDODof+36LMn0K3QSPvZH0t1+IIzY8yGpq6Nj
W68mTvwUvWf4GhSco+dP1bwcJAZI+irwmw0dW0tZTPe8+6xGNTkRafRcXuVE6BH/MCPMar51t7Dt
Xa5HOiWcMI+l8ycP0kQ3aVp4RexU2M09WGhHlz+zddgixJ7rEzFEX7r+bnmwCm9fo5QrodEVlSf+
wrnFEeSkSsuJOCe5LvfTniI4l8JwgUf2boiAgVqD+KTp6sJJVhI343Kd8lJq6NUP2OSwRkoGxHU4
BG/JU17oCNtTU48/wBXQo0gSkKotxX9anTOJfF+bXl/bKiWd4ouvYHvDDVmosXrtLzbzFVOG6ewl
15WbH9PYbvvJXOB5aTrIwNjxraKnhsDUzXWvHbVT/8QEZS8PeTXwGGOmm2eUpU4zMthEtdFAL0YQ
UZabfGUL73CY8fWXBCNYRMLtaZNbjnKEZ0my20ZrAZZgyTT2pnfJeiw3VlBSjsflGggHnRR3t3fr
Kczax6DFMbp/82I84wyg3VrL9TsUCxcQZU6QowwoKestBt5sErVSd/ZoxPjGuTeZSaBqNfYd5yh4
7Yhe1quvYZ+rolPHx60kA8bx5yfjEk1TTi13wRNAeW0ndHDdOh76lisFqzkCj6fWgXotTZ0ZW9q7
e4WpKN2KecV6qmVDtSHXOkJY3SrRxLfe6ukemJpH5VQAQWqw3jH1vvZjFaj8hI6W7wyvLuHkoG7S
Uc8lkGjAwAR6RXRKQ/+86qhQfEl596xQbEBS62wRpr4tHV4eJgcFPG20CLKRx4NVyqg5DhXaLHY9
jFopYGw8jU/AZOdgVIEe33q+dNXnVREA2pXyoDcCIWtgy2g5OjWkM06cLys1neFVBdgyOXRgGz75
F7lvIT0bIdfyXkKps5p97+V6+vBP4zJ9cTkKPVGHxkMQ7CEvQD6jVSScDfF+yjDBIbZxKku9wJyU
IYVDd1Pzh/pNrVcLiTMhPMWmq76SjPCEekLjnHHuPcDW50x+P0RroCzj6xPPIKniC0gXn/8S7AYc
Eu1JfPB35DC6bsFuqVYks8Y4mbFGd/hm8k1UpQgEDzNYWeuFvTg97MTtB5OmKJTGjGpvsun5mGk+
m2OPvAMvo7B8nlmKIyxaK/JiCEj/ZC4J07P7res3fN/jkxyHcrUC4LTCWFPN1X3O85ulhstdOTCz
jDnEDmKRjezcP6MVb6rnpZ+EyGSDZ94RPNTkCpB0fqIY+Nr8SmF2KeYxeT8YMyhc1hG5A47PhIQK
MYxUan/ahihIDhMN7Tdn7zsbQ0HcGoqgWzobg5wGSXUesN9VFuFpwwvKBKieH4L5kI1r7QuyRzQy
VNSw63/5MOKityQV9/rvtFwyqS9wl0t0i6bMNw2zFKsUikhomtjsA85lttkOEwC8pOnWNck5FHV6
1sPPcM+yh2ZKF7GU7o8vpTDXZDlllh8eQpQVI2566ZrONoEwzrd3ueV7V570jzF17UCq122rCB5N
eaM1wpACfTRCbJU1jtdYj69t/skmRWkbY5utsRw/C2cNOluT+CyUU8yeJtFyqTR5tSeMszJtE+9Z
nrtUrpfla8NAcsoAMMUZGJske/ggBJ37barvvPau7tCcejvp7GhjaoUofc97hdyw6Jn7iBmT69oI
J7/xrpXtjYynKT01JEzjECX7uTCBRdlwW8ZGd8bnqjDT0by/u4OmxnJzYyTYsCJCsjcfe5Ud+ykH
5Sv6rKI/yQt7jEhEdxPBQ+pzpJ7KNTIfovZYuGji6qmtegRLP3Twsl/8zP7IkkfUGzGiAWZ19FtF
+ePfVXvf4l7WEU9hYm+SRZKTxj5dLWbBGFcOd4ASxrMdWPEGUFpwrHSHq23mliWMLDnoxu9y2WAn
1klDyL4qqKRG3kSpzKbgUqsATsV/LOzdLzpT3zec0R8wOlWxXxg2KHKEU2v+WnQjFYzMMfNP1F+A
4peWHl+zT/1yZ3/RFAfdiQDUERPaySJaIVXmCmGeFBHL+55qwp3U4lfFUSdG7VrJ8lTwuUrC2KCG
9WkAVPR6SHMq8FMyemrHNmyT8QoQJrFaepk9qLp8d+1Pgq5YaZUJy32o+New40OZciFegfsqhMc+
bblcYlF7cGqEmRnPdQGDQfqmL0DxN/SoG2aL4q2Lof6Ze7tIvfnfKPT0Cn4b+BJIDfzfdZ0LqTXt
GM+AS/vRk2LNdJ4nm6hZnPRJuj7GSQ1J3SEjV34jyH/aOdBjAOgecw2CGnk9WbGt4YSwr5kgGT2S
LZCmSVv+wwzwdbkndHx7L5CkAcd9hDaotrwRmSqJ1mgDuzo7HD+HxBbuyMOO6ausYTB9e2OFDgui
vjYMh8SBfpG97FEVjozZ559+e2/NgM/IKF9lOBJWCQapYnH8f1zx9G62RQzA2Perig1KtIUYoRjN
bt1Nt6SRgrECKUVM8YGLbTBkNONT/b+e+bz1KM5IUI/szcweEIkd5p7kqYHpJMll1or2yh585S1f
hC/Ex7MAWcm/5r8joebLsvCSwhV0Du2+WZV28uOz6+d/853cHAuttJziGTnIcnqYCw8/XWOR+rPx
6Cr9ttfza6/E2gG9NRi6V7LCZGxoYCedcowv9nfp/AL6DzInvArgJtXGbc+RuCnDFMaKjGmyK9v4
U8LbzmVX4VCWhz72c3L4CJi97ARxUtCKPw4ukxJ5I7aceWkqf1P85sN5fxOglHkyTRn/sO3jPR/L
3Q3v5vpYCvPc4qLIaEkM1zF0DMP3cZ1+g1hw/SsabMBLwHoTX0DhpCbRUDTzh/P58nbpEGydcoyU
aw15XKEHqXd8ZMhRcEoy6YTuR+QWRQt0m2vbBCYBxK+P0jJMHuriJOKG4A026IWKuOi9cimDTDD3
sNlS737rBrj9zRuMbrRJOiZEhM5fP2MY077MElkwbrgZ/kX/5fAIDktItcNmcERiiw8M6KJNJBDW
TFhDozhu+c//ZK5Xnkd+K0FOA+8PFKZt03uQ748YG47I2dO+Hi4LEkjpaMmvmm1q1QFWS88XCJWV
A+YAnFYtiqOqdvcN/W4+dMKi5YvMQ0T1JnzxYkZk7P8HAZE1HNjs1h18yZdrby7YWeZfEKJwOBSY
d8GdbWT/cRJB3GNIECKAOMCD8+geP0EDbWZWHC5o/l0MTd+GLGiQ0jR9t31cLiXgiAXvisdRNGJJ
snEPWm2AyY3pf2XaBvvILUDI/uysLPnA/FbQP9Ns6emn4rPB9CDKeSXxB+xKivFkgqE1IgQ975U7
Pv/PxFnp/z6wIf8gOH0tiZBuXdvXv36z0zMqHyVB65JZWaiyWWy8geYIOYp9juJ7n8317As3VOG8
zR4qLQ6SbpVIvY+5mBbrf/eY9uVN8n5gMYWzbL2+Ok4CUrLE8L3Qc5IzbAClfQUlx7uuVUMnx+S7
GE6cAlHv3nYIWFGWD+znoHCU60n92Ii9JNzbOglTGhvZpZEdbrCWvgC1bufPpZblcF+jMDkIzsaP
cL0rFTxBw4gbl3AsBQc1OQoIFXrFvAReH8bZWQOlQ6xv1Q2DnV4CCZfsKqSXppjEIc4c4BILgZkI
EGKQkExApJC9JlJqYxlqiB1REOdvSMOypxfZFPGYicrkbY53fzn2BJTs13jk+D0hic8fvU86LCA2
olPZIzl0Bq4zBP7S9umsfNOu5Gv0v6JquBKUlZsFoeb3kiN3k1oBywMS8rSInTxdIfo9mnh3aTux
FluqTPoXPXLVIU64jlNz3+raAEwk6hKEzxnDJitFTjWtDUZXGTC4pe5/DS/6kAVqf4iRmrZvcOCV
uSAKsa7n76ffKrSrFmfuYLbEbxaHenaqw7jE04d3p1jeEQNWmgrTzylFbtkXlkfQDwxWBtYTYbq0
4j3BjLsmuAJcNSO3MI4Th2EwdgmR/CkVFT0sJMMujBurg74Wl3BHn+aYoHzrroxLVP9/xWQ2n8w7
+l4lcrLtxOHQ1FBxfUM5YKGVPrI8g8iafieyIUhyJNZHB1L245GNK7zu/WRXcls2w8WWxN/73aoR
gyYAvRMBOaIPUvU7gaVI4X/ntfh5EgzzY7qxjC2PQnhZaH6k07in3JuSIB8TBLx9j05tVe9NWVnC
+G4iGABAGQSYcBaT0xF/JRB/BBxpEhys4C0/0xRz3CaePOl9nP4PzTNl3Y1dy3SuuATWN99wVB3S
ZBKbIbd1jOkNaxjSD0Oe0+2fEhIy+lBUQgH8HFWJWI7YVEQBWpMllrMxEap2GqzSHLl0uQTOho6u
6QlYenjoC/09AVvHJNkVlMOt/0fE0NLIJFVk9BsI5FDH5IIbq/jt1YgPZM7Qzbz5iKA/YqGIvksH
u8zBl+g0hnthqfLxPkudWhgqc3NuPCFsdkC4gviBKDNWr+7TFuJA5NUHHbiw6i+fvrayaNzXAlfb
Z4DZdc8+QXkfENU5Y/XRx+AWGYb9O1eVwyuQan6FdbDY794M6XmdBLD2S2KVg2pBeh6wURNHn6SD
ol7UHC4mGhR5hodQ3YB4JeJ28JGIaYvB8lXcBiefKMW7M207kmNNR3MSdpDoMMRwpISOM5jxc3BU
J6R417T12XMkY/yQ9zFeHrXvG2Ix9DTdiK3RtdhfQUizAKqYwHe1bPylvAPMrBd26/er+vOrBiO5
GYPhFlI8IozpU0PZzhveGSqy0PO+dxNGQ+wRSVElVR9iQolD7rk4yHF7EKcckpbP24XCgjgUSM+Z
+NMVkYGKGPbwg+WgobnfimaAGkYbkng5vj7ET5MezdW76JEQ/Lypeg1Rei3dlZv7Cj5jWl85CsDI
kMwLx9DMOMcLUW3MbT6nJQsqVDO1igyE3vKa3y35neVkTHnXMDwupRetEvtZbXCaPDj4B4lQyrrR
Cdo1+Q21mpjCvq+10Sms11ojEQyas9fCqJv2Cu1x5sqlVtMD2SHoDuEPiGch0rWe4svgPa1sRdM9
qVzk6BzGAUb80gw2ZlB2DRLtSJlj0tql9ONcAY6r6cyKPmi7NcIk+f7M0R/Y7B3L3dhLpv7TU7fn
ERWC6VfeYp/XKO+aUZxUKrxZoxsT9K9oJ7m2TnC/lWtvF1rmJcmq595yTAtn2Amq6FrYNHF8S5pN
izqiEtmo1ZEnSlQ1K4ZuVMGYjnAMpXAweGsuXZjLCXn5u1gQYFgBStHXwXDzvQzMpdPQ4wAXGa7v
t28rPNwBvpERSfG7K8WdOFwNL2g1Zv+ZdgDnfUvir4uo2kzDpm6Ja1swx711K+E6O3nmqxoreLV2
nq5LOWqY9kVRJAq5TbolXJEmgnoJyKrxvWTRlRuHoGx1zemcrNDje+xtXQL48tpLYO3g5ORMSh3O
E47tTjgml2vElmwZkeCBafQ7pnaBPNPOXv2D0610uEL5YsRIqwBIEPX2sGYozRXgOyCMFVNxckqy
SBV5voR5871IVDCpI1i3klYEuYSA76C0OgjcUBUbRYnJfFUBVIfhRnTSqfXZc2mpQaUQjIdJKo5N
chuxHyRSa8w5ClwHx98V6YZ/lgcfsrmfsfM+tPVwOAA86/Br6eF2Y1PWlAVQUR03CoeN7ibJi9g4
iKCpFA1jcmOPDCtJto+JyCuQ0DoHdW1JaP3JhSQUe9cpLAwNzS5W9EKabsqA72/Ri3wimD97hfHL
CAvjcpwEizu6wUvFIv8ael1TN4m6fJcP8+p5LvKVkMHnBpxm3i9VIZFr/SirtNAoYxVkiheIraHd
4f+OhAtViYUfAwNvr/EQIiXmc1ZYMocYWkebr67vOYGOAqQr24IoK1fztDl8faiDAKST1xoPrwyh
WaFNtB5egLKg89mxepV239CdKhhROnUWOG7tfEZFWEqZFEpsrufQ/eeZYVYYuffHv5d8knlsgDiW
iOKK+Gs25JFfVdTyqEciMx7gDG+ATLocqY8NUWeaBawdqtg+mSFJ8SY7oCNaRaGyGJiB/H90ccE0
3YjDZh53ac0FHsdZTuZG0qKLdecJDHg7MiXlUlnpZK2X4zOE69xIyiiY/WRjZ6TZFPfw1DbDGEJO
zf5bS+0KBuV2XdCp9LZ0iEGnNfsKwxf6WecogmqMf8kKizvzqF7MpzgQ+ajIz/RD+uE2wb4InQEg
BUbOaZSHjHXoJMYxwmNkzeYa4NMdqkWJ1/SFD2PKb8YhLELl4LOqM5lvCJXOCJRdXTVurFTMEYsy
PvbHb29xcwQyBKd5OBlM17LazluE/UMWCfMZ7hsqUq18bXjfriB6k42f/0fPq99jNp64QiF042AZ
13TxFOTAAbyv/QTnQ4IL4y9+og3Rf4xqgkc4k9BfI0Y7/5SBgrl6Nz19L1yjctmRuZSovUOmZMaR
mpbmRNnjwmttfQdJrRFIN6HANXPu9/LwjzQHjRubUmNJTn0vOJwxhvKY8bxRt5e5jzyWEiglw5fB
MNX+nPdqXeOXjcw01UHXOoGer91eec//X/z/LYhBrzcz0ljPa3sxQv4bq1eYysf/JjJkjsLfL4VK
Onv8g+t1cLKzGZXPd7qyKcms+e7su+O1ekqGuNPFhrlFOhVDeN0YqLJTEnk+feWsvdNhp7yHtHF8
XsPmjuFGIGfGDsvw3Y5+5/C2RzY9zmolY5s01YzlqU2ZElh7hXb7EH5+UqJupXiJIHJBL0hgK5KR
7nkY3TbsRERbN5PmQnodAV5+zt+vCuqxo/qac5NywOlW2z/ndV1uqC/jxMxyzs1gWRVbHiAAMOUZ
Q9xy0zovOP2yYNpatck58kvnqQEJH2LurFdnEtguyhc9Mx1AlVHP5RsNL0IAPw6VK2ge9fK1p0Lf
fKTsIx1Jzva0mbCNZlnETjOWwrk4aNt3xW9lq3bcTEvReH+yWtmQ8LzTJG1xgZbNQ91hE2t55XnE
xJHz5EI9PEh4wKU0R9cxcfqzF4P/ckiRg19zEZD4v2LKzLWeog55W9vya2U2ww564hB0ybyRbZ29
J5oNsYDBhMAJgtNVfBtyL4/2NW4POgeChbWwJ9X9gc66NYM0eY58QfzMn5MHXUJ3LSHfTZf/Go1w
1ayJA3SyD/Qpvvgo6d4Ypjog7LAaKVCemaGz/q3x392zX+aj2B6yFVwo/VipZGvopeEbYpElt0FL
7l5WvFxVi4SzVb1cPqWGNyzzkdWTm9hVLMmRPCSi29NXe9NYszY34S166fDVBftcvybuj/EK5cdg
ZAY29i0haKMUUi1hwdhVRw2vD1egAIJyB9CTSWLSOQQRQRVe1uhVxVP8JkZSoT4hfJt0ksX6hYG+
3DsOayLk8981zZEPfy/cau9eLt4vgkuBe9/EiJkF/YIdZ9lwYMN8mvr5JRB/6lBxQ+i9V4vrxaHT
ia6b1Xs/I/G0lGyeEnNKnAT+cN8+SkeCEuXbZN35wLf97BfiCDV+X2wdVebmwvDhkGtxDOWzR3lq
Jh0jU8ZxnHFDofJZVRos+Ur512sw7RU7zQHASYm55K+IpKxnilrtE7Ua+5Jh178dH7yeIyYs4G3z
GZfCypN68TWMrELhdjxAtY5kO1EhPAZoqMqPaAqrvBhohYTUGXtuYi9z+xtKU/TeqrNUocpXMKY6
gqh4rvdm/a3zlQTV2qoZJGyUxcj5XTAq6FafeemCggCk8gU6L8hy5vydwO0Tt4vsUdPlMBJzlyB4
alozT956TPpSZdVzRXSj59BiUb5Om5l+Pa0wckEJuDdkB0MMrqw6EI64tNiOvvDYNSCdj7BzAnJN
zdOK9Lz/TWLyjggYHhkT2OVNcMCJ8LkNSxM7RV4Ov+oPOflBg1KDKZF//arKHK7AawigTnt4bHP1
1DfGRLcbgtR/Io8jtfQHOyNvBv0gJcm4LPR9/3pr8gIpqhaf1ESBSjNprYHRTo5mMKjXbc5YZ9ul
XuJ9aTp18IZe7iZq6SMUHzHa4sS9sY+/p3wpYrDTgFkONAZSBoxzA2tkecTzTGZTW3GJU6y7DZEq
X3SF0MjNe5CbriFK/fRE51nRW+kGV8jMpwVQQKsMjMP/fkkPCHB54cLQhi+J62Z5sssDOzkGGOAu
zSrldEX5t2nWYGTaeBGjHU/XnewREXN+1dAyAkBfr7Aj7FnB5aG6XvA11coUclwOvJX8HkdGDN9t
It31EUnS18KOKnz+EVYSeYDj6t6AMEdpYMrL+jRy57Vg02Rt+ko3YPfe1jjmAPfaO9PCWPVurizq
pxDT35UPA5m+ADXpueV+5H+v22vmqEv479cwgE7ZDS6cB02FD+22vyaCBg/17Q+gcsYPbDrJCLhz
NO4VmTM1r1BLZ0xLAsjE2Mr/43qmdhv2gA9XVjAExTMjf3Njeat6xnQ/R21GVQEBe7QjUPVSL9Lz
r8wv4kktanp9uOOljpLgAP+RwqYWqKrmMeK5K3sbUQSAvedWBpS5ShUJJC5fr6U8Gop/hqb/M0/x
RYDpJ06a54BQ6Z1KfT5F1ib3mxulKZ5wLRHvdXMTOpO1uYbq0ZaHJguVtSiZiE4xenmZlVKKFE1e
C+HSW/shLEg6RH9LGvnDPMhWulOZFbMUo4YPbwZl7S4KbkiCktLC3qDj7VfWW50b0TSgvm4weLte
+hSUFZ6we37SOhGn6BpaIrfFQ4WN1iO9h1SiAf0491AYHIOSdYdWjqL4xpaIH1B10sgaKPi4rzek
kohMCPSrejYQtBV5D9RZhEM+e69XOQtviFOh9LVlxK4lCFukkJ6b+tlVYuWrv/Q5wSyfWHAWaaIG
maLHAvej3AZqAESOdLmt409KpR1Av4DNz3HGgfzUoCd2qKoQ0vh0hI6ztqJJIyClz4i84l5ha4UW
PTSf1mHcUmQ8/tb1x+T5GshCH0bDmREDX5lPfqzs879DBuhrrKsWnwIcjeF7AtJkANEIN78/KVdT
5F4CqP16SMbDEv7JiNZpeEIyoTDSzmm6gEAik3vLmxzbYa72m7zhEZcSYK1YzP/NUaa5/jAA6w+O
dsVnbYNRbqSH0y8l91XgGNfyUOMSuu56B0IKH00YVi20s1gDETK+Fs60qXDcBvUKVg6u819J0utV
+l7zPJLWthgGNPWimtIQbQRxhkrdwd/DahNbdW2xkmyF5E4tGGfE9raEW4yLcDjbt8SXlXdq89bp
kx9m0/7AyfgU4gf5p6FUwixztJhLH23YKX1IuB1WoAA4soWUMQgfSi+9OvaS2yZo51KvzSotpet5
/9r4S32XqwtO4kT5R/JRX/Hdh0hwt+fmoQfZR4VWt26I8Ksd3s0O9JIB4p7Jc8GYruNzwetUzNDZ
mrPZlILxZtMrs71RyZlB0/6RdN333XdOcF1/0EgPEj4VVKBPzZsvWv58yOzbbLB4mtYLazEb6mqq
L9Dz0fKL12UfH+m4FhOz5U+xSl+X03UyciQoSmklRX2JjPTJBCDVUeSQGInGH/ZbYMO2YLXZw8wA
4A1YZiXN6rj9P8M75cu7eOb3Jid42voE2xoM9VG+pHWQ0bce0pqCbr8GiiIHsxqGV9MKFokA0kKN
rXKDFbYQP6ThwKXlG/AH5A+bTIduFYXxbRFMmpR9cciSqSGZsWN5o3iycOwH7P3K3OtDSRI8jw/C
863j8Px3lfgtXCdpRaYbl45iAVmifV7GUYYf/HVVdZ146PbvSoosda31R8Nk0Nvapxf1qd1N8q2e
CKjK1tjJZfsVGD9ps/di6gBsyNMRhPJwVEqGyE00iWv9qKRUhQo2xt/1292Z3UTXfHbpoU+M72mT
AuUMLm0V8ExULztqhz0Ip5zlXOAGLrSanqUghjVEtsurI3P9psBtpy6mf7MweNs4gFSHwowCiX9a
md+2cRM+jY/1n86PstAC9jnvbFZt5v2WhgG86HR2zhgbiRIalPD0fv1dVDSWNGu/RKmtkqKnoOFd
60TH20zKGpTotBNhi8qo3BmvT/BEVDSrL1l+fr6MHgonLPAypXkCADrEd8Z7XOwz32ChD2aVSd8j
ldnKzJnmuvbUw+YIgdqyufZlTHSFQ9x2uwmVwVi8DlVrLMEngDdCyU1rHH2TmdP/i2uZ353m+L+r
pAJe6j4JhMGSnk39PMJaG3Ealfs1wSSvi/5byo5oUKd5OeAcuH0LNrSJ5xkJiB+VvPRRT90iU3l2
4WP/lQfeApIBW07MeCOPcOZzs2kyjJ40L8YOW1a8w/f2AiXt1Rx/JzSFZ2dXY4UG4XWQKAhBkjGZ
33KbPUKoEkXB5LvJvPg/zf5mFXYjjfTs7S3p6kaC7yE7hK665kN5PNEjO+dOmDvlAZ66eY525pNl
IhzcpvQFVK3077YIq7xCNNoQWgQ4FDEQfQnS3h1xYF5m7VfDuOIzbhdCiOM1MuZNCHvO6Ap0xx55
QLNP5tYGgewtbbAe75FDlCgL6TiOBMpx1kGq+HwVblWLn08ru1SB5clrPT0JQbU5n5gyyP4Fuy+s
2YvHUOH5twqBG4630IB+IT9Arx1b6HsvN7IEweCKbwPyPbvBiaHj83IaJa1ADo2QGyyZQwBm+BkF
L4PPVpeV+K5CHFchxW9Mxrlyv8KCy/pDILHMZJ6vWccLlRFuGumQaHEms/OEZv65wNv1DUMjiyvp
HCAr68iOMF1DGWxaZ3DFRn+xFrRqvnFB/9wBiyGc9v6TQU2Gv5QPa6Y7sEPAbdg6teH95yk2xKtX
LmenFTzcHLhbglxfbHtrmHOy0wSgNB90nXInT1afExwprOtTnzA7HzmPen4AY7ZPkLbh6CR3pTMD
av4zCdLO+wNiIceTpQO4pJrXotMZws3Jb9D3XaGn5XWrsTi902OxXTRVAfetaXgXivziyz4iBd00
EVaD4nJByCeTKRW2evQHpO1Ef9xand15XSG9YDk6MPPQpY+mqASfvSJ9Qb8R/LxAuwJroX6L5Msx
c+64PHI+j6EmTq3RNuQWmC1lcLJi0g8565+Xx2i7IJnmcFhwLZgC3b4zwX3SnrbSCAy13bT2kd1E
CccOnBKblJDrEKTMkpwdwtZIzdUXf/sKWP6xUkARcV09ioruKPVBWvwfI/Bq6SIaY9ZD414gPEwQ
u3VD5p2OTW2qU46wryIk7POv0pj9QVLIGbv1Y7tgJO8n/aT8kWQZPUooiXVPH6aXeiPS/uC3P2xK
qR1HfIVcQWLc9RFY2NxSlm/chNRVxX+DlndS9h5rpOIaoX7Z/4QGsUpPGwO3+pCkISQJLuYBwi40
HP4ii5gY7Qmhd26B93nPbza2vJhRR583LF8bHFh2zukgpHVvEaWN4jaq8mFNAEKJWdx+QSK7UBkG
AlFJDmfRrZ1DCzYMF5jssdthmfeINDyIx1D+qr9j7CJovndboeFOwiyH3qwYHdA+P++4UcGenq2g
4O0z5Y9F221HF8wKjv/ATs9XoQ3W4B8lxCDGqRZqTC6seHN1MFFAZWvhiK2cKPz4wKCQjgtVz2JF
9iir/IoEvw93ZkV8vKj4dXItnil2jEBpCG4iipJgJuKS1Sb1pf7t2C5ivdDrF6MmQeqn0QZouO2v
qyXqn+LRZ1eXA4s37scDVA+0KIGSoQvbJE27wLdNXz9I0PkeUFRSUjDRb1kIBKyAEFQVicW9MN95
6Fdah+hXDET4RwrotAPwh7tYSGWw0TCl2+7B0fUInqi0Eo9owDgn1yLRpjDSj+vh/NaEQo/GjL9q
NFVbbW1vCuXoG+zf4c/IMoxzzeLkfghmxGdztqhLJfX9SBCpSTpdZCKP/0iuocRs07FJzPwGdfJG
99XbbCr0ZcDfvLQzvVGVy53MRkGjkE9CV5/eIlFMmNMqaDXmfacJ9VoPw9Wg6ofh8D/yevRYZxKt
Rte2Q+zbHEv6w5FNpbCcfavHo+bBpqhlbPByNw8WFPF6y09VK+NrfGNcOZDleRynYAu3Cb6Hl28h
AxJk0G9yzdvR4VGSfiJYSobDxVB3810Jg4Ekn477phfYGsKZHQT4Wvo49HWISmrGBuPBYxwRGkgt
/6hjGzKGH1huJamTLJ7+KaDD/p8pcg8YgU0pq1txCbtijzO1NUfCFPH/Qy//gZqEZpEvdYUyZu8W
XYSQCO6cyDkoHatjYZaozBz3BfNTzjLLYHs8GlZ0gI6MG+kdLwvUNKBeR5m9jpG5khrniqrlQGAn
bFpBCh+W10BTmU/VrEaAXJJafYAyEQFI+Rawv3xm0u94EQgq1gRylZVi9Uxiy9Qb/PaV6lawssBL
ygZvw8WxfQVNKPdGi6gfDTxDx4fzl2qHGQtQQs7i+mjvLBe5Tk8ebqSE9TrjsxY99ari0wyftm2M
CDnaXdDmqEictp7OdLvyVweTeWwk9mLSJf2tUsdyTIkeZvlRcUcP2sc/IZFtvpWZZp+sHAQac1Ol
vNpLgzRCCu9Pu4f0a9ABPV1PzQ2yaT5hf10qR/V5obKZWrzlh/423xLo3vdIynWw7cxx4xSMMtjj
AF3J9QjJz/35Lv/JJdfqDQro5RGVbIyxfBPwEGCVd98PU3yWIiKvPFmfuEmtgvsRsXhCBSZQVSML
86xTnPpAy1zg3heSpD3z5ZNrkVoux2WvTxd8O2OlNRAzwxw9i/iNxAbQ5bj/oqZqTvm8yDJLhB3Z
OoGbtb31iYj2xKwpZrIIX7kTy43dRdeypbXIqeYuAMOLikztCRl2Hjx9eMq3XFNtmKdsiI9PhzzM
2uKT8uF/+KKKZ/Kg7dRcWnFXq1M4Wt+vzgUAuX/DCg7/n8otwZ0/RqfAhS34+txS/RxO52ux43mk
Mep9dy6UnGs9IcZstVo1FMO7lsnxGzo2Eq02vRVqqiMJ86JHb78TPW0DaIxve/Bd9OROsOLenXky
+8OuIdr+hr2+uRuitlAfarU4e5/CDnCMJnKCqgCto+Xz77p74q+xn3E7sm1ea7sPPInNxkXijQDK
X9tMbFLjQq1vIAwLoGjWIFs9LHRIhNcdrnXlY2I9gobVXPsVxGrZgTWTADUlQG0MYLb3VR8hffRc
Zc/+JAeaMp6wqwsUsMvAjtm4uKT7lDYeHFf0ffUdIvHMM7jmjjdQNRl2hf/W8WqzxDucGLA0LgwZ
HyKf8cqFkdVKh7sNmxiCKDDbHCtw3IQNH8/KNboFZX4WrUrHrQ8RS5TYsAf3JH7vNNiVHgYwII41
Q6qAeoEuEDPLW3zO/Jn6t+vMQrdwPQnc5qgQqrKyOWVUKfJx8TUOA00BCx+1c+J2a//TXQQYqbVs
1XeS5F/6nWJFRj0SLy4Zeo5/8/Lzt6Lz4gmVvYd95EFcPeFiq9K42GYpaRJNF1R64FtzNh7QFBYd
xuIQkQayYMiOpxTQmxoN38nQ/C3ktQOAy5EnkZEg/Kr4LpNbLkT9Fp+sz9TMGzVwJIUwtE77T2Ou
+1jqfQF7+VVK3k0wDO65ofeycyxWtxF/hPAvnPmNC88qBPsbA3ZYMPaHO5VRR6j45/7uFvz+kfxr
uJPJalLIC7pvqL0UosygfCzoRkhTfhs6CtmV6+9IBjQ2p9m0OSDufQF/qZsmdtyqDh1ZyTA3XIn0
9hxYBoV+tSPrx2SBXsIqbhM6XdDN9GFgpjFAaw9cwQWuvSIgPFH898FaGWhSj/Mj+JlIzXB84v2s
jSzsnWpXyF3Y09ruvAd0J6CncunH0388YXrjJJJ+F+XmjPVnlFdAVJ+63B7UYcdRwZVchypCR0B8
rytDGAhP6khzmf1PYkpuVkfuhMQCHV3OT2AwWAyfmWpCh8HDbZq9UAtkpz2y7s/rx76N4swytOTI
HldsJ5CLR4ib7nK3iSUh6STTHVcDktVZiWo68NXwvW77JQl5W33YSguLiz3fMBd5is93wX16vNWS
/+luT/wgouYPP7oVTEDMzk2eQ1bMbBfpAOCSZ2+0/8kS+WPaqbb5N821WJIQEI62ZZcn5p2HD2bk
AAOG3JR88DJfJGdCyQ9x675Uf/yD+ZL2C445o8ZeFVUzPkFO9sWI2wP5+FQYHOR39kT2llReUXv6
tRBKS6mfI9WkgRWsSFgSn3NWbYtoUfxl/xgEwXI8MHlbMRVXNXti0Angy8LxfrhUpm6VtWgZ3q1F
imYlPcL7koizCTFzEIiSJyNwMBqh/RoRgMqOs5eHUmoVE19PGXPM7Z1lzM2aspZu4QIb2VjWDzoo
rKlN2dE4jdGoxAvAhjDkkn84egQatVA5TFfjDaHD/UXKvGABEPPlUD/jPWuQP975RdICY+4jyAj/
KkbjFYFemQuP3cCHRT4DO+Kg8kRPkasNWoTQltkxtcNigRyxNd11ty6Z60t44+X/xrTHPtsS2AoO
s7IBkfdqcvnsM1lV3c05d4Wyw+lCHMc19gTCnyFAISEihYFLEVk4QUvFnDvXE1KMA1MBjFojkLQ4
tV6K+s8RFYp19yczdOnIIrgC6sfDPA86wjJUQeHBOSY7ruUiB1e2bunOV70E+FSkKoB0vrZ8kGiG
MO7tKkDfpi5CmZg+Qr15yG83XTgjPBDQit+fJgLyPQB7DL4AmlaY4hBzkVDOgV8ZPCw9nuyHRhP9
xbPztcfQzxjN3QuK3h2DMJBcECInpZrzMjgfgkb35BDoJchBeUikI8YdsfcDPOf7zSbqCUhgvraK
kLjFGq6YTSkDE+iJMI3I/WdPzw6NnWkZs0u7YkaaUVa1OdALX3g8KR0/6MELZbbGL/XDczSVultl
ybRHQ28YNSR6pFtQ7owfPsHv2H4qrS4WdATwvwJheeNUmS7nG8oisr/5A1LiBF+rBgu981OWrNCc
uq8tVt1N/fc7lQBOoyXxsC5Lx5fHIKnAUwk4ghktJCOE0Adig1OThq8YmABgsJ2SdR7dO9lo9rUz
+rzBBIUKIzEsOlTkNQuU1uVBhhiQtjH3xWO2IA9+RZalNB9kpCEt/17YleK+WkIM2CYQn6JsunFH
c36KZHJ61voplYrThVMx1gagp127r5vTdjZPKJo378QzXBWL9wFY/w3xFGZ6Wt4Kqf18TqFbgZhp
o85zfkcHF49srpOuyZiMvYl6WfxVx9Kjj2YzqSUVW4ksr5TshbM4q9qeFuOuAFTrSWjMtxv/qxps
aebWW7s2YFcjJG4R7ksI5mvVmTiwETju2/ZRUQKudX7Jmo6KHcSwHC6FVpQfTZrvLDStvpjtSUa0
jEeJ9A8M4LkFFwV2pg9mR+e8VgKk0WfDHJFn6NBVhzedg6fShSRIfjEHXluoIdy+Jo8QqMcoy0AD
1Kt+zBD/owdPByeVlye7T04COHrr76sea7bgT8AQzQFoT+tl2LRuWijmkNRJ3CVZAsxKblNLdeoh
79c4h1vpCts00XMV1WKXto6lnZl0OeeR9zNiVw5/EmE5leyDuYn5vg6H2nwjKAyYbhofRBdXW3sU
IqM0c8Vw9yt7yyoeMIw7sz2zc8H53J1DC1U/0MpEFqH8GMOjBHO0TiFsf3GI0tVy/NodX0pohrRQ
qQuKDQzW3gRBM6CmksC1xrawO7AB6bi14R8ZoG3CBLc9lxdziGRyV0n/ZXB0gXB7f8tYIZWctyT4
PpNHQx2I2AvEfJd8iEOvh1OtdcsBVq8c009jtgEH9bjYJqczwTrtJXDNxg/oY2gMEOLo9vWa2Rdu
e9yzUhz0we99MsSecjmGl7jkki8pNzD8lkbSBrDFj2vs+cJiHZXkf9jT9NNGN1TJ52oLuv6xCrXG
QC3WG5wuOgWZNtf94+o1N9YiTahbvEjKzvgPs1eSiqWHMcBT3IEYeF3fr8sMvqdWLfch1nr7Pk4t
Zu/bi5ISnEP6FAhJoO+CXhPIzyy05jiXCFWlmPuHOcnVI84COVW6DGoVk8DGhzUxywxgGCfzb+Yg
M8E/sXPQn44LUi5zfaNZyijmqTcSRMKkrJHQg3/LpkEF3B+IGepbAMW9ZGPOlCCUlfrIMJnTIxuF
d4oh641V0zvZ6kACY0hL/irY6ZNN9Ol8S03nImRF8nfAlnSFqoSR3Wxuma8WpsiKplofjPb/8ccP
PrmJfiahJDmKWPXmq6INz4jJN8rrc8m4iyJvs7+6RiMai9wSxTDFuQqvkedZejeHseJOuD/Bo5av
S/TDJk1AEF0b3WrQ/V9uY42GG+ua0FxgCyuUyi7g5oy4Kg20jDH1cmVU6dTCVTgFSVOrtiZMoGk8
EOWDN5ADrTDn9B2r6zO5OrwW7tL1siFAuSeLpRTO6qu4NTa49lcqwYs6GeorvcE/9GOEVZQ5ckUm
gMBqcaMFvMlRHtzdnkMfleo2zr/OWaNl6NKhO669hQz0xn+p83voNVVMOmWZq9dBg4PI8mCuo6BI
dnUdxsJ8kJJpIbUm8rfqe9JksONcSrVWrnQRTZ5oRS27kIOLTvvsCa+LNPKoNRHviU2zX96bQYUU
qK/W76PvRMYs4Coo17vPAaeWmVW6mPucN7XcOyr0y51U6QiNFJzpup8YeV0tEH3GB5co0DE1qhAe
q3Lk6ZyMQU9aLaDLpZQA5B4Yu6aJVtAVE8IY/3xLuBTwVTakAtHvRFkHBR6zjzYRPQbHpiROgr2o
FbL5/8MF5qw2hKY0XNgP1/zTy+ljGqOBEtdHLR0HE4XgNpkLmlDmK7uqbEUtIScZq/2c3cc3bS8H
PAIzYuGretNlZ6131p2gqkgkyrkKpk6V8yVYWr6o3c+Ztw4EQMGmiigdsDQaReMXmgTyo0VPZle4
IMenYo73gMo4mfdDJWmR5nCOF1e7NAu0hvW0Qa0+9WjyVl3Z/nc8Q8lN7CEY9YJQG2zoQkpf79fy
qQFt/LBBKt5eWEA6BNKnTyJV1p6G2AYeNmV+nUyOiGtqy2S75QWeEgXAInIEx+5CjewE//zGN5hi
88kIgwJitMkpkCh+IQJKrZtNLMidw+5reKFirbjBNWbxrqum5S8vMcJ+kEzjNvNqUnciHbp3mzZn
vDNNBXeSSGi928E33+asvWi40Vpti5i+bqnZN0vkS0y0Ublj1tJDV0Xs/mXtc9uVtQLQcguRB6La
mae6RM8018YUjyMHz2S4UpGDgX9Zmofoe9cKcW527gFAJLEAV1Adl7Gj6kzA4CZA0m/a0FLb8No5
/O5+To0Sp8Wnw1+5Iqv6Nx6KvslhelCVffCbp91m0xY1ro0g/E8CapEGU1oDZr+kj2LNkN6LFIQz
8AWE18nER6wuN+neNoQSGVvpI1Qg3yl1++1do/RqKrgL3196Z4eWdhpCkuXzGblHWb3hqPiM1FRy
a6ji3kngC9fdMAm6TPrnWO9nvYWR+HSyh59UTcZrT4gnbHrM/g1d4wYxWtS5SNR45BWY0Nz9Qubj
C1ojA/es8uey5hIFakyHQl/C512S77B09Dibn6DibTcUz6asXtoEjm3O9Tc9juzA1SAWQq9fPkc8
LBwvnGlV4CDBYjp2Bg6X7WcsGsrm3iPYX5tqjKUJCQaIHjvETp241nWu6F0puBhrRL2j8N0DZ+q6
8yCsq6bN74Pz1WOOag2bglYprM4NUbrzkTVFzX8ZPXPJwbqnUuHAPIPZCSR/KmSGoDle8ACtQAsQ
2fnPIF+SjhxUdAdb/SQ0WhojkTusn93zW6TtGja+hcWC8DB/Go3VvDRii52gK8Z3ErvwVRhERQ1v
ZzBSIfr8tp8uryjwniDKVAn24/+R07uuRlHqokWqzotOO4qf6RuKxB5ogrZzdL//7gNZPsXENm7c
L6aMciXU8g9wm/O8jjtgfIkLaul8ynX2g4xqvsB1ytg45MvRzwztrJQeQVb6lJygjeKRyHDAb3Ji
BJpedkwCDODPYNJKIxI8H3SSZBmFH5NgIvFAD1pso1c2UlB3Hi8vM1RksxTDUxJxoi7Yvi4z/h2D
nv3DtNR7Zawq/Vs8WAkHTuHMOLzW7piYu1KGTaUS94dcFVtSRNEZpjPDGS0YAXuCT4qY4DZdLzfq
Sun0APVrkYUvc9ScSMVWXAbpUbY3JIUU2QFwbOO62tKdqXoFTlspvlT2Z1J8emzH9A2wGGQiXd0g
UPp6EYhruyaYg4MyBRXjnzuUe8VI1VrcvuQ3l++a1ZJ+B+hzWtn2cJcpAi7K6Vi7HMfH9M/YZp/4
6n2t7iXQC+dMW9KyvrQI1mHN0HcMOD1HF4foyxsTmf8KyInQ+YMb4pNQuzKuu3jtT7WEfnudWgWv
ghFOChPubTENUHO8D9nXndLfeNHghehJI1/gZ31P1huPy0u1OLT156dYo03YCm9HvmbtNoPvOZrr
0R8rTRU4KGmguREj5wWNII8qCRB4ddBeODORYpReuL46V9gCuF6ykF1kFd0QsezSj9MJ/T+sq7UK
aRNKikoo+FKfXlT8KCcgvvdHv4glJAnTkhysshbge1nS86Qqt0wScaHWnnvOxELBPCNGygQxueRo
UDRIB239Gduwy3PrKGe7Q74IrYfr5HWawCEt3l9LVDhZi0v7JL6fVM3RvDOfmSuuEMoiymhKf8Ge
DkyGyMdELqvBi/HJ+DdBk3wi1K+lMLi0BqxmujSmAkv2OUSclUbfB0ryuEpj75DiI9DXhsUc7WQS
aCc2JUw4YUmuRn4q02BMP7dlqQfTnr5X0W64XQmLVwlLlh03up3OFCGsgNT0qRiN3oBSt8sp8DSE
CqOSHRoZVHTDyc3sZiiY6/0+G1e5XHbo0FKaD4P3IYRNsfA2EIgbKb40MlGal43IqAkWXm4ms4Fu
Us5DJrGyf0WBD0HrMfMWfl15rl0VF2opXs/4Jba2f0GKaOGokloqmwsVgFbIvNCH90OTaxFloU8J
g+YPuigTsvD0q205xzvRGF3x0IUEy3Am9GXGkytNtcqHfgVn48YqJdE2CIMVtR+arGKrpHh2BH9U
VxrUR7lNsrliJ6UA4hdjEuKRJXtP/1YZnNNA5H8DYiX5vL9FCdkiVj2UJMhwp3/E9gHZ5hWvLBxP
ez8vZdiaHjKUnLdXfjLy+iuLXPPwUL1Gow2t5BO+vp43IFZH9dlAkB0G0Oeq9QvrAPlJrVSZvH8h
ykNIM1LffiqHDBZsPezUyNKRoeoxPwNk4QKHs6OLn/z6J2jhYMQHlA0pcEKvr56+nIR+YUj8N2Jy
TVRED7QCHdnQ0Chw6qUOg1lzJGcAl7IH1mCxLESIznEKU6HoecJram9lsa6NbsduZ12hB4fVstYt
elZCQhMjow2ZcoTSKrJmmUxGJJOhQjg3GxdHAddkvFD6549xm2dl3gT6aalJc0ayiFMjd0WT6NFq
lpEdW7X6sj/ZqnAJjzJMuTsp5Bjag6cdXG5FMwPHHDd+C1wYBbNCWyB2CdA4ojCdh2xRaFHc4+6i
eEKypi1VlXrY/WQ2qofiavL9MVvbqJZK1QVwn8JqPoTGLarSW+9EKFKm9omKIJW1p1JKApRZhZWT
aj8puHhC2uNaggad7+AYUaF6y/rkefnQ7fPf92vARRqEdXvhpfT8/VUTdDOlkf9hdqu+YUbVZv+z
0vRyRtmRhAjnPapK58lqayJYk2rRaImgTeimEzdwGqvfNHKDJ7oX6ach4lXKMY51e+x6OkaC/ue0
+bful9dk9Ta/6nzqheu6QzRw+nB4o/yMVB5es5J355JpG9yvsrXffTOhZO2YKRdw2bPMFJPSDakx
pNauvNDNA3RegFxnylOoZB88kKhAKueLZEinRzpKVMc4u0PwEeioy1uS9QplP/pVxUocOGW6w6M/
3o1Cq7NrBIbKLph9Do+fHF+GI7KkL1ykUDtIkpDOt+xOJ7zclC3OCjHjGOa5ECKNAUIDHs2KObUQ
Y3g2GQMC29Irdp9ps4NjXfkfQQ9pWC23Fu1+lAs6PUZVfOcJEpzcTP0Rm1EvcPnVmwchZxEyvQ2N
fvXBztHiBuyIktqOW52nu9marFXpY6c1VR+A9sMV4AeBrpHywg/Acrc8qBnLz+wAYNESWs894Tzm
8S4slkd2Y+3/ryivqwn9HJodBRA8ASo7NdL1fk+JcFzAgocl4FzZFoBmgEExlFmlBQsR4cF851aX
9AQPIRrL+qFEZ5Y9srKIicp+pzce8M+TS3fF5QOO9bWlaoK0scucWWbS0aK2X7gYdtTiFIQyhEQz
KfPOjWgfsKok4GOeByzxbAVsYbcq6K8LDIG4HIGH1+iP8vjJjP94o4ZXbnzSvBqPbv29ZS1PCF1M
YWlsxM1/Hn2sP2EoeQPiSE8WycpXvOR9XN7CS1jyQFxAl6wFzH0wdm6T5MVUOj/gp7y9plmWdS9O
942y8BiIADu8puhglbyqLhDDBafpPjUb5FzOtlA2QuuY/ab8VGhzjiKDRXvYa+LA911tQrq3JEUL
4BeNzpBnTz1XU6hjyuPIqJBCuYTzKtAt/axLkoPFg8zIzoXkxtfdZjPw8adcpCWZhgjJDsjAP1Jq
6ulpcGKZkIiXDiG1kYivVUv5ZUW/TpcXr/xL1kqwmt1drohwZtfw5d75I2nVBmTKP74YlG4AZflZ
o6RINa/G6fUo2kGuXR7CNF2uiqPIZ7pSDXw6JhiZ8Kbr3vIlze9G1CEW28wgsUPZ2KnRFWWAu9vN
Oj//z6mKoucCNACkn4dIl+9fAD1zJurOQj4eqqT+PF5tSiSDdd/fmrNVc+P04FSE/y0c2E+i5x7S
hmKTaHGB6oh3+zr8Xo9fJ3cTJoysh00t2C7t0IvuVkGHFQx9gveFIYm8RLdW8ObwatkUrXhJyu/m
DLbcqsqGSUIu6d5h9uYdYjkTeJerQKfbplx8yxKm4vlkSFhYASlX/ZGT8b87fQxj+sPgPED7NDZm
R0RqyigTW+4f+3kKTE4H9DHlJDkGUWajL2q9CJgRtBJsPelMgOcH5TZsWH/XaHARhEDEkNLmu/Xp
JZ6rKPXxUMq/NpwjY0NwBdR5TWreyPcL2Lx1K9P1iO75KAh9ew9dNGIx69H05H7tlEMsM0zY5q9s
ya9uCLeWAB44ficGe4cbIQKrUea7stzl+xE8i3ldfn29CLqiPzgGpz+KiQ6b9/a4XCouK133T+rZ
htN9/93GeH4ElgTUfBdjcJSyk7i7tGlTPZyOdJVTHFVQJzBZJI8JEpD5eFOBagrzz6yK0Ske95d6
1rqUq20X8rpV0WhsVNZN90iR+QxLzj35/lPNElckjt4c2k3KIbdj6DnDcppS8CTS+PjzqPXSAH/o
UmLKgHntsIQiQWD8QgxUU9v7zKC2EXMfvYSIqH+BgUAOO7ka7UFzmUiY3nsKplTQc5sgnDVBxTIC
PiwK+GbZQFRoaBPfH0Ltumfk6aaS2Kq0V1crdrkTpCcvDBeTKdsyT6KyIME+vSefy09v1P684PGo
zR8ZLwnAgcfCsGdvN05MpRLKDwKLBka2jQ95H9dvmEje1uAOG+TOEvH1JAOaYp6RwzsIfGihTrPQ
+EBuzcS3+pRboGeNLBpZIekhxfp/zIznc6EUsFbRbyQk/DLHtqD8QGwvF+KW8T69LSaxfDwD9zPN
zvDcJB0s/Sik0zIKzTTaP65t6FB8wAd3zmAG1/zCZJMu5A3yOByffZzW1JmcGZltQp6GKfbkFfiD
k1UJZQoeyMV0znSVwDZFX58J5Z3EytFwgvfvE1jx29lHReXQG5prtSOov5T3qVJ51DPvCitqrjTj
qBUkvPeG8lb35Q0ppViLUL04Sd8a/vv1Z90+aje1NqGKD2zcuKOhG7NGrAIH60TUw95n+IO8WL6C
0Hm6pmXyi9pQt2Ys2v6DgvCtYfkh1TgHVvlMF0f18XVwa3sabRhcAsIoLbHn3ib3NOUZPsftDH0L
9SbbUj0YNDsmiXwDfxFbD9xM2oY/NoFWQwVSEYlpG+XLD6NRlh4NRJyj2ST1LKa8vbr8HOK7DjZM
009sWXm6WtvYsYRs0CQvFnAfvDx6C/aWN3VGtZTP8+hl37ZtdbDdzRedMCtp29I68c4EYtSg+1jX
R6B5njs5punEK+TYe73WgBDHnYMQiQg+hkyd4fJhv8qoBcdnpir+vXA2f78hTfJS8v+jih/iLLxL
Wbps73saW2eenGgrr+2qGKk4wrAfQixXVrvaV9cpe5n6KywxgLAkqm/t7t3fjfhL5NHAE0szwrQt
8zsv3h6zytaqmQGLnD3reOVeakrBQWJsshrbBf7lL9u95qAW8+n2GSniHm1m+VH9I2BoaUqLJkSg
FDKj3ZFjVMV7mq5SgOnDKfF+AdZ0x5DFU1LATY8xEAqtXSfRVUvV/SBRUZumKaBR0RnGXutFTz+H
TQly/VUzSgJOUIqvfZvuHWE6+ntnxwgGsYu13ED1+0RsDu8QZeLY6la3A6k72WA270mS1uclS5gv
+l75zKEU54RIGioiOwlQM7NPTbwUOuwKsAp4bI1MIj3Qbz//k/ZetyD7kkdO6aksq+ZvpTGTTyEi
AQTkDtgGedi3fjRFLDR4JukR967z/k43RQW0fSK6n5XRDSSBaVB9F9aN1bcg1g9NsTJitvVnNsFc
DzAollLi5vdj/3UsanqGju/sN08yev/Gwqi21ZtkvLY6Y/9HS0VmZWLcxOISmhNZ0DLhx86FRV6q
uEFY66+QUBMM8v58zfG7An7SUFOlR+UXpHxi9Sy83amlqyGtF1dtVzSq0WJYF0hr62hRpjoBdSmo
shTOZFMbfUDBvXGqS38LhjiEd21g4kVB/ANb0iQL9dRlpZXVfp2M/DxX585aSZIptu/VuEZHMiJw
PxXUnefWHhMPBvNkRYSo3twHMIdxSc9v7ISkz+x8Ax8Mdg9jfNtyqR4RhYm6M7VVOWsff08Me8+W
QwamdO5DqWfv6c0B2N8ToZDQFh7snIxlgdh/60XvgSsduY/rbGsMpX0cFA7qSCLHGrR0yjFUFw8F
DXk0If3N7H7Ec1o3+73MHHSIy5tDNxNUfN0evCbuOh5nnJhrHm9dKSAfk4WyPlo8gaqR1gvLJ8h2
MrfpuzPtqIp4wuInzl2mBUoB++FAfKb4Y76aFcmICQyMxnPhwX7Gyzz1t8MnXhr/1JmfkWaOfWJV
oLwRxgcIWVh+jtq7+8CA/RQzj0O5V69k7FDsDRhxnichFLTxieMK13ceB6wS4moci+k9QdQHeZHo
YwHtdacIPVXZ77HGjdanPdc7qX2TGJbUvHOR32ZChvVPJ3sIgdOVOI3UeJpUb65Qqav2NToKSKm3
UuR+hK1GgYV3pO82j2zicGxqbAd2BNoRMsMuKiawzVCmIvoOIcyGJnoUuuLmB+E3KYTR3X7xgxRM
xsAxveUDhNuGYRPxqFsOhr1embeg4fjiCB54b5P9Gf1nHNlvmyyO/z5QtZaBRHxIdcRhF/nEfwTl
Q4Xzr9IOwi3IQa9kSmHRLp1pCJk9hYHJytogn4aut/78M3lCvycYoZh+4dUvf80hcLsEhz590mOO
tOX9QD2JzpjQ9iC5L0cEZftUJgx0eNfK77c99WDKxjm5EV96Y2OJuL0jeIHDS2BELSKR2PFJ9uHO
LVgcI6yGsZwDkKV6GFxwdKnK+D2b9hrFqcdHmoPVwlELW/VtrWPXY+qe0D6DBOa1tl3MdK2VbQwQ
EyuKshYDqh3Du4OHqEx9k58l7nDoeqJl0w8t3S7RvNsOQ9UYkgWe+ygTp2xzkJ/S4hy/HrmW7nRk
570kiIeMKkECAVdBTovfIrTTK+s1eqiAttokucJeGfNx5c0rj0EEtereRfkjA3DRGZptMJPYThBp
6sdjl6/K3fc6Bta5pa9ULNW/xCStKB5TbQKzRGhhv1+dF0vcd/qXkzwWcjY4V455dfNBQK2CC1JB
MIacpjBpE9xbpHgLNx4Reog1SF402zCQn54HBK+plJHyx1UoM7zo5SUrfTmV9C2qqu1ZOXK6seXt
aEDFa2Ng7Xmw0p3Va73yz6AZnzg1sYIUNz1utvc6FCOEtqoUzxmjQf0eyM8nOfpwjVBGurpfh9zE
8xQdpQmvQPBL2g6YKzVEAwpsDHD6QxnM1PA5L17k4bHYGx1LCJwt6mIb4N75D1Ei+sK6xx8mY5KZ
DWd3nn/CZJT3LhGSa8G+y0LHDwGB6BPs2myvembZG0CChtVa32DxVbdIo6rTOKeQoNNczoOy2bLQ
2b58bMC0OHF+i3t0/47OfSpZF8F4/N+FMzA42fJkpa1Zkg27NvmsJKgtckfElTAe9AIlF/6zeUE2
6rHwFmoOFXduHqh7ov12TLttr+2E4o7+GqbGdKEhm+hpqBkuaVh2uAvF6fjZ05MCkY4G98avgtjp
s/SYamEqgyeTGDlBXc1a2fDANV3j9tgKB5L4qm5UjYpXV786HRvvX5x5f30Bgm26ABazqEj/yo9H
g7SXn03Fg7IGjBrYFeFexXciE/ytGMd4qpu2e3wqeKY+p4fkAZri5fXtDHncSTRk1/w25t8D1/tl
sScIXsOtIk/KODc8kfyR3CNKBjxgajJPc1wwYzBjbSSw7CPzamQzH8/8V7HWWUfg0U63kU0Ao34Q
C7ArvSZ1/sxj0ZP5qs9wuOu0kvFVrjs1yL/m/Giw0f9PM3rluq++Egm641YzkuRS9YAPhrpqsssS
LN+mcP3RczZcgJvjs9FvhN6FOq4UAVVZl5LMbyA+6jaE7Cs78hzgEfEdRMnApAAQbnt4Rs43dzal
Ku+OU3OHdAdelqZ+dK/yyPRkfYQiB6ScBIMB3Wf0pNKwRGAvI6O9steagOwOEum81+/DFUdvmCEM
u4zbYy0dfMMDRNv/mG63feojFvEh+Q0g/60ZLU5p2Ijb0ODsQHzxdqESzwpcn7R+Rhb6WOB0b4kl
Siu/txZ8LOVRSNSCCXDgJEllmqqLFV0i2a2hnltfDnYk2bmr1c6xSPbQ+cIX8qoUoU649D3PqQeJ
fWDEZa6Fg4IxqIdvV5SDpfatbTJcHL2ZoHfqYnIVmlrPVrbiUyhDsOy18AOss8zNrxtXxPDqF5Kd
C7rzNDW2uVjuO8qs5rOyU4wJjr2r/vPpVsewL6fGrFgn3nwaO/J9uxuQYAjsPn66QdLp1h/p7LHv
QOlc2h+2gz7l4Pgawojga0+Wm16DHNPf4/9Oe+N1YcjCRf4fd9igWZqJHAfCeKjujNf1VD1SCf+g
xEZkJz7yEmAhNuPQgwDLukumZYwj1lK2s3gciCj6LscPp8FnSNVywwpaBMAEeSHlwxpLxlQg5Wg0
qBvpHvnVmdanMy8rGmiQ7NVWZ9l+ccTPD6HGTPvx8wzEj8+FdHWIBk5WhZ0H+xg/jEQbQXpAU80r
49bZwRdlGRqXefA3mvt2HX/kmiNx1Mh/9phlS+NlKIb7DkG5bCARKwhOij9iTj7EaremoxNX+VKU
ZrJrKbLQM4rV9bR1C801hPoU4NVqsaabm6KVAbNxcrZgvv15uOSt3Z7UGGThQa8u5RjONKXT/0d7
kOjH6vNLHbVScmKmGK9WtP2UISgIBs9+pPXLuKMI0Jjm9UlJIgI+vD8OqRXOEsnjA3XfsS76ZQi7
o9k9MBjBMm7Zo6ikga/jQjPYM6pmnZNG7xxoXAMAZJ++cNvvHBWfYQRZqQABRCA5Xm0rwBqKAtLp
/NznV/miaDXm3pf/FL8g3ggpLlmNg4r80xxWf0r/+gJR5C0mPLbLcx/coAmPgiiAhdVmVAgon2LH
zsRiv8ixZoic4c5mgdDdDGZ2X2hIlw4t9sZRsVj3g9EvLUm2ixxKvYe5Gbr6SToMRM7FwTdIX+sU
KtT4+6bioBng7+ZE/yVx8wLlVvSdnZnMMlhb4zJhznyMdvnM/bqxBvRqXBxBckC5NuTwxZenQPIz
w19cq9Mzqh3Z+Jk2DoRS8FbIxKuWXb+AEUwHwF24nL7GVO1FMyvdmeN7bFfwdI4nMm0r0bMl9maC
06M71vZBlS86XG58hnJe4q3wVoGJ0xlBW1WUgDzV/nuC3jfzjtCUkhMObgCwLBBs4hbpVAmpwshE
HAMAWxHGcElh2adKuBCMR9ncrV3mIiT2RF9A4t6s0LVtPlnOYE0lGQzk/b4AfiW8ksWAD+ShNARU
nxVYqLN2ZKCNQTlLPuXaxqct2L28dGVsOLCpDB4/s/CSrs6wLSsVnVdCcuvnI83JYscLV02Qg2ch
Sr57ndUdzrNb2BDg/bWAo8ZTTYxCKGzKhxaFYC/SFsFfoOxVJfY+x8NrfLnAVe//uEhFfyp1ORAG
CCnsNQ1bJFMYasRVxn8whru6xkJGB3HdfVM/YKA//HaztkjP50yoRRnYKOivlf+/4I82h6TVmpDY
xPYV/YDxeBEv7cscgHEg0EbQWqn0tsCxV5/iTUfvPl3kcR3+507M2MvxTbVyzDlJcKcvObiN2qvL
Nmt449xmnkIYy2ZeLYRSIWWSl5YTdnODDUeooi90kbNZYzI4Z7N8d2A00MWHGHgLLYWZ+j8hesGr
6nddueEgGBQY2x1tj44cMN9dvi6sc2IUfaxbc5MoOqd0P9eawKkm3TBkr3gFowed+6g+o2qxSh0R
vRx+87jCFmw3sRtjsGX8S/J0UAgG4zYiYSgDwbJb1j9kXk6psf4O2Vos9NI+rouVY/qSggqTr/qO
x0GiLRCAT6QCe/B+yPuNlxBkUEzyXlUDE6OFZyi4PxDp00zDmKOTp16hXfwed5esqjlccu1Cw9Fk
M6/c3bOXZgd2z9yHWBE9nN75KtPj6sR51ujrx28ul8F2V1oplTWaW0rcw6T9eWlxukSV5yfY2ZET
0RjAw1eM1tlnJrO5+nWPomUhDfSQNpEXrdBDolzPncgvHAvox5m78T7PfZoHv7AvDAtokUjzqqH2
Kuog7smbg+HMwdYTQeJECiFppf03rc8qKtvFBSPe3F1Q3oxBxEcuwa3Cd4jQgxRe5vHsbCC+2IGk
YY+hk7zc6oJ5Ad9knqEqTaQlssjPqrwFa8bMBDefMK5NAP3t6eZzBQCTcJF0X2Qj6l75+Hc5XqpH
E5v+mWStR8o/dVVey/XWJCHaC+YgvMiSK9esN5aB2pWIX74/MD3A+mHBoh9kGdlFFO3LA3mZ2X7e
1cIN51ZfGNwK5YgnlPVBcLQyEmTxHk+CsIlsITpTXd0VTvN2BKLYHyetX83BD1YlmizH89Ucr1Qb
yNqPhlDN7MQE2MZ4D53dAmVxnr8AjDATuBfSlqdb4nvT/ssq1pHfhCfTX1m8Nu2Y/nrB3YQyitsi
XDGhtbuUrTqfl8jkcU4rCbEJkVP6lCcIh27QcM1Pef3nnh04d5MErvjjCl5t6LE6NJQywtGHHl5I
XUSTqa/SOHCkRBlIXpL3sprSyu7vlJX7bxWaLDA9OqCMyF5BqyyQKJGkIyNNz5EddHpd1t9OluoG
eqE/T0Jc1AdlA3Jyvyp59szK6OYTOhNWJ2rqiA7rDPajzgJlN9qxODaSmoMnoggNfWfU1X0jBPtK
H44oAJis8z1qcrRGaw7/zWFirKQjLqHyfoyNAD3emaFk8j3pbFfIEUpBGFvDAQq/ujrVIoeE66VG
bn2xlm2EZkgJA6C0v6eywuUIUbnu3xpfc4BVXN16EEzvIjqzq+NYhBzBLKJu3Z7rH6Fz4qXsVJ7p
Q+Hy3Dq9B1JmRoeVoGAFZsBO+7zcV2vYLS+vQjTQXZbfH0cDV/Gbh1TR18w3+Bk/GkOcjmptai+p
IIFBGR4GZRJ8G+QAdYnNokhEzuGVhmV1XkHgC6++XUt8HfIBqGEINcACLttJSckWgXvLHpEVJKwc
oymrzl/tokTn6t8S2zv/JYXG8L+fhmUX4g5HxGpm+MTJQyH8tLPEefk3BNdliU4FnfVvho1bfNs0
ybv0NjANX+4JjMOJhOOH/z/21hP5jqDZN7/vgElndwiVbiBk8W+Z0pLXfgklVTdO8ThyShy6ya4u
ZynlbiCUEPChKDXEBPto3W0AXkzbMHuyZ1asuhouDKFHc4bY4d2QzY8r529CcVYLcYiFs8q/XKp5
j3fiU0XNZCcG7o1OsBVPnf+icyLSaPdUbtRxlz6yvIbV/LY8LTg0CExkUrZMbM1awKw0hRHVUDwV
Vwr8/FDsqKMupHRLq/HtBIT5j/ZPWcxMthUKnL/fpzVrrB0gpa8hvg030eCSaOWecA6SSNVKLQOc
txdmc+Q1ojfW5QPubFXu0la/kb6Krj6ZbV+tsVyey2dWge+BlVecxiTl4mZunuPTDC7nklnMNGNg
D7jrPkD7HmG3l11bp+VpK4/6guNLUeg0KgTeEjVlPS0h8p2Ohu4EdkF6D8AzhEAfHLhVILtt+LsA
iCPWFNT2Tmp/lCGd6+Iq5qUr2z2GQ6CUYNd3aJoBkVzextMWuHzLWuLT0EYhhvmFFh68qGD7aL/A
56JeErUIdXCOCsJpsoollTZBZtvtIcVpPsyP0gW459s+SOFoq35qXnNwMgkuovNOuwkacrktnZdh
+nR8OKo+XRcNxQ7cYcG1zMZmMc6focmptymjBwnPZeKykdxJ2cOAYs8EkPrlFh7UQMqR7N4NjrY9
yIef11cBlchKUfA0rmxVcixa28UaJskSUR5keB7lgmtF38HB2VZsfYZeHcDwgisShHmklE5g5zqv
802pghfxrLHO46YJe16EcqZJkFvsg5aS+5wWQDwxHLvkR77UXbPq+fRSpW3JDy2KXLfe8oWeGWu9
TtR5yoMGb9zANi1h1O5J71vY0o19xpWBi6vIBp5PmcW8GiFKbEI+l8SRD4w870agLVagKApRbErz
ZWqhLdbHs5iIs+KHKxstLxFTeYi9Y3LojeIrm8LAiCyeMIKi+LXLQaEy3E0RwFrkj7tCTnH6xuCr
k4XbcBn2VCxlI1NDfcR5iKgPHp017zDlMBwUVMJ+7/Emh+KZNrfMGqdVvxj7wMZdCW5rM9W8xF1b
vgPVV9mC1PyuRu1Z9AAhA0lyAYmCln4SqpN9yz+/Ef9CHaR/ELH7BtchHrd4s1H0zSvPCfzRK5Qd
FbguEd8EgdOh6kI+uifbXPyOO/XPw0KYan+73YBRnpc5M78uMlOT8p0T82tVYEJkeYafHCcLLPr1
huDL2yU3dB1ofNvEJRGQiPlhGVgKKTz1zTYJPyNaE9QjmSgNBzHtWiHKXzRiftsJ3/oSCCqD2uBd
DVw0+wR7xscuvIrTrD3rVtbExDEeTVrvIIbjnCL4TmjO9xYhaUNha41PFSEjaJpdyTb48UGSzsef
ZKIXherGPUowwN9oJ9akI/+aNeTXwx4NTVG41qM0J5necUii3+i6Nces/pQD58jw+vNPjRdNSXU+
RIuN3ssysBiZzukKjai70Go5IphC274cX09Z7G38NtVoMpSTXLliewgwqD2CLyXtvNLc3xYpW4Z1
YGGYasJW1RRIZtkA2ouq+2Hq6en1/1HwjSr9Fn26LpoBkakTEiakN3BWd+Z2RXGMSSYVCULXtMoi
sFNl1lzNZu94sW3IrTfw6MaeyR1X/smaAfEfRWpt9IP9zqLqMeIu4pdLG/4By0nc8Jr0J6Uo+Xil
H3e2E6Bi1Wr+ICn+jX/OaPj6Laf+SoumBRr6DpmsbOzE9MgYTpgAC5N7MaTVouzeSmMlIBBdhJL1
SCvda1QrxUcmCw9M16kd4m0n/1aKCF2KVlLvNAznzcH3G+wG/anHVcSy/YOyAwnhS/jrubmZh0bo
DBxLhPowF6PFRfVu9UjQo1wmkQt3RdDBaoAQiOBUKgj31QDiZOG9GvBbicU/AA4O9u5W8h+YD2QW
Qd4L9fEIdvu0GxBIAnfWhlb8cvIJ6k09HURPW1kSdp2gwQTqjaivf7q+JKMoTMTbvL+kX79kbkms
Q1rDc3ktzZPrP7mee9auvDh0xCWwYpWyWOIjR17NCDcKswzcFEvtwiZgHLlc67PM0yI4EkmfNRtp
cFIihScnMWsKwXBwE7BorRUf3wvU5lPEngLAWOosFge/LArif7ACD8YnDM4X04ToJQN5dEHaYu1E
7op+I6F+i8+HDdH0MYBiKqhkzdXmH1172LIwwysV/XCgXL4mkkbhBnAl7qoPAoFLAqVwpXBnDnEx
kJgKEZnM/om92fFwTUyr4CgnMYGF3yqK8MmTQcES2NKpbEeMJgu4BzrFY7v35RtRSkm/QNJ0kRbT
YisFsTVGpv5OiVDNi3DyspK8VKyuwk/Pm8ggheo3JSc8dO4914MgZP3OxFyqs3S29GWZaOlP55fm
92aJcGUAEliATFVC2zn6hLwiVw5gUU4d93CnpR0CIqNxf7CuT8Bt5P9pfsQe3DRXni5apiT/croG
+diy/7ZpblZK0atCiP/ZuARq3OdaIY2qkeNZXkXAvyn/YyYIj1DlZTFnC2MKTj1DWEC/ezx7bw76
mjyr1J/pS1cxYaS7AICm0tLInjxshXwCg8SGFTEyj+XXk3crN6Smcsm+eNF7oeUBF5auRXH7FvFO
mo76VkOfdtmz3soac8Crc3lb05enqLRXdWDnKbZvPsG4cZKfgxHdtCSgwU56A6yXdBczekkDLMq6
ahDDa6664Ru3hOGDsJer7ExsY3t1G0BKV8Bgw4Dpej8c2qW/ct9LVrxjbIck9xGTabbfT/ah0OEU
BgtWsGdkw26pH39kfqHyOhTvAiaP6R65JJgEVq6EWfPwcsdam3b/YVpC8OBLduXM2StsZxslT60M
kynaiQ7P3blAUPwI0plS3JZTVeyegXv/DN3y51oCBpQW6+nvy/3w5UPEgysyZ2VsvOg+BW0KlXyo
2sfA0HVSIOpPJy5Igcpj6VGkbsGaOm6i572Z03wUx2snJO1KOyxh/Oq9PmiyZ1bRuCjY2zBAtB4e
uaFLipCw28Tf15fEpQZ6vQOdrM9xRTZ0kuVZgYtPy+tzr7iuwHvQl/QinRUPRQSJ1XZC1bY0omlj
O6vJjeth5IhF9/IlrtxaCzzBGrYLFYfWBrab3k72pfX8a+jSvL/0oUbGIZChW/+Pwvfunw1nSjXF
PyZCpwiNs2X1cKZEoycliVtGUZ0x34RII3l7yUVspJwLbFfgGinjdVjibJfC4ZoOChv8r+pk088l
Yx86G2vGiDib2OexWQWpRWp8JR6YY6MgLjK5KEF5L8jn54ogimaQNLMpbEzKRA8umkeXO/9A0A2e
Rx3OCrZtyi9vCBJRsaCmzXDe76C4luFcfdYeYlhq1mRcO2Y4RufefYN+RSZwAiV4pBDN92m4QlOm
hkIGsKlZPz69W8fWRgYDOC0ECPvfUHIv3DmscYK1y1tZUpZRHi0KThEHK+7c3idjYnWzkEeov0b3
LXMg8cG7TJkMvtDnJ4HM5J5EKbDntJkbba1aZC4TQfyLTmAi0Iuk4dESrNoMdJLDwjxOCy4F7mZ3
hN+kvnybMcRsdQHgcwCzFJZmFmgGjPI2Dcp+CFj9NfVRO0PXB2YDkSp2NgUrgEQeS85KZYZFLuMx
k6uwzoApU7Jsssa4UUO3CMi32TIjgZ9LBcxeWJdc29wMi+is1zTO/D9Taiys1qwAtTChj8JIVNxt
J2icpM20v/WRcc3gC/YbB1Ycse+Jjb2WZ14j+ar5eiyVP06IcG7ub7mDovvT0dDPnhexz6duQzj/
SiSPIoUK/BanUDai0YKWDOMtlDbDXN9LxJZjNKrXZHg81mK61/vc9k24Huoy1XVig5W8zQ5k4DWE
rjnqqMYxHr3sG3PmELTVXaDFs3NWDLXtpcFDdVM91bq3GYgaYoMZuKxNLqeN2NEJSZl8tT7kF3wn
IJNZgQ5u+GqIB+7ML2B36MWzapmr5MLXHjwVcB5BbBDFh7cxSOlyq0IeFzRC5b57jssda26AT6+K
mBq7M6e27c+UvyO1HcX9NABCZPEIXQDan7FAfyXdqFJw7LtYxAorkgDcmCygQBS/ZNMJfz19HMD1
He5nnTccYRvDarDt+u9v62f3CsQqOQi2Yi3KvWs5yHz5ZDmWLC3hCcrcnG5j/wVpV9eQ0ffJ0PKW
d8Z+8roFG+GkaVi1iDfUwCIMeXJy0Z8jS/wtjKSz4/+UV3SPNRstiqI+tK8suv/zB9AbbmkHL7Ft
2Iu8bh8SL9lfE3jKV9qdI62zbMG05YsgWs++gbFHeVlgIgj+jIa5u9F7ryV1Itl3rMn0hd2IsiLh
x0qv7CHvPFXKxRc0cefvDwjlaKzCUnbQDzw5HxFYmy9j822MHeLoi0+zLOz0K5NbIVFV7F8o+YAS
OKUmZrVVB13rwM6QpdA81SaoBAvHspjpGUs2EhMm8ewdhvfIrwZGP7l+A3AM062pJwiRL5V90Xpa
d7OMviIT+AnjWLSKaMEUBWhH1M79p5bBoEwFxj89Gnl+u8kp3kTd2hpiVhMGcDWcjPSDHMlbC83W
UeEBmEcZGGUCeHgxGP8RoVklZZMYT90D77G/N1ZCAcAAYGucsVVzHZuMR20GEgsiTBSR8l2Zjwsz
OEnHgrnT2r0KT1kxSsyosALPgQkLfwn4pZkjyAoGaZWs8fq+mOQ2NKGnCQMN+6hBBMSshOnuUSAw
x437gC5HA9MiScR/6ymEqskkF+TxhEWxQYM9QR9/EwWijQjhHMPOA0dRmVRlIkxPx6R7OpqT2dgb
urSnVzyj9Vw47bc91FXSI1h6V2WdXQhXzzOQJSvnjYHpcc7JG2FX5RDAyPJF3tN8CG7Zf/y9WD0F
/1PCAJvlplne3muPO6u8YEi5ap7dKx/hvqzDzabUQqlk8+S6gSVLnTGGPVj635IQeMl063QGlD06
qhA7fSVxXl29RCswlB9Jewsvf8ZsfszIux4VyfEix8EITKUzbI6jmqK3kWmnqr6KaZNVOjy3qClU
4Tv4eiBlDrczHERo/Cbu6gLZSVZ92SuBl0/vP8MVNtgNSO7598UOIsP/a4AHd42xgeaoxdN/qw8x
TG+6y5hWynpdyd96YdfOz4owoOuusF9EUVttXmlz0MALavr+BYF0EGYTQVeTiOSs50hre+xODkvl
3o4xJMRtwOhOUcluTis9+1m5o/RhJ0gd5kTyLA+647FWkIX3IqDn3e7aC1pXk9aDcxDdRbMelKwS
KbLUcnTxzF5cLRbgklGZtunvqnR6Asm09wSMrcx22kd+Ka9Jg0Ivbu8j30x4jKLOpRAJKjgshnyw
8FkPAPX6mZlBCMxrJNnBsAX3lPZZjigEtVkLQmBI/pzPMMQEH1AzmuV+cFHwT5Xus2ryHzLmPWoE
kD8HsdNfLVx8bjvBg5rRETNzjLLdH+mfeHFt4RpEJ0bsXmFO7r5HiCu+VnbNZhi8OLu9rj/GuUOs
kPnneCLAZQj/e9ATmHbGnWpytuxpqaba4NRQwWb+3t3fIs2F0jSr2vXhwtlc46qmj4eMOYioKz3I
huaiT5nuSaYUdcd6I6SyVoNJLJ8vAS3KzehbNZIhmS3qQeip1VYeHINXp1JBOtu09aeL/B3If9va
g6zMAxsRvsU93QlUy7x8fZLkI/nvnlpKRCHS7FoNslGxTrlXFycwNvqncgU9Xek5JqweuskDYhZe
q5GMEo/tf6JsCFihJ+9BEiFhyJBgbRwPL92Vog8boH8Jki8fmg0mmpcm8sXpUWpPST8zhgqTArHJ
Gn3ycsIbDqeD75mlTOb5DJlX72vMJJBYP2tu49GhqqaBixldir8fzSlTrI04ygNab8hITR2RWDeu
2zjTt571uph1Lqc5SvqvCkyh4j8qTBWC/2pU2Lp34eEviUDmBSCAT4+OXBcE/kVboxovZW5PHfKX
JJwuXNipAfJajTF/SIOXChNsiqe5CLsE7MJqcBqnWUmaN/jFMFjtiJMuXMEW/+8AxtQx+/hRoPM8
mCvUDKdEllo7bynlorne9E8zbCNRHEaVtxQZ3yLpu9EzhMdZn1i6Snv78YbRMyiVHVpNFTartCUB
4QRMQXPEKh61gU1jYEHXujw93vdBNqi+K15/ZXkxLx5NcWgqRm9KM82sNf24MVlku/BfXWPUNTSy
aZRM9os9mlD07tlccQPRG5WWK1/WqQNNJ34pR1QYDsIqSVXLl57iLeAk+0Y4qWDoVKZSrH0q+psL
LjgYJgOjdZwtDbvSKJyVstp/fz8zllOWWCcj53s0GPXQjwqGU+Si0towfUQC4wondJrWHsMVeINz
nTp2tLD9IZXVxQWoQGusl5G7l/ChgGfbkG0C4Tnq2sq8WmPstGZ3Gh5584vluAwrIl+8kukrbntk
Ir9jbPAd+2cfc0sKjMNr9TlqRYW/3r6LUDBUyjsHnh/TApwQOKuHtG10gMnySxS8S70VKUTaHVYF
K8y1GvPwkJNeDp0rS9O/LH4w0SCBs/nqdDY3dZN2VZ8Ewl382YqSbtoN+X6iEvwImaQFGCnlNMUu
ujVXnBFUxlOLa+6piB3YnlHuH9SNJ2uB0JGFkwMoXISsy23n4VbmEuSHBRGCickC9JATm6M0fDUQ
mWBmS+II+RFB0rplCyttHhP7BDftgdbshQJDTqJM17XLqV9rrXmdGRhyeu9G3JBuyo1AdG3dJNk+
TQ6cGxbI8nfCnFFfyZlSISfjouXfBAosG/HEXcpVxjlfrVAusyW71CqsI9YZJqUmLzzp0stux8Hz
wauYmTd9xhdV9AK9tJRp4dkctzOloavRuIFPMYfy4hAfisZxehH5BARWpPDhPTR1sZ4Qy6Bs6ASn
OzWgyLJVkt/uwSGw4sbrA/uUN+/+yHl+CVdxQ4qmxwOQ6tpVIW3D+frF/KYf9KzB5GxrTbiWIADD
tigShWCbUi8IxxP3v8O+A35ygtx2YnZIwBYm5I3sb4EknZS5+uOtvLqTwzE4fLGuX0Vej3Mtmx/w
ORDCHM1wWYvlWXr45Nfnt1f1QHppdnQNKV+/HjNRRcJqE4z48HmVI7BFMWn14GdiDqJ13XO/qEuQ
Fn6GomT/otQuscxFXpVNO5tH3Hd2bwjwZN3soNziq3uLQgJjUSDUd6PrK9J/g83qHfejCN999zat
wK8CRq97aE8EvON+Pfq5OcS8li3fR1VWwsBGq3gw5axkeclaqSmHYOqQfRtLGY9EuBH5TTKn0WlR
QKjvfJK2NqwWX9CFyeU8h1MfiYpIaNo9clLjWgiGOWNT9QUbPVr0y5oP82SP+Y1Cxa14CDot8VdU
bC4fLFMgsGBBAIKA8nZdGyrY7SL/h246Ajo2AKbB6A1FvTZVDqEf2PijR35y/QCn5XdcM5yVUc4l
K/gHvhHUKy/gtDEB3XyInXpBxKwec7SO5lAy1KfG52f9RWHyQv1kaETu7mDD2sE6NPwL5lqfdGBU
l/JEftEVcwKTheBkcr4aaNnJmuJTp0ci7e0s7crOf/lhUK9VhEi04BF69eKEsLVTaUuSXBzP5ZKU
jDOXLtRx26Ih5kubDYzh8mDAX9a81MrKHaKvoi3zkFk6kOsxUUDO0IirjkUtj2hycMZ9DLxPmTrP
P1ogFCIJ1hQcglHYH6Py2alMKQFx9souPoECBipD9XVc//Y1Ufz0tqbir1gSe2IOhIFzz5YIfLwt
d50Dyv1OoRrMR41bYQxJJFRURhT7SGQXn3Rkh4iu3vAsWNXeADAylEvjz4EIpaw5UCVxumIALkB1
UtItLDKrm8oeYxhvkz1R4Iz6eB7iQSlYMnycTTyY2w/W2XX0cNCnwkWfHZXfUIrt6+OdBomv7vwh
h2euvnpS8q/T4GKd9croZ8drC2Yd3kOevxFrG7VeWPaqeBQZuJf0rl5DdqV7SNiZom8/TMcmUKGo
S5BowXv5e5oXF5bTqkyafx9+vEcD+BAlcXTIpCqiolLIm1LAyVekZNTKS1SOy4E6pW/npLskTC8W
8vBhFLBdxXZtFkBbF/WGUkzDFy4V9IS/c2toZUKM2qgCjOzmsdGyTEaP3Cal80MprgZSOsDya0X0
sD5DUf1ga7mKurzXhOXOAie5IxSaDlbL/Ohi4LL+e3G+zjMBG1TutzIb+vhtgDSPr8zp1PqGoXCS
Sp3C9TqCUFvcOYGl28HSui5A7jrdeHPzmVbzqKa4nvTxuV1sLkniBZM27IAG0TV5Q8GzruBBFPhi
D6bc/v91fIpuVXs7IUL/MuRVgUpDosDYPnAZ+X5sA5pcjJT/Nr5ZOHUkUr6Gay5QPvzysJmRESLb
5PGIaEg7u1y49uEOEYOkwW0QpK/a8SWTsVQet01Sbj3X4gDUMbstqhJjg6UWC04KBBoZnEiqpy6Q
aNATHV2dnhcA5HyD3/TtD2NvTVcG7f6ZCicrnumVmgvfw9fsu4A2I+GCjm+EJ0JtVbU3NhqimAIT
Rajm8tmTGCoS47qK5GXIwb8OncIMpI8aFd7hry9niFIwFDIP1GHzn9U2zhkAll6GRUf9m/AjUQIO
iL3QM3z6ocUwaWGPXWxpCdZfsjN1kUrCISEpawJSdM/Ijoeceju3hEPr2jeALq/Ek4n7GUu4wLuE
1AYNA9DKKMbpJYRZyUN/vR6n6OfE/mjqxSTYNEcb1RlK2Pk7EE/HWbAjAf3VfPXhCJCCi4/2ec2O
mtkQZS3dk/3ilOIYtMapdr7wGNzW5zold+bbzbkH9pTw+jtLZ/FAN8cUjNFMlHsWuO5u2m13rZxN
717K9DxJlkC460omDRxkNOCMiD2STx363mVxJ9M1DnZioAhcoGEaX8pVuq+be/PnOKXMZBwgzFXq
xlZGjxcnm7NgOxXr1cZshmdHd7vWoSO2oVOuW9aXhWPKorDKAhW2o0A6fnBnphAbCfqiSPW2bjR+
ym2WC32vIO5PLWs47OLcx3LjnBXXtOk1Fsr8ZHk3zyM7pn792Z4sw+DhEC2KQ3BKT1hropqd+rUt
hfn3RGx3I8QTxK5p+kMV4D0IKDV53SGF76AH/2eI27fNV1XJahGcZX6i7WIEyruRN8yTvJz25La9
gxARJwq3APdfHRmDVaC0oBIzXmVC0Ad5dw1fiYm60+sIG+itUhR26oyWxi6wkEJKhmujnzSSFVd3
l+g5fsPgczOMwxbgfDlBrwHCVU+8+unElvri+pv+de+ZRI/FaxplDoF9FANrh8Vaasvrl92YGUvS
QKI3zWAaEBWGm+qDgjnn+XPQsNPqSnWeLVKcNf3BHqsEnWyMXzSgrZQpEKa6bMq8Zy+7Hd6NuG4n
gE3KPBiFaOhf/4IVAOYqOh3JPILmayhki8zwtXr1nLg8P/TiKP7lt+G9VY9HuYyQ3DrlPWDhG+VG
IIB2Z1ObMznavPpeU/NX+mVZzSg5EAsKxpvyv4JY/8695vyQ7HHOAwhHeBCrGZjS2Z4/BEluOXhW
J0T0TSI/IKKA5ZjVHPxWM0uQEKwwfVq3te8RemIDThswe65BDobpF3ZDWJnJUfbGWZ4ZVyfUpc4z
ZbazVZ++8fTkELLbbXsevdBCSbJte0gbsC1XMrc+ph8su0jiEJ1gR/xf3VbaNElRKERCJ+m7O8Ih
DvYElzYsxP9ReIt94fCBOEKhs2WMu7RKLnugne8ddw8Woeg4lHXaB4pvq6TYD0EqDpEDYbrzyP0r
nC6ROWELRHnB4Gz2D+hgdHue5ONPlPJUmy6zJrUA8FyLm8twRkzBGsSjxu0mC+40jDo/QgSApY0c
xx1jbup97znULwl+SD8CaZL/uKBryiOECD5z2mE4mwLYkykstN8cbjDLQvonkfHWombJTNyvLERM
d4yuBtX7J3W3g8hdx9kjk0P9mab7fsYV1VqsL4rkIglYITXG+ZDqkXQ/pXdCtZUNm5VHgafoN9/m
Z2HIo0QZo4xMKjhxgS4XBvxYapYyVRujXrRDImawVCNXV8h+eynNkhxRqVFOONSuvXJWutgWoTDN
rGfdwd1ZKZ2LIDMH+GpRvwlVWoEtG1rm6SRTQmV/O6X+9yf9Lz+w21bbsUZm0kXIf26voLVAMIqC
YUGzuFwgfH2kU7ll5RiqspM2IcrwPSYeULl9VXqBnvahBL83C/RlLpD4gCxHoPexfzJzAoPAE+B8
Upd7FEPcYOUrzOTUjtUOUSPC1V1BDRWhY0cODMglqBn/UEV6FG35ql4SXulD5QYwjOvXVrPpWlSb
S83G82gjUIqpNNLItzfvDKRzb7IiXj+RA/KpvgIYHmXBWzu0nl6bPPbnbJPD8lR+BfTIMDDknZsb
8v9ArWrxzqgoRb98/bKSl4ANHuqaq1anfmbBhCphvG01gzGcknDKsVFzPJBLFcXQww+NPJcPfaXE
JfO5z8kBpQeaY3qCPBDJOmvDMs9wDy/Bc0ApFbiiTAkNxSQ5/6MPS1L7hMtcwGRax2TLya6r6bzL
f3JWOgWyQ10NFhBXfVvHdIyRwD9AyoLZWRVS3JmC7VoFo1miIrocjazyQKTlRAhWO/KlYx/B41BC
I+bF0ME9/Pd+fg7cp9nYv4jly03gut9G210zpXHrplXU7XExjwJEbASN0gLVx//yqb73LVGKGo6Q
RZI1Lzc+OuT5eLiQRg7Vp5Bcu/J9q8JlsG/+QI9Qv2wSZhdkW3lEo/3Q//4bralskQqpVPu6loLu
weJUKFNe/hvAwkRB0Xd/wPheNV5JM8N83lB3xgfGCAzTcXpEzBUEYnG56IIU++/H/B08101nAcs0
i4D8GkVnAJvGAxq6WlI6snuaMfQhuaH07ISaCoyWLBiY2pHyBK+9542SELMCSynKt7cFL6Px/C7j
KeTm3NugGiu6SCicyXLX17oH/Kid7oM1mM6/qsINHKrA31Bu2H0RXA9Udqyqp3XjK5XUYidf7M2d
C/FdB7+deAJDUbhUunJtH+WTa/hb0+jLU5nGsK8IM49tMMYfbR0FEGFIU2zq+Gkl/qdoxoV0P+vN
yrZj6vkklsbHgX86MZ1cCrVm+a2+kdbV4C3dCh398e/KkhdLk6cvuYo6T/1V/Nfhg10NkEXL7IRw
MNaWOPzBWet2nFijv4lvW7meL9aJiNwVtr9x9X0qcwGOO4qHwRRGsSuu8OI52dvib63BP5lJo34e
ey/yUb/92xt9sZawqr1nWJHweoab7GybkDWjL4S6Lru9I4EYhl3TaIQQEs4BVmuQ6jX3sQ6ufMnI
YSzTVrEhU3TEwwUa+5I9fPBtT3Or+R1hkP1vyv3QP1fNHbRls9P5utWRBXp+PpZBvG9lKzIYT3sw
MiKOGDYsUIMBh/Vaoi+LxkoSwLAAejZLY5zfyN5nrSDsMChL0dI9SzYf3K+wZhfDlxFsOlxXtF6Y
Zvw2IR76fAsU/7jskq2K4Gje7xr14fdZx5SfWXnzv+QFO03OrtHE/blQ8QKk7jNaz3Z9uEA9jeD+
abmpF8jcnGj044/YdKI9z1cBqNmMoIyTCyU8RvyqTA6/WaCeO/dVyxB7F5+sUTo/5U7JHl3goo1p
ZQlkLodZkn6FmYau24nKAs31STMXDuSxdbesuE8WVul36c0D2p3JV8dB1dZJT+0wL+Z3Ey52bMO6
XJKQV3U2WmdgmZzhuGi5PVZ0hb4nz01ndx8eKhGrFgTBEck59PbzR8LegUIjLEp0xxpDW8pNxltm
e/WI+TRja00AHU8CguGYYmuAt5/M67elLkTExArG+6w8QjdwdvZmU0mYr6aUWuzPUEc4dsFVkD7m
PX9T+VLg18mzeCFe6++Hy+q7m0h8oXmsgej8ErIwgr66tL5lCsAvzrJnZyv8CsyN6kY27kZRlezj
gOI+mU/pMO+lcjzEYa1aUkbi1EJUa10zK21bGsIaMPN8QCDEWaP6+2Ef7mH26FwbX7iClrrv3j20
2miA+kgfHe0b5KAFMJfbHzN5KGcJR7U+RJ0epETkJSIlnjhjmvLEBUrmbfdMn9oCGMZiNnzYr8CV
JKmG4rc0JKe3Fz9puGpzxcauIAKra/GPlVfsvaDOWflv/mm/gTPasqyEdqHtO2rTnySct4QhZz/Q
HG6cZknlgeVx7bwwGVJ4NNywb0zd2Jh5fJUqmpk3jCG1x1HPYdipDv9E6nZVWCtRgOE49UoWsBTF
7YdAcLP2pBfYB/JMgwX1pgd01Lf2hyNHf2BLz5MzhP9c25dTlf2XW03EK7HpDXrH7fsUyRsFPd6l
WOXTx/MqfuAO9FUme9tLVPFDqKcfj8YX/jeGEk0kM/FcR49L3DtY4q9jK8sslSRbtWkSzdhgrb/M
pNyVtM241NkPqQSEmmpRT7hwbYaBSRL0L7MWpn4uVeAHdQguhMnoXGjz8/QZW92CISCs3Q9Qdvqj
l+xObwvP+yFXwE2Nc/LuZXOczysPask6jbPN+4foVQB35tmRjfmyUpS7+OSys52qUre1hRsRfEnP
6ghmH053IbNcNkY9z8iDwU9ZdPbxAaAKZB8VbB7zmyDKIjD7KURVSitY42frwIMsRXmQrFMkTKoc
u0ExPA/zuFB/PDUvTwT8VJbkUH9/dU0QgedRSbCcb7G+oWkb3Pa4GC05IceOwFe9UWPab/g7PTmH
t+aPVDr7qMx1Gg2e7Thy5AgdGf1dVNPvMwKXPJhQ51ZEPBY7IAJcyaeHqjUd0eFScaVRkPMN5JSe
+FmbfOnvZ+cuVEOm+dybe/4nPsQybgQkXpdtJH8szJPpR9qB5+A81518LX2KM7AqLV/SP8gbonhc
UqVEzRdf7g5HJ1aPW9YutxVzhrOL48VAXEC/brrceXLKZ8DhEQQ4vurcbhZE4wtp6jLu4tINKI/J
HAyKy2l1renHxOAd6AVat9oxwhU5Kd86FcJLKMeff9sze+iCYs5z31Y2iV7kOaJLbVMUEnOXMrt0
OMdT4a8RZqaEg/p3vDe81i4kU6E8LsuEoc6XPIFieMkHXKlt5wHw8KOxyfqhiHvlcJxLiUmyF2FL
Gh6ZW5LaNnpgC5I4MyHJjPvid4rMm8Jg2wZYhUzwUO02l+4jRJEjlvka6kLHwcmihgGca8uC6R6r
6RyGabGCiLhDJXa4E/5x78xFPrPZmIu85R5sdzDdj3sImNzuGRTOi0bWAfFfoF82yWw/awKSOAe4
hv/aBuTLf2QLKTKqZl1qPXwWrjpdAZ+Cc0l2WYdwZO+drA3mtGB5YDY1se5UMCfXvQMwSFltGsHy
6W7yI/u37Gf8YaPAnlzHeTU1oaiPsagGCBdH0b3OIpBMoqra4na5SDlWf8e2tffvr2A7IOnxCQsa
th3KMJAh8CSPEypb6RvjMbyju6VGIPmog7q7bptoaByDe55QIHcPp9HMiUhF4btzVvj7npt3RRdc
uyxDWagHrhFqI9jr7/DjeFNNy8lBSWL8P5N375QyUU6kjicgjJtCk3tXnTNfIKyoXqP/uSa4LdxR
jCtj/IbT4Skna3o0+ajg6aLLFzJM14q2d25GslZzovSpKfv3k9LHmG8y19EgCpxnsKNS2QXlLqgA
HLKqgwX0O77jpCyUIQvh1Dc34VttmxU0dfAfUouArZkzLCj1PQzwt8Gf6/bCTG0JcWqeT8rH4uf0
1VVHIsW+45PBV9ptXZtWCmPT3UMNOD6+9DuAiT85M/uDGu9YttKzZmNMb9qH6Lzhy9BmD/I0oiV+
gMNJi/jOjMpqQHgwDxucjFAviESPVTQvnZZha1sPmX0qjuiK+kE3ELPXY0todv72NGrAyqXafvMj
bO1lEt1Ll2i91NJflJhXYlWYJfE7IQoUxlNP3/3Uz8TRiakk82j8x8BD7DBeCZLETvKgQljvM3/K
d2++2QlhW/ekm5YFHw7PAFwJ8n569Wz8kiUWIZf5qSTy6cbDftT2v3OwzkgJkn7oAD/2xFFCormv
Ai5FbGWl3zLRgNReGsFhgGdyLY1UhERp/RTPL/qxLBb0BfHPlZzc41zMANb3TovO27Iao3Zs4UuE
IgcwB3xHXYkmG4nBjuviDZqYwUrxijZg+zPSwX1JjQtiRrYgkMIffVwp5O0uJ5ZFDEBQWDuN2BMc
o+K1/JTGyf6fPgEeCA2buEim9377p4wrRfapWijVpq8yVQ64MfdkSXrO7ch9lYab6ucaIZZ/BIM3
K6H6Xwq8u0hqOjswCbJv8vb6cFZGEA1JhDNTVusKVxUrTLq/0csYUunuS/eMM9baXArf6tUcl8HN
sFxZKZx8vM9oxxd4gXhBq5tyvY2rtB33Ufzn2SR7YNFYbsqVTODJT9Oi6ZFCQDYQynNgsa1hlUbo
jWqn0gG7/etefGNjzpAaENH/NQ5L2ND6R6sQx+PBaFO+KsKYQQ4ngq4pSRGKTQq8/K1nfQtlcqCe
zEVRgOfQrwSg7ITMZ1uZKSnZTsmy9XUhTCkEf0ftEzFomH1tfXajo9RJ3IT7H+cTY5Vjx+XW4pL8
uyWQenFsn1v11/KJw2xprqNk4HYPBglOSWdmdqB2+WcGE+MCE5KxUzW9g0NOydfQtvunGpPfMiMb
A6KdB5xsrDhkY2Ts7s6pAUC9bJiyJg9/FuSaZqgf9lwOCi78YvwTcF8vbivI60czAajhdinOdQ+J
78rG9CUWa1L4JLxSrnW9gmr5R8jJtRd9VxSYO59+bFZiPGGG0C1WAk3PXECuUiy3a76EHdBWDh/Q
mh3n/WzWBjahJNrM819KysAkMzEtq72iwkaihpD45ArmQOSQzdTwf8WIepGJYrqr7KURyN6+HpPO
2vouyEzHdpjKatoOBgJrKCSGN7C0JLJ4MJeP+SWg8TfD4i0d7SHLeptMTEuntYhab/XcL4omyc/s
tdPHukRhmcWh3dXAGQ5bGEaVNB2lxGZaRZScbUHPgZAdyhcrb3PfiQXpAcLEVjxNbtZsRY3wABwV
Zs2pM4hBnIC3OcJWMjpJKMOd3YdLwKUSQP40PycbAIhcCS5lp4LeG8uBnqkJC8yH6tzf+Gdpar8h
WTevDnHofCUNPSAsrbkdVbw46g3c93GAOaoc8mpAUSnA7V9lgn8ipuZynBlvWLfnjYjDTHYSvj5i
TFsh8Ooumn+Jg7UZz0XXQkAUzZlp40IIL0l7Tx8Eq8ksYNjwej/XnsCOCgVZBRZEs+jpv+upGMlg
8Nvel91Mk+Ua9raFFARIAUl2nlk6iujfJAJVePJQfVNGwUS6JEFOt52LTlbe89doBCrbcu5eeTai
ZNmOQMeGRPQRfGMS39g1Gy/5teyF8tO5eBfd0CjOMbrWvUloNbGjytIPDuGANTPD0Sj/mQE0Xv1t
hL4HX7lDGO+iH9VxdTBabTviqdBuHDkGMJmFvrrn3DPm5JBwT2VdadRAI+BwKY3P+wmynLBYKot9
XfgHmGcUaQrDg+TiVW49pOB/4Zn8Pf7DxthRzNUA2kEtJK2YArAPA+BDk+F9ErWTEXlTDkoR3H1m
IWpTDvB3PxMImUjoAT0p+d1L8l2yxK19i9szSaYwkbkZEFHKIFSKj7JdgEuSLUzXDPQvHt31ygFW
gJnWynKBJUwWWTLdd18IPDNXSt4G42Er51TUibgGTaQ1kaCTrI3JSpMFXLHgPOSLwT2Spk44f0xP
dIKgo1TJOHZ/Uy8bz+cxnv3Hg+klEKZC4QU5Yv7j23iTsQXrB1kuLXnYO/IsjduCMQEMPkluvJGV
WBJcEpeLUPE+4WRNC89efKjZnMnuvWhxEaTwpA0cZRyOyh2g6/GhcykZKGgGa+r9oVy0SA1x374s
UhcybfFYUe+LQitDmdDSvxs49zaqcEvJwWVjMoiulcVWf0ZIbifQuyUWnDIgntuhpchLA4+a3llm
fNtYj97/hX19uCjSBLvkE6M2fxjas2Fkg9T9u6MU0mT6IWAp/vi1W5RZsLa9sEhpwoAP6en55BBQ
hOyYll/MiYoGMJHjSxb5MP5G1VeWN3f3/Jwlp6nZb/r/fDbg5tPLDxvSvGkzmaZjiU6UkQ48tkgp
gBvqIrx9EX/La6lzTORELGdcC3iSrsmVJlBPRqebFGUjCsgSHPOEQbqWRnqmglsqlsYlExW0ZTf6
Q7vLegAvvtILRbTecPW6esnXJWTYJ7PV7cpQans9/DsQ0RBL0XAXYmZuhTXhuMzZDLPCYsvFNoki
tPv6g85MbqhGQinnhLPeVIGSxDFysPrJzcKPOyOYCL+Oo5QtJkqdmg4wJe3sLNJujhQB2r2LqcBM
a+JuORNl9wP28iSM7pabZ3v/PMbsdXj2txuVVSe2jp5/vkJq3hdGCOOXejKq72ExyLDoqMhc/VnK
dAx7qHJQ0GkhLWqPgRJuCdwiLaNqU0TWeFYP4iRib8kzN/aQ+OGsXtD/cJaYijQ1roiO5X0CeAWe
y1AWD8ErBZ4UKlQBTHuordMCqIQZyExt56o7a1zAAvcEOwdSADTUKvDHHrMUB0bH3IVDZav0iMsh
4u87MhWwqRU4avDKKhRnPqHmOp6roa/ytC0FDObTAoAxKGsHrk0RQbvzl68ufufMYiqbIr1fPRzJ
iK4ginadKkqfuOqbEgzVlcni6OzGrdFPX3AZgByCrp1Zc9n1BrExachuD9eVrKtPD0JSXa7pEecY
bDr+K/wXXXzY6UG6QpnfG6SHD8iWWDsF54a2n5J0uNZwRCFDsfer4PkyQ4OGZME3bgbrWSRMT9wg
YNtXudzEuGC/L9/CvaXQXTNGdYuwu3bVSyHKBFiNYuqg47tbzRL2qSNsZb5hvnS3fYXICU3HhOso
bXHg+qrA0T5kRLHDXifH2EmZXlagQcj5mf6BFfQef0E46Bxcon5LxOKdCbCJX63DeBHpqgwJI8y2
6SfpCeHBInlBoCisIfseLIoPaSfybf+CsbH8bVEzfyokVGp7Aqz/CEq8scBqnqvCDgP8I5FEfGdc
7vqZ6hASrVPfAMBvlInxKc8CRQvLAGGTnGm2/QNXdOMdPfX1UrfCmVyLXtKQbo8TwEWdZrpaM5+1
6pmag+V5EQ5clYef2QwtKMKSG9TiaLgmO1w84pY/ilJNOI0d8RmnFzwUuQhsF/PU9byo13rIwUR2
nCQ18iOwySSK9KC+J2OH94OMTwIiqB+lZ4fUSnWLm2BucSMiAy4Qbcs8iLPet5tTkZ3GLrSC29UE
4L9syulDwcrr7yRvwzFAbNKAH6QOYflWml35T1IuA47IfmCPysZDCDiucSgWHQMiy/Rp5FpL1xRX
sXtrjb14+4dhJ6uuw8T7nzR/Vi+Dr+nnkp4IzQzy+NGQ+3ELZq9WxjihbwhgnnWCk58aPg/tD3EZ
5bTzUVQ1YDhqRznjuOj14BWTZtH5tRFq/xf5R7S9wn/B45kIVy+c1buh9SwjfH/TsTvxCxNWKWif
U6kfLeYJ2YDONnDwN73TGmBduerrHH7cH9ACW68ihX0XzjbfJab411+UwPWpd+ejNggkorqFFXaY
5VM3L0t9Y0Dq1qFryYkwbxpSJtnPuBc1NG4NqgY2W2fg0lKdzZCIsoC8JWlzou2jlAF+QqdGnwmR
zLowK5oDYvLfmAyDP/oHYS7/jvSR0Ik1o+NJudEtTp/B3lj+JwvfspSJqVez7S6n5FCMSsN03US7
KorO7xEmPkUVevNE+RWc4FqniKIIkoIdW109d7KCgyRrNYIN5p9vDxRp1leAWWccMgzyKqrgab3g
cYlB+epWvsbLvjHAyE7WX5UVdMCtpC0lk8xBhPKirjx29NII5ACe8YIPT2rgJSAQRgtTX7S9h/2l
H6tvLiNCztsrrE8RpSSV81+dndPkelmv/qXxoQBVhzBTAI90bKzBdBsxN+JKB9hFsDwiYApMZCSL
KiD6a0lkTeqen8qx8+4ST7IfeQR0sLDHBB0OvW6PBTnRdvKHk2BJAw8bXZQaqAuVbEQ6/fq8XU4a
LZl0VmYIOR3AlNG5ZygT6OttaeNVJnkiPnouaoUz8zfsIdwPGRJwRLjjYbmBNZYDz1I3wTrAyHtC
IEpCdM6tPL7u1QPC8rmTpYploupCMKQarISN3JCkH66ZF1dY4lpA2Tvcfe683VxhWtgpg+bHPB85
8lQVUUjgy4jIQoZ7QzEU9/X1LE2MQp0J38+w5EGBrEa85weBkBNTMgmeiE2pTgvnQ3BIl2+JJYGE
RqFBvCNW7BwbO/wlWQ6Bjjr2pCiTOAetku1Evx0+s6fKcHJ/3ovVyzfgINBkxl5qesOvFBpmmF9a
zSjEeYIYZ+tp8gRiosb8gWOTxMGOEzi0tefNWCFf9F2YxIZr0HdVrD1EZkf/etZQ7g+2aqK95eE8
GkHFrXcMd7WeMwVOvTpsoOTy7C4EbQPm25T6Z1KIux0mhacTDfPODd8+gc1CCYJfigcGYAbJJoIY
OX92bCNXsQ4upCnXajDMvMAWO9eims2ZT1AD27Yq/vIoy0CMRrDCHQDxSwc4g4u97Pha7YvC6aGI
sg9vbh0bnWmJVzYH3fVJN17dSXa2jpb6PmPEhjKsUO5xXAwpl7I53dfApAa0LP+a1PwGkPSpwu+h
wZdZs16s4OwrmDlGanEjWVg+Zam7m5AYQNnz9XtGHlS4JYyJJgCLc6rXRdmC5ebFm9wawf88Gvzy
KgmmPAnwdRwfHYZQNqTE2DMxrAv1AHS2kVIymvYiobhACMhaQOu6u5cpkaOkjPjkv7o8kckXBzxV
0kvb19GDSkxCfOd5bB7nHGSG0rRJG4fCySZ1mPTqdt7w1n588BiMQX6JvVmOefKsAp0OnbQZTBQ+
mzP+wb5x+eXb7Q+IUrPacRyf+Qvyl8No+wHc99FXL4UDfPn57RBhfqo75F2oMhLWceAHkyI5f0Px
AQBWx+A5M5kSeFOL7W8KLM86oZahpmLdY8Vzr1/CvYiUMg5WXdblzl4EnysES2U7gKlUyp13VYrP
xLcOoNdY8IySq4AkAt//8HehlXVBRu+UC86qaVPqcMSlu948QON4YKydWS/jO1KWLWGjxglUGPyO
KUDfZXtQ3jZKMDfQP7k0ht/JBGk7LBJmpWzizxMtpqz6WJg2bPFjHy4GQ4Dz/cWYJCjy7hErYxyC
SIqsvlXY6sx6mrdTopsnQwL7f7uNq9m9NPdFSn1kU5QD/cDkDgF4nwkW8p0DEUJxd/xO1hzyEpGE
8td6SpsafeLJMNImLnP1pEns3WOsuhA9Vjw8W49kv80JqA2lB9ph1gRcmXeojTf30gIPv7JnlXth
2tUgcD5Q/wOpbV266wVyX9nKzh35+1Hz5CI0xTkho7HZO/+zzl9h/8zPodY3F6bAsjEJtV6tQ9P9
XURcv6t64G8eSTWuuC+88E8mM1m2rN40U2hMkpqiS4+HkVdqvgZOG/vGHRroec6kevzI1E6SVihY
7lnMgjd1F3NS4FeKgvCZvP/VKg20/uUKT1Wu68jgNfgiK6y89lQef2xT6acelVOsfWzeUNg9dRqE
lhbpbKK8PDwyOaY8UBzFsF2ZC8SYfQJdTdnC3OdaEofmdxE5zz0X48psuasIBCarGR6QCGouT1wr
5vA5jJf03UexCx+1b2qFfvyMqSSboR37ncIc6lJYp1JEIEAVb0h9XlS10fgwc7jg4hwUvkLob5JB
craNTiL7R7RYH+sFIYXUiTfIcoHfUk/aCMtzjkHhgMsLssY6IF+pxBoCUJh/wLwCR3kbp2Sda/p6
nOakb/gVL6npLIA6T5EkL2XhshQVyz1pSjEYgIK6tQsqqw8KqZgeB+DLCzh6nC1uMulLPwGaLe0Y
er5a0OVqBlSMqYxY4wXpHnDIr5sC3ISeSJzYKIqW5iHw++LtEL1+oEhmv8pQu8/5qFfszzqI9/u5
5vF8KHnxzHVe4kWSv27RcPLiPEl+156/WjorWeT8n/F2S+niQI1w//7RHBmLMFrbeS0ztK7CH3vr
RXlN5Ea8d6cfj1y39/T1wznqSB1Cke8U2ys09egdx7X5Uj5RPiFXqPv5/eJFndykef7T2SkNJEy1
+csr65cn8bfEMQ7DltP9Vgqio0ZYJZADMB2XnPa7nuk/m2AS28OLi8g4n20uHoZKE0ZGywOQCusA
Y9yUZ3TFkVy6bWSGvvs5oe3yBuws/ukQ/e+AL3Rq2G+VSHvySfsxeDQ/C66n5xCNeMLI2folTM30
IPfvtulWGVXliGM2PCJ7q+ot4xHeAoeJGyj0kWj7/5EZrq2XTXa+JuP5FJf50HajcYbyXrKrq2YU
Ockptzsec5KP0uNby9Zd50LcelRzW2vRioxFm9Z85omE0Jzh8nSi6rbMplA8wKr0mLOIlbR8S1yj
r28BdHPm9ufYf49xymycnt8Db5Z+T7ugnlH/ClHvHVlED1Q4/r/PMQ8LzmEw1pZWjmfUgqosqubk
03c1FHLqXVgx2Dpejng/QMOWMxHLhcaWwZYQRrpnJ9Z280BBjVmqjr5iWEZ84UsUIoZBp7DdJMCz
O1x8PQJDLY/sadFsqCZ+dbKsvp8rJwEtJJFhkjdigLZoWBobR7+xmXYWCnZbl1rzy7ekovJQjzNp
hT3F9Q+yly6R1OEpZFzm8ZPVXYRWImo4sLExk9AitfL8zQ13KeWSan4LzQgtn7itBn676plEd2wf
LLBZlFTO3xvxRXZdwJfUMsRTErAdrDA3qIcIuukOLMOURpksnWj7TMBKkf9iXhcf3O4Yw1N1HiFw
PFO8XAMoZd1fVa40ulGwJ/2W5fKOuW0NokgAOlShAS5KEtgK6bV5iRvz8iHbuBDwDLgaEtS/f02V
hxeagWWntxv9ztt86Jz194xDhjsRiyGb7zg154uWm4MzD4uTjJMMiWiBy95wSDlB+N0qOJypOl1M
knmU+D8zJ4cEVqFH1ehORI28ta+Zttk3BqPsZeqSEcLW/3Np2BfqjrRfpo+cgT8nkdxM4zGpkhKY
6JV1TtY7VJD4JOxRWnZMKud/GChF+JpRjFi0fzSWjZjFb+xJGa+ENYcZajdfZwiLyxpQ8dAfAGgt
VbeqpDGSfDClsHpMgkMLR56zASoWrmkeNe2CGtxMoyZiyqUXOetD3eBnwwcHtSqeYjuCERuX0ikf
rNOpCbukwOVefMxrJrR2ERRsVu4uYk6UJP6cBYw7/4TTv0Wp+qZ1NTIk5to7H18S9JHxQxoL4zNx
0wiOvX3rRcofPsGmLBN1vETgaSJ27PUWOfak+AYRRc+LNFmyxseRz24hJWe0VAzdZv7zikrmg05X
jQ2CPAVSF17Xgh77aQPhICA+Ks9S9xAiPLNgCLWXFhfrD+CFGj8gWMXvwtXvzHX4ERcPi47qz/Wk
ByzyjSTHC7pJ1schqUmytVmUe6YbVPxt9J/7GJI+eW+zTUQaGDVSnIrGlf1ST0NK0tcPkYqXLmMA
Vzf8GgOXRSunFbpfti93MhhDxv+29vtLmNXze0DBciE22hoLczL3Fr+VJ5Nn4rGzR0ifgzu0Kfib
zp4DWWCS6dg+6SadCpCNyrFIJzvvO+JpSaFZH9X6Fhn2SvZud17E7EjXwQ+lmtukI0fspPLki7no
jW/cRVvVgOgBK9AyhghjxPJP4XlVtFcgVBrwo521KMQINAGwFjDLiZbFLVMTO45H3x3ETWc1SWj6
BbK+7C9rhXoHVMcB8C8TpbQdVzzFpX7eBnPyR0aMmzMsSDyoFbeDsARUuctPPb/ilAt88t3OfLDz
mTXlyMI1wsdGQEXijvHyJG6a3IAybRoGbX0nJ+w183k5qvkiZ/wsGHdBHzKFtwJd77xz+rKqRgGj
L0iAE+J8w71eGr365Gl8umEWBy23DvOGTlkTWiyUmwPLrYUY7m68We6tiyLS/jpigDmO2brt2CGJ
WmuRSdrzCN6ZK1hvSQ3pm6zFRzis4LhjXUFxqcS8Hra26KGXz3rYPiSPnjrjNPPRyIEXA7egpdRh
WgqvUyT9+4cc0isyGiDDjh0DbrLvJetML511q2e6GL0mjye0fzuXh9bTybYJhe8m5NDBdwFUYtXg
uB6Xvf+K1syq2b509cVph+UysTB/mEc55z0B7WDcGGhIoIs1RfaR/mGb/7GqkqWPajEEkbGBiVCI
y01sld/AFN1DDSlLj6tLnc09D548sEQOD6xJvxFjJarOAvCFeJInqMwV92SK1M7Icnme8WJ2aXxb
4SeiBHiOwrbdHHZSrSmXrhtS76GUffSfLcw4VHMH+1VzYzSETNZQqIZZCOuuzV/QkCN5pQ9Cy20U
gmz+i/tYGQkTvSMVhVsl22BDL9ufcnvzbT4FUqW3VusJcTMJgHjvXyBu1ca+XJhEmw4wIQfiokw9
tmf9Tm1kbmCubxBzh8foVbqlv7MWrYDEqDNpKl17u4IbndjCAGBKDZG5PvR7a0AwBZqVJxcCiL6u
WUfFxqW7rhxqknLBkBcdjBE94AyyV1cjlBW+hE/TgQ62QP+5MXGsunBfnVMEv1xg6kieT30x9xKJ
bSZlft0J0pO4CmDNpu888EiAiIIvAvzWI6SZ0xZxk2nCetBR9Jqi3+JLzdHuPJU+VrYMDrUx6/02
2WTeZrQbpC+2Notw0zqyCK2uxHUqNnR197q/BKLBO4GjUgDceumby42t/udz063/wzYr8UQ1PGLg
1hLQLqnBZ3ZXKUsjUQjg5I0hZsL+fNR7r8ZEX70PfIpbsYs1mYJWqxMeKBsWT2GHas4yzVE6YMrg
fl+TTmXU4yWiqR4l0KN6cR2SZj2SsHkQC9aZ5RSraX/jzAtOBhGOv/gczflUhDA8xPZS5lf+v51z
srYkTWxRXwmFZ0YtJ7Jemv1dq3GQa5eGL9wb9bjxFlAbnAS4G6Dad/QsSZb8i0tUuqBxCctOrPmn
KFNXLJokxDLfg0/331pvYTRCmvTGfS4IvNVnMvHWwwSxrUlZ7TOd5Sa9RIoxu+4cVIOIqst2Ww/h
XEqQywFi9GgnGRNslynbXEywwNyUxGHeUAg/CC5qw3ED9xavZmW9yGshGDFHP1DOzbCAFJTl6H4o
0qeMI225rNkwcx6xx5xZWmGIhMJ6v0qk+4HtMvEhO/pk03Bc9m03CDXDRBeeemg91uvvEvEwwKIa
yKAzArH7zxunfF1riOT13rW/QbDgRyUYQ0RsO5+k5A1pTJMB8wo1r2767+e4G+OXddK1ZQ6uImNN
CQ8gPgcT2n415tfzwQS00TnzgOW/BO4ZRMzBaUZ0JXZaGuupIUxkPD+vxFwbJNBytR3ETuljw8Yg
XXiJ5lTc/BP9L8NS1fBhFr358QuyWWrpfPsth/pI7vOheCng01OsuEx3FZTFQSd4ScARXSqEUWna
I8C/Dv0h8BAD8NTX4p5mWeKLeQWRmI8akMHbJ3kP6ci/cDpBReyZs1PxxR7xOA64ehzLoGzobK8A
wCg+RaV64GEn01iMI6OjOrrq7HADCjwSSCh1Pt03kXjN+DIq2/JONkg+d4G5WsJ5D8DASrK/BD63
3AuPYVVAu1Gr0jUIaHllk0iXfSbHvNFh2CUxK8XKxTkmgzMXdcTT3oJWg92XlR/5ZBcEHN8y4hbR
r1k189kxC2Stv998bpyx5TQ4sZnuInxOY/UvUs8dSNmfLBdJJXi3mJUDb2syZHFX/2OdpVF9Syb8
RP6p7mIAYLU2Sfa/PHkAFqLXXwnjw88Tiln8W9fTVp1oZx9soI57p3VqhaqE7fdRCtd3XbeDxyS9
KCBXbMB9o5InjQys4ADf58OdYqdF+CdzOr/ge2uuxpC42KEms5akW2J4/ESjYvtXZm1oIGSrjur9
V9GMqSfe2q9c4Qj2/ptRryuy3l20bAul9AFVHJghn2lBlym7Qrw3cufPsvugLyF/JdSaVSquWIli
fvNPp72Yq70oSR5YcTPfZg93sEeZeHRfAuKZUdqleHgkhm8fFsEn0E4Eb7qLnCfOj/25pRWj7WOt
GZO/D1rXd9h1ofplKw4PLAIvuwab1kv/Ruc7YtnndoUZZ2nJygSeQ9sKuD+quECFtRoxft/DCaWn
SreuUqJleV2t0a7u7k9IRMxMpfVPZ1NsUE8gJfN5hlvPh5DPRZcvM69ec5lxC6g5FaHFYjQMVYAT
Tdc10vSCk2ZIjWwaotAREG1iaB8wD622XDq/Nqa8/ksD88gQP94vhMO00AF07WqzuOTyGSh+fMiT
5AwtwXCPAKNuayePVM0dhRi0f/Zwsiqw0Yw6pcJWAWM73Z9rJ9awtc35S/k1gDdVEj9GRS1//uFK
5YekTbCB1bMIszC2c5tO0cjXwtu2BJmTpXFTWP4oqTvZh7MATsn+y/gJ0SsLjCEH52qxMhLqNEuS
C8Ho42y2/ihe1zayzI4u1A4qFexrKVmSeclcKd0H9fhZzxrzxMFLBqv7PQs8NAnb6tCOrHGZv6+r
fxMr17GN4EukWF+jUOLBUWnsUsb4S3d1qqS8723G8Ck75yCfgKg/Hn2Zyy68x+4iIyJynO8Pwf/0
jzg5jNJjBtcWlCS+yn/e/J7wpEUW2znSHji+1nOCqqkjkQVH2c9xV3sNSD+rVueFMbt5yXQYQiKC
AcYmqYkOM7GkySHpxXcgaOcdNoNnkqSxEdi9l9qb46E3US6h7AcKbN9RgBZ3yHjeuOjs4mbyvxYx
BjUjLOu6dFmw6y+GeB4YoXX0LpvNhId+5SpBS0ca2ButU4jWFKjviAbFjDOuc9545wdSmnPU9t5o
StFG5OJ3tv8ygCFVUPtstzx3LbsVT47MIw3qWhZfvvHcqVOaKefX9jD4xQLcjsYgJlzRJLeBZQMs
5O1p54wBC7Ozf5YlqmN/0Lv8ByzQ2nCRWSCy9WrINBWRaqAG1xU09nFW9KBJN36Slfqi9fecsiSj
M3jD0oUAa1LUcCQSYHdsjd5qs+IOjX1AoSYbXLSJMGCApObtRbzU2qdCa4ZeurOxDqdIXJhnUmXM
ewLuZFyZ0AI3MCZetGUwCkeWvBmvs5feRxsoBLQd2M0jVFOyorOEgH1pNMY548vPhIxffDnKu2mA
eMTkNXRJsdD3wgmEbINWjy46FL8+173fym0nMO0VMTJXOHmwwtMWWWmG3tcDdFmGcShZ1bbshvRK
gzRWDx9xRbV67D5shND74OyH6gs84w5plPPMXhqa4M9mHwPwW6WgVUNGTOG/kN3bzdCel87tWwtx
VtxOc4/vnnz3Ua5s6UZNq4LnTzn2sP8PEyg3hTq3ypEjitNePtrQoLxM/l4w0s02IabWVOPNhtak
1Ri3PRQ+R1Myl3h1kC9yOElgPgCDXmD6/MzjUqQUM89s9PezkEM2Etx3YGf6Z9Lh6K1L57HAEoKY
4nXlLn4TM4LukXUnoQZSkdS96/u9t4IRQJtXBU9/aQ1gMTp9bbfkSAyJ6my6i7KkMlFPB27wVmMg
3GMee4dSGJ0gcALLzKMw+ZTD1wf5YD+Po9DIPXMPNtAPo3aSX6GOJeAgAZlysayzoqPlVmP1YMZM
cH09O/PjEVA7oIPsv7bfVelsx3tWbbxXh7o9olVhedqXu4X2yY0Wrx+j2F5wI+Xr+LsvWJnKNqq0
TWptdfPXw8bucGvxsuWqbCQiOAOQhTzd3cnpkl4k9Seo50693wNQJwa8ahHwE1ZD4yXP8s+RW0zk
Usby3vbIWRrKKwHwtaYRHuPjG800+Xrb6K/DfWqoRjnO2o1TNCh9gyG/wKmfhyi7FL6fzei97KNl
KD9tt6mABy/rNunN/d9sXGpk7k1/62x03ELdLgdSPszp9jUGTMc/4oG5Vn8obQ1/sQq6I2IK0opy
iAKbXAVQv6JboJnGa0FkrMVXwtaN0qQ8owyH5qwO5yvfkrfywsyQCJl4h1xK6CMki4zFe1knNITS
56r0icKDIh0B64tnv3GSH43+tBIJ6QPiHVWPEORAEW139cURJ3DLXikpJhrhkLkyVuSUqzdbRdBR
7VyHTOHM0x+EQ3yH9R5kZiAdoVmE29tyC6bRlUQkBNpfD7qB/Kj/hBT+CV3utfM3xkn8WX7I3v/X
xLUb2dAj2zTLcuo6DOFe0DjgX4CXo4gPRjVW3jqqHC2rtqcuinjG8Og5Xp/OTPa9QVZuP/NuHDR7
yUoRD4Ph8pr23sL5dgrHBa4ouF1ccxkoOO/+EtqqeCngKbtOErcS7WPJhNEtucZkH+KNZECuQeMB
Zd+dzQdJd4isJzhFca1SDR+u8VWRLIw43SgStBIEdj+eVUtNaXCexfkJ/C4VVU6JbMkDPMb+PqBj
4UGG/cPchNvXUdUr9YuMAgf70f277WmA5cIzTxy0cPXEe8ifOP2DajMQXvIBpM0dRyq1A9EU7Mm7
y8YDt2hmup/n/ihG1gUr+5hw/5JvH+zJ8eU8tqb/fOXiELjLox15Ezy1zupxSCkAyRZWf0nmc5Hk
kY8YKlq5mth4OlWP3GuZY0/6MNbmgQOKQ73HpSY35mnQwOFn09BUbkqRho1XIfXXyZlstK/hcp3U
UJxHw5NKjaq3LP/2Bo0FRPF43nPUoMs22zT91KY3yTVxO5PmRCQTwJP12Cu+P0Ncefxn8XySMj/s
mxQTrmGQx2J8JaBacRlvsrUhJpoufVd/hPItndRxgr88G3/ZB399EJCkvhdyW0/i62TvBeqiItb/
/WESrbcdX7+SNU2ezBoETTMg0Xlc46R/9+MvP0UiogEjQvN71GPPwmH5YfAxhBGVKCsMS6ApFNBO
gMr+8Y3wqG+Ll3oLjRGsia0Q5E6bMR3KcJpBsTYkeKaTty6H0ZAI0ATWs73vxUxlawS8F8WrXls8
9sWidAu0bktvI7E3xTyRz5uVyKmNRdwDULoY7nIit6r8yEkEcxJe84yxvuYjadDKhNVqBfRGtiwH
wVwkzcCD5xwTSGjFvauLGl4t66w/DDXV+5u3gY3N3eZsMiTH1hTPS2tQNs7VfslEZcqmrbxWmaDK
a1ctBK/0bFlMITFpY2+xVO2gAZO/7rJipIxQCSRyLA9vwbtmX7Ig5JJd6MVNGVYSHUp076jSlYUx
a/peQOyCYdEqZ0GZum9728duFyW1+L242S0s1djFkxOcca+wQgzfZAgZiRrMHAOSQuRfntXK3Nyl
SIdfKsEToR+2BQ/D56+s/zLXBZhTtbJgj/RiBHsTaIQYDb3F2h/7kUJ1VdACxBfyFn0FUu7OXx0a
phfMzy2DM32zoa9QuI7f8D7LTdXu/jRdBff25nP+Ihx7KtIIab7GZgrvGicbAsE/UA19BXwHec4r
5Sf8YiLt6F0wKSKqgMI37ouDOhBTMcsRbGz/gSqJ4v6lhMLqKAnIW+Qstq2q16DUdzdH/QcsY0Zh
xIKifHqOzOz2Vu7ez/mq6eolErz/D34sYFSNGfNvWmmCJKuJahxul2D44SYCy2oY11XS+bj2a6DO
NJtrCxnc4A7w928RtXLKoxy8KXKsUrYl0KVbc9Q/IYOMm0pXisW/6yABH/lydF8//HPrbonGyIlS
YhiBpMNRtRkTuqNs0peKKKxo23oANwok3YI2jqB63gTX5Yz5hCXDtgO/s7qxVAdENDDMEbyy9DNi
jYxdfSF6C1o0bfzr9wV4tAFQtps7XqqmBMIceYfsrjiC9ZBB63he3f1+PL+wCLtHCd69vWvnT+JK
sjhChbDMUjzlm58HFVbzhjTuu/unNiQOfLYgGBgJN9V5wmUIvZOQ2ipiwa8IVEpSekJx7FoM3908
EXmlDVNfwq1VPAANoUD/GSGZD77Fd+s4frHjw932iCKmk534SI+jLzikQujJGfigsfXbNZ+vt37B
F8dFGe9afUWa/JTfGkTJzyZjM1rFaZZI8tAV/bT5jLLIPXIObTxm4R9hIJRZKCrSD8iDIihGlLCv
mMBNx9IfygaGBLvUqpdm8mYadVGZiPPa5+yYqPT3oCLd3ouYHx+H7tRnZvIzXbAoHxS4lGG4tvm8
YdfOWJ9fp4eA+q7QqZyHkn+B3EW67v5O91yiOL71qVj3ZIUJ6YaXbBTziuWAg0CO9FY402rjgIaC
29UMn/2fdlPaL3oDEMNL091Ukrn1cF/twm5c9SifLJv93WgZ6Lzz++W/j9hIGT2qrbB7yo0UaeW/
QbIefFSZRuixjbP1j0PO00ZqxbIQaYXJ/BSPWqnibXDxv6qyijPUIOwI0BOnQTu7CEgsX69aFejv
/dY56p/O0r9gH/ctKifrZPS4y/SzhLrYiiiXgU3SSempdagOFI/1GLhfAGVPRPxaj7gVaGiBOVGE
vr98V9cWHY+zA82sORjIFWXFK9FG5G/N+WKt8Ov/7sVFyUtmWj1Dz6xv3JQJ7EJH1NOWw5tQzftS
w/3RRcQgCuC72LDCwepEQ4rCwzGw3CajF08gA9DUza8OYkgQjYhp8+u9/NOyvCjBrk4dv+pxEeSe
ggP8xq9dIcTVAWF1ElypC6cF/mC/+U6wcFjcBU3LNV1wZ/JawG4jpUqnSmig+xYT5MLOqkfhgin3
U+pVW8WqogxfKmY0Z4Get4dasNaPRnmIeDxlWrVpIGJbyjG942Zlm456E8W0y2AIINPwu4LsNB+5
HUGUZn9b/51hX6/lHh7zr2sCn1863BHMcTaBf7ROs7m4vvv0o+ds6rLKStvNDTffwCdjEZUaLAqp
LzzealOSlubro51VQyNXCJ7om7wZNYRB5ZzBKIjPcG2iFJMbTd3k4jAdgq7Fq23gdMlvp2K3QdRy
WcWhoiadEBEZ4aUOUd7CnZmLkUxIs57iAbbC2A4WcCkUNvO31jO8o9dn96qAR+RbP5/tiutFq6UB
TvIQvhYkPPLUBxPcr+lTzwXEQvRe3m+M9IPpW7yOVY5X3LxEzlgObIRkOSR9+Fds6N3ha3dBZ7fh
mJ2TwNPcSZ3i1iI1gDBChAqyr6PGu8/RAdBUnUWyQaX6lTg/Inu6T9civy4AfuN9k332i3clL3U2
Adnvr4NZ7OAyOktasA1zX2PiwOQRaowlu6IVODluV7PQTqD3MnmrmjP8iyeH8guJ2yd/rv2Y6IJX
Kl8kYZsDC2OmgVHlKpL4HF3aqlLxfXGmFAIPkkG2cKQ56n+D/QmmIXuTapF5czSjPgDZIAvnRjKS
IEr9YtZHBv6t3MjP80/a1iP/UFY8K9oQp2SUREU65DyKbBS7Mu0l/a8S++4Qcx5bpJSaeJwsmamB
YlnOKmtvXue2AYJh1OS6+Fp2LyCLnGosywVLXNzv6A6lRBZnj4w+ZgJ15XGFDZPfFVOlQwOPUgub
2LgWm9YB4rX7Al5myl68NqEHfeWZp1PSM+EXcilSXCqxLEtKohFmWxnsfD+FRJbNjBNozEqa8HnO
WcYRkEvpbjpJ98IY90V6F2aDdppBRtNWb4qbwtS9OHIHtc2bb4iXgUgBxcua2eFzyRpr+zWUbSAb
pYWT0ffZiURGxLiYYdRlW8fKEHOhy32I320WPJPbCEHS/9gkn4wSQS+4d5knEOeyb6JJkzkjRAxT
9CFSUSCaM4SVIWSLsxVnsQz41JMj4eAR4sRF7BcWI1exVkGsNNPXLd+IDc1RNgH0Xq/5ZiHM0Ug3
f6eOXHs60+Q1y9Rw4HyJdB3qmpUdRjxUrEuBNJWu8hGkWSHLmj+9ujtiWhFDVEnZWU7wC2kCofb6
JJms13Pk9+F6cRrhfITNfMARSugZgIknrqV4aXzNuFU4FlVJ9TVIkZHybNfVuDzDOs44wvQBvsKg
RfdK7YXtwVvvHfQif7PFB41mR+7uDtxgfxCANrOvGqDVCHh8mmSCJat23nSgMfl+47bTGmZxRw4q
qG1fhFpBkYv8UOyG0fA2J5fYozmOBI3b9bRZFUgivWzwfwitkFGBb3DvgMFHUo8t9HezHW5g3hOv
MgdahpKNViS2MfyIyMIkDhzvw7feztRLKG74NIvUPxxDizh4q3tuKRAZRzGX3jfjehPMll4i04Tk
oNoT7KeVH9dJ04QJj9Xw0Ff/BM8PD5TBBL/pzkbeZDkM4oEkbr/M8Tc4Ij69QXPcDaIf2mkFseFK
S0PtP6ajL2hHNGI+/uid3V/rgVvNF0pbCv6T+dNDKNiv42uZFXJUEwE7ig5Jw7GlHBFZb2P7cTIx
PAS1JvhEz3pXHfCrSBGEN3q9fKjb1vBXGJSN+lyvaZgywd8a+1/tURRPS/iNaHhVy+8fEUmfPBP4
PjyoyK0a+hlM98MBWhIedjPHXvuEcZFDr+iE7eWnbDMgmmfm3J8KaVHSFkLxBQzR9eBdwnsAs9a0
/1ueafK3SZIzx+7ZawCNb6G5M5hjFMuU/CqvF0+EatvQiM05DVn/m5Wx+/ELFzMamRZJzL/FycSf
owTH8rRxAs1dzfWvkbahGaILAPr7AGJXCTVUZoiFrvC7EVZryyPYTJQwsgGpEE7U9RmPla1FPqyJ
Wy9oN0VKMRYpId9ul4ztlKGhZC50fJNGCc2k9ts907G4qb8hG4rk/HKSvmgRoCgDoWEEE1YXU5EC
ogoRNSuUbd+pUiZhvIKsGLDH9EDxLQfohfnzadYJj8suRkc847Wb/RWsKJjUTqweYF+5s9tTiNRt
lA7ZqGrBh47kU5RMx8sT2JRw6ioZlyoycG9BD7HgnPxH/99k5GFAeMglNNyUpkhFmCRbAD7yp8UZ
qFc7in0d51XlgMU6DnUYHnHQxvLpR34cBOtyP3MV6jz7SiWxAx7Wy76py2Q8uhEW3Hc207wFByT0
uZ2YB2HHeu7AH/F87b5Hse3TbsQQ1Jb603gt+35WJLX/24kr20YaBsSABiRsH41+rnkTcx0kktrk
IBc7d22HEG3zgg8HFTzaGXB0+quVWtkQ9+ubUig7dFdpTY+E556w3faYJ1MCnwXqagJDfuHcsRqf
cVhgfBvDAoN3dCjQMYoQswyy2Nt4LYLj6i1VfRIRR4U9riQbiQ4Xmd9y3v0/5YBHHmIVSZr1Oj/F
fLPnK0gzl+DNpO6NyVghK3eCD19ixk2WeXmQ2oBIuGNrzTXIkGQ6GxU6zzmxAuHyrj3R3EfAwLbL
xHKS8/eVWhkCiAxwspawj80LVVUlZVv2cRTMNIhL/pUBJdA5BKoUo3q0Y4WjfWbll33GCObeYtDI
NBiZyjHR6qglnOXnC5OsvaCT5gYZ0z/O3yCX8YTcpdPlzOOwodN9edSjIoQGmZUMKeAy9yFmLHkt
FnCDegjD1d39wxx4OGS2yJy6+CcEx9ejRNMmovRvk03DjgUngpqByTNcqjQs9/ZHjnW5dbKupG0Y
2wHgDejrwSFC7eLUWA8mpjnYAPMZILT2Bv8y9p4IG76rl8hIZydRyzvZkpB7rAtUPY5CPImx9VQE
gIRr0R4kBnKKPFEEod9HR0fUgYB6vWYcFhF5geLy5qFJOHjU0WV1AzqpwWhC+gcVUQhLa26W3bYn
GFTtlkkwLHhbqYzIr+H5KyK0KH8GoM0QAhscfnqhGge9wDS5AfIhg9wb3qGUXIyTtlDJT2WMfJKe
fBoKK9kSktldlqXggtVsAB7R//3gDpMkUvzXfsTNGuI/5xd2e3fgOUXt3tuDiHA4Soxc8yL89CpN
r/KBNPuQIfXbXYfyQDKyS50VGS29MiasdbV4mK490Vm1tvafkoN6Oeb6s0eE1K0gs9xEVDhrSeLH
aq76ui7R76u6cnYR53WPKxX3GrzyjR2NyaffidX1e8Et/XzIzmLgN4I+m6rlgzLO8h+xEqD7WhVv
5E7RmprLCCIrgyy6fE7kSaUtvS2bdaZ3sBT3KIxfhnsKlQn29Bl982f0n1PqUQu7iDj7TFFWWGWR
mcc2SPqX/IqYHyoWloxNXIENq29Ym/RAgAa8pLENG9/Gj90+f+UgNganmC62Y+oki8TGyoT8iabK
lgGFklBw+05hHZM48cHd1yzJ94aKEadPFpgH+W3Sd4mMuDW3ADgWVDo/aOh9v6IYHPZmeZrdKGE5
OC56v9nepRGczGrSZM+sZLBoE2oi/C/p6zUrZYVer83dyHwoC7UKvJIRexTXNWe/I59Y+NLmiwiF
kXYAzhOhJdLFbUm3o6Kv4jvFs2Zn/W9DYhvKo1HbSAbEV2exiEt3d6e9th1qwjirJ3P7U/on8pSn
3siJFpIcmFhOXMO+zdTZYlJ+EDAlJJ714iJSX33tQsP1zDvefUINYv7a70nrojxWc0Cmz60Nxczm
90elmUnVpJdokOEE/xJAhmvMND76WEweBPY40xvDFzp8zGhzO3/au+CZMMQyc3HpfxqNitQDyfyF
NWEZmft8/rNHBIdyykXnlcxfsw3wGFlsvsny8juqP4ck+QFV7SqF+ZQa2lQOQQWeWiAGSCX4A06i
mFUKbf9k47NCAgyB6eRxsSqVB5wGv8oH4lhzo6sdKLty1QRa+gxuelHtQp/7mlbZZMw/SuAS6JLj
DmpOaOXZ/pqsl0JHyJLQkz0ihAumaXFDOVKCJIAFpS6j5pDK3Rs7z0liLnV80OUySqVKHEJn0AEA
YptCuQSDC54LyqLYcb4ZNjZIiQoe52xNlLLKddZT6IwXzvoL2DUmLpfVlMidzHEVzWl89Cc1PuUC
hpaH10LLiGdzekpDNROTbWezT94kT7Suk02qrhoARsOi1XmbV6YQWvSnhd9n0TmLB1rglCTEGlzU
e8Ul8BIhimRm7TyQrGuDYLJGfQYxwAwJtXXyMwE9SD62FH/uhDX0Wm2pANim+6bsuvHwEmJDchth
oXU4dH3XoTkdprJGct24Njduj3m+Wqoi2rfLCp4dhjp/J/ziJ+PnDEVmIUNKPIpjFXpZkwkhS1nu
6+5dvZWtGKZHdqIRgkIQcdKf1Mcd9ISRnrXM8EdqWloB1gBffdYuioy4ZKDBhJPmlNOxkNK7Dv4K
OuiPx5baMwezc6Hk9Txrz2OtVgOSP6teebwAI0bQHIYpCTLc8mSq8gRaeflFXEG21UZU8wkQe/3L
9y0kusoLyIOF0fPnbrPqJ3k/87zpQFvH+soQ3anS6zpzFE3QL8Fzn3zWCFeR8IjPOuQtdFEdYDvl
nBotHanm0VfMYvRWdVc5FQZSTpcV5SCXr8P3T1cAngqi45XqABfP3WFk60YKqjVjm080b7PhynKC
tFmYVOSYiE5R5KOQTPNQaDjF593H+6dqT6C7QyzqP7/P5nfL1KxRsnWZ0ltry9N2NUfrUQoODYxa
bDRmlZfoSebM5biX7k8Kfnxk9Oa0sfMPZLMV14M2d1F2hnOOQlHBZ1vo4GkFXA4zQSWiB6vykwY+
2nmwY5F1hLjzx1fo71GVJ6+rRlwRloCH9IelOYModFV5MIh3pzmWNrtqvS7/JLKpFK8b3PyhIF0d
jwXUeOkEIg7pmdwHMSL1fpCKXzGXJBD+yGt+z0QXMtGLP3pYv+EvqldbW0I2tF3hrG4if9ejbsF2
VTbiOgcMhdTKQKGU8yU95JR991YwBqSOf5ggUojSJbpN11KILtk0RtjM4odR/I2dVS1cHn7FFx0a
eN1+1nSTI2CKjZ2RrHY8IkSvaqnIdUA7Ec7/XC2y5FlSFutfq9aTxfVQxbXRePDQlo4cejSvRbqu
VqEIi8FycuDZ+66cKkrnOXrQWECQujQA2DCnU4VuydrQ/3XYLSYbQeiAdHUGpnOOLyD0zWhtw77k
8zpSBpEjdLObdcm9aHZHvCenmqYJeXYpixzqGxgSphf+T9UkYiMr7Mo91hdybK1FMqj57OHu9Wje
kqDjrWe/QxbC3cwmeKeSoEuo0g5Vt+dodC3zYMIzHi81SSZbZ07x3VBEMgQpCptiidOjE0O39FBd
FiszP6cEzTA3J14iQI4Mw8/zw1ggyrbjDa4jGL2arBt/Fp/eVcvuoh/LzPBLJcy17vFJXuqlBEEB
7s8DAoxZeZ9lDirouTFSJwatkVNe3Tx3wmn30JDHMsxwrX0GWMdklGRY5ZrtPvERX7a/CWCQcXdh
yRDs5GCskn1D+5Q8K6XC1lDHGo2fdFG8nLnyLA2LQgiYJfnGa2yNIErBxRT7+14z0s7mVO8wPERF
z0lzfftg3cqWgKZBWBp/PhIF3jhuQ1vBuxiw5KnPBPfkphGkm42aXdgEXUxfU7LuTZg1R2VwVW1t
nYbzPb6BdQVC8xoAP1DL0dfGJK7KDlFKjoJld7+MK1n193C/pXmiJ+dwGGNNSY4Z2g44PPSwnUMe
uEeAdyWCy5yRix7Bn4Cv7tD8S8/Kz2mw5Kvu25lY98e0A4AXfLZnL+H9aHLBEI2yjzL4Mvj4mzTc
O41b7lghjpZBk1kuYzpb5bglIn2LcsyIvt1H2FsQoW6rc+x+Nf3bhGrk82OwxvR/LY9VSqH77DUn
4wKahXYPBKlfr1JgYwOmdOQCyn/OByUSJGzBSDG8V7TzRuQMCvwuzBc5ZPXW7LlTL63PDs1M3hLA
xgyDfLfUkV4tu/TevTS4pJ3bfRVH0H7KAtAWxNiVQxXUJJs9lQTiW6/FExBBnWWcmpiyc46nYGiU
n5SaN+dGzAACbxqpynZ2gRdq60CL86PfewXtQnYIY+fpvz06q2/nzRYMQQWZYTbI+4F1EaiZMqQL
HuN0f6oL8+O46RszXVQA8Om5dLgCy2qoQ4B6DjhoguhezstzbcQcHHlGpRY1mvwIT9UQ5o4en1RZ
9PIr5VGaFiIcbpWyo+pf1Ht6WNRACsDwNoN6NZuPkC1tDYkdrX18j7cyz1tnoq6v2gyWpFBM2WuU
2t3Ucps7Ntl+XMNbGPAQ3slh0SdCeHzx6qsnCQ9Iqfo+3tyDkSKWIky5UuJA/dFdep5+BNWFsvvd
nG/nuCg1ZVVNKzzFtA5+J/qV5whezz6yGhZBAdwDz1ga7ZGZIGhzxdD5sySCwqFw2fcnBVsgL0zA
26MehLKaLwGMiC9EqNfzJ5yiCQSszn3Vg+DsnXead6OAdY8fSy53C02AG4veck6EEyx38CGe1VU0
KJK/jlIuq0rGGuLpTg6+w65qBZalwqOccCJSRzfOVfLxZyNpSUh6xHvT4ibB5i/8yp1xvKrBxtGS
akJafqLtO7j1u3JOxnZqXCXwU9UYVxZzG/d4cBDsQZyrDv2Z0WRM2gNET8t40ZMzUbzN69wZ2FSs
Y3H2NjaYLHLRNM8xr91um9tJokuzL67LE+9sCtgWlxPOcOxHn0shKMK9Pj8jM0IHBoC9WKZgBOkB
EOCcIGFF+vYaRCgV/f/v+XA8C0cVZmEjn9QfNDscjLoh+IMcSQBzqTYrR4WeaQZ4R59gjBmsQ3hY
mBeiCmKP4dVdyRLvedKzdnZueE1s+DJDRtX5t7qh5Tw7pwexqTxnBq4fRGYDDSrikjdvuH1jMuEF
ADaIb6XRaSsWZDs2mknMW/RE0VzuG5eO8r847OmyeIwXV7ZGZzGjkQ+fzSDgB5EUlz/ASi6NKOLl
6DtuG4aQlJHvNA4kcQSqHu0R2Piy4UBIQ+IFxYq1z7u/6a4hq7vbnXneMTd9k6cFHLrbhMljEgdG
IPIFtlYjKH2fX+3rKbtuSGLcc9x6/kOypFleqJUiSifTCv9G2hKzhn/43o4VLRHCY9tUuOuEJxRT
DPTCwr6cRiomdEP1qDTO5aM4TxOC5181wiD3OPgQ9ZzRKOhrWUYOzfFbWm3H+S6fuCIICxVLnQjt
8AVF8JrU4TbtoV0Tj2/diyCErn/TL1xMp0eImycmEOOIGEnJmGYTVYWbjenuCO+A9H0YJrdbp8Ib
e5aXmvkD8r12R8YO5R454FH6ndTpnqwTKUMNicdnQBdPWv5uX9q8661BxKWiJzqYqex7ax72X6/G
CdnCzzK5fcPbBn7LFrwnx4rE+irX7NBLmVvm6bN3Stzbo430A23O7WrOP2RUTL7dFaLB+0MTjrWa
FSSrZiyOVl7O4ea9qdVUUWw2gdNS1CiTosfcytQxU12JbC+Nnr7wn/tWWrX1MNMekV9OZ+3ngZ8A
2PI2nCEwl6IbumuacARxUSoerlsWffbWigp5iebRU8HEu44lJWx58D/6DydQmjFDpqUsghjmCwC+
zCGO3GXdyNNAJVKuA0eDlyXUJh9JwrPLXTB8cv4nwyGNukQf/wRidNJ4A0hhrOJbVok/c1DFzR3c
2e4aUKXqdEI+bPoIMOYNcWVL2fPyHl7iMR3W8RtByFq5rhiceyjKnhsgn3Zicm/Qz7qN9QHcHGur
LDI8KVngFFs2PmXOpeyiCWnimQ3tgtyvDBEWfWzyPHk9VoNNvZSBoKVSAni7NTIn0tOrv14FP/ge
R3s+MQHsy5Swx1Nr2Utch+UQar8j+OgK6iyk/Vhb5g+WP+QpNjhDNMyyoqt2kK2ce5F6j06Cbt/p
R660wqdszl9howo90ipqwq2zIL+68j+W/1QRRuqNQW5m2iGIdSYc7588sxws6RSD9u870LO1zLi3
B8kSl/zE2Xs2j5eUKRtO6me23dgUJ2B6hRzh0hBz8rJjUV2HQEDbvAi/TcIp9yEH7ipnx6xVZVeA
rm+15cjvSP1ddYjPLICMDrnznyDNICfe0HI0EubZ/+VHvtzRwEEvONWtYWauHfa1hbo6uo3LJ24z
LYras/0ZDu0qeW4CYNbSnB6/EH07lwrAR76CtCISjECG2QFi59kvUmizQ+hQjod27TOtJKB1bEli
akeDeUzItzj8Jeshu6aew9ZOJ9/1uaWuUUoqj3UrIl8wbJ+gATIEtRWYjty4CmftfWCGvbTe385j
uWjTTmN2lxXSUYx2M5CrBsva405VilAYbsvcNhQNd+m3qjM6PO+Uzbg6CXJIjCo93pH/kxF0NGDV
ihZmMD80qkm7uNexZM6JtLq97YO7zTWdmRsMRRSJiQON4ytF9Nx5eAU3vxEvcT3V+VWMUZgUzSTl
bt3KmxvP4O3lHQK9S9hX/Gc+12ilibTEn8TTEgGP6Sx0jC+usDDUAQeHVzjUC1nf5aPLKAZ9RD8Z
dO1OIMen+rx7uY+FUUZKtlvOCePLhlUaM5wZbXuh4UMryT3CL4jEcb+RZMURdwvfY0UeVcDWK9Ez
7Wtc3XwbESKB6m2Dglx+EB+RJId2lrNnbVwJ8mwddgtP3u9uv8/xUOakHtFTD86IEu+zIT4FZb67
9ckO1vHjsFbnE4maXuGxxkHtkSfj/4bZmunAQsDFc9KymW4fnsIg65lB/suRFd61POzEfx/k6Vwj
CgMRSKFUFzSdOYLCEn7k6EXUbavrA2d2S+J/0lFZ3YkWorwgqnPi1ohXUCfu3yT29vORhqcdW8v2
ZEddxD1u8NBrxavQAIUoPAwzZEz2qR3//bwMV4Ox1Hdh3FUK8xx9JR3wLgbo8UYvuA2jIlOOI1p6
DwOYzOAS/i5/WtY01RAYZrSdR3JToPcB6hSBCohGm0MjEatYAN/m/xHQoo2rerxgIqQDWsKfactr
d8QzkxNDCQ4VkAe1MP7pOK4dwLneXzKO/fgyFLNVTOxVkFjW79YqAzSuW+uHBVeUCB6syTgTy6bt
SeN/arZXIpWucR8kE07uMcxUy1TlXrHP1hBXMz5zYKxMtybr1526Nt/7uEydMn6pd0Od++PRJNlR
juDlVSgJw74TuK8TG+Tc73sbfkd2WG7h86qm9GFH/ee/lXIbF8aj2jpx9cYGH2vuDIEwvspbsYdM
hfya5VP41r+QqhdvyU1Z3+VcWif3PcTf305yBSIU7nBIgnPy/2jNaH4OcTut+PomvBZd+4t3OKM+
wJWHcw8eepF5nNJWjn86Q4ogTqIK3GQ49fiOhkn0NsAQ9u86w/sVNlrnH8GTwg4YXoyOSp/cPQA+
dhrFLfPuK4fFQarGT371lBnZhcdGiXfFP8g0VzJZsDtJ+sRvfjY3nOBxLq1vmqzNDKA3TZw8K6Kq
otqburwCiQ3tEce0fQhgy3uBKxokyMJaWYakaHPbt1vC4yZQg+cXM2K/Xt0TEk1eisxleiwcDcaR
piplu97MKa9Sg2FLlnsCggaSsjrJX5gk/IptWjrCNmmDySVH3TWZCs3/yoJEmrgkr+mgzMHwMRYP
2RHN3x5oToUFKUVjtKz0SmGg9OrUBIvA7ngjt4woiQFOuKuPUIOe++vsFvc1Nk60K8eSzYuwSW29
26nsUxcGnF09Y8mqKfHv3ox7Ai+hAhwi1d92CI5EM8o6vflblL+dxPCLEv8v1TnYjpUCrEgyZgGP
jAhLvU6iTX3LiEUwST68OuMRUX+r/ULblW6MHvkcm+JdNrsNiAsFGWzkruKIP0CoCP3uoSlqvqap
fKcvg4BLZ64UcxPAsiAzTsu5xDdRnxiOEagHgKs4rz45V17WIh7cCdF5y2d91loz0vYG+ePEt7mC
uKOSpsa5SnjuX/UbY6eY0Mq9rTLuQ1ddEj0YZJ/ThVn9jc2yzwcb+5KcqQ683acNfubgH9jZ6gku
57FFFMWHuwR/38FCO1F3F0FsGjNcz+9Q7tqiEIHSiWK/aKmIUTC1yDkCHVx53jZHOlslgvWyA4dy
BEfijbmHwre1k2TeqetVqzrOF0FKxmnks3F342q3q/dyq+BO+Qh9y+XNAXrxU3F+OQzaSUxwNChP
yyFVnUiI7F4YTzogEt+827jrpRyvGqGYY6CYKysKNdJHdJ6GPBL2ypUO1Q/a422CROFBxNKAngJh
x9nZXzqTteDQiJGZ01u/kePsKNX3DSC2nuUopJuL1O3lSbxex4whEYp+pLgcZVHvhjt3CvGD86vz
u8zKHJ/pNh3vNAptjCOGAkGlRansaLVTQ0qJ2mzHh6hfeKmV7r4yT9SVnQJQ0ZcdZPuSE/ERtzf9
SmefeCFCEZiNgEJus2uxDDeZoDpKe75MR3A8vq9i2+TiZmJkM1VF3FmGiOG5Mou5AEmheQT5Qv/a
yifdOThegzl8SD0seRycl0t5Nijj7aBz+DJrv76N2SJ/FvdmJb30yODeUYZPCQVzjZabIxG0RzfB
mROKszeLUirwBasKp4+BIQ3Pfio7wetzfs3q17BM68DxDI04v+pH3qKk/y8ngA7Z7yrxigy50CYz
qVD8+o8RC7knqYTlV9dx1PYzVQO9PY8XSbHzhKU+Poa/HA2sU9lh25Su8fvHQoPLf8/9znQMKM8o
kH4wFJP7QgUBA5l6krdK0JcxDBRKLnm3oQTlLi/PO5NnF6oEW3R/qV/u0at+8+z3283968dUPe4n
9sU1owQiKBKBW68vDladAR4L+w566SqP9lRwhKQ46RrGRuJW960+R24J22fA1Ga2r1X9Yn80nDnU
f0Ep/C5YdppqJ+qtLg9GWpmLuzfyPwvvYHSEsfCejO4LMb84MKi3VBVIQcnf9TOUfsLNyDpDQTi1
RukBgCPvxvN3QdikWUp7Y/rphvOJL7QOi/M/RhZk47jkADOlmRBk16nIWVTjHfGRS1sqJLwi2cmX
hBWlL+3OUbIPRy2+GTVRKjxX61huFKjoYDM9n9eN7CDc1beU8k7VqPm39NvtG/Ptz6joQyuum4nE
imJEh+nySZH1SkKJSmJMgCqlBnUagL5vkQXI+KEC1Le3PAUyLdQFJUhjoUQlBPJPsa0v7Z6THWXG
8LTWr/ciwBTu+M0XM1m+laj10AkCiDph1Jq+SH9Vk1OIGOhGDemvn6Di0Lzk4O9tNKMbNndKvtW1
KNSCIS3VAJ3RTYtS4Ll2AxZJepc8TqdhtXKueld22TO3PqgYe3wpVgAEqciwv0TnDMSx4tx46+3V
V5AKpF3F/KY0RLwQNZjXtBnIoNMVXyY9kO84/dQ5hw3LG7WI2x6RbLNFTmeIvYkWTk6o7DVklOFd
mxxwv7XJKfRQs6WxUs+Hr5RoAzzlQvT7rgOpxkh118adJflApJICxPQyQPFSU1tYHLd+nkxNVAG0
o5H/a8OWnV1dB/JLoGSPLX9YO5i+djEdoNO8YIrBldYQmdO8bnfJ4QnOPALIbMa7FNLcKGUzEfC5
NR6bm6gbOO018baBoz9bbKaO2DP3NQpPo3PQb2bwklxd6lV2Gxt697CMA8yGZZ6moa2FAyQFoHyW
Ke0T/XuA7TNoy2g0zS9lnQsRP4b8ckT/1OOCgwwEJwx+mXfhtoerijMMTx7u9pTVBzW8f0rd4clQ
Q62TdanoAjpESh/AvbsUlwg08iGdDSvVrt8uTMc5Zknho5gufXzvXpgYOB4PYuXRCchdZiQMciwD
f3CTPJ57xlhsTJAYX5rQtx7YqQy7POZShgJPOtM1NKbWKJ0fh0owrPPsBZX/c13FJVHHv17rZRRc
Kxa0htQC4AMxpKzM2Cm7Hz/taaV3bfEsymo37vc8zIzGNxEUXXPYi6vO4ugEpqxNCkODiUo6m6c4
FX3SwE1Vxqtsce3YWIPHFMvJBu2k3wd2cKY8+SbXFNJaB4lkFBsXJgkFLgdKm6jxq0yT6IWWBsQX
s4me7QdLXJGEn98fLqVCC6yNx2/LBmcTZq/3A5w4rtVlBxXD63LdvK0Tj4KSifzIS6oRm8QZp8tP
OyvQK+3C/RYK+341HK4jIakb+VmyHTI6OrG40gWaw5A0TAXjIjZpbzoeuTYvzHecOvwZuTR6s45U
KCwP3eseRinhCmKdzJz1xO6LNCQc6YNY6F0O5ZZF1JlNLMwBOyaZZZj40jOyMNC3LaS+8+l4ML91
yoBFYgCg2UBx80aVNVl5YCDBxrD1Lm8fX9CmFhXOubgi1rTtKKI9ImgXctsB4kaaAGGN5bM5psBX
vEb3m3Q0QQ6Zi34B6LVpMEffNW4dFNrWFfXddqRx6OcHHX2HPTPFE7tajIRrdRQv14YtoRt5cjgA
kaOLmDZIZI0a+xNBzG1S+W3BSaTerpW1AJJjEQho+qhRgQTQd739oCOsYLIYuV1bXg0m30vJjaeK
ZNAVf7I9ezB02H1i/7njt0G0IWyItMTTyRqJl3vLMfyKykZ0QgmMc3VNLp3yfZNbL8Sv0HEwDIk3
Blj5l+wjmz7lIc2KANhATGs5PJiJ8j/JQzoIXgB4NemvW9wK8r3e/rkzWACYxWwg5a4oEOKwyt7U
qJGsVUMjKnk6CtSjbmFFTG34iTfnmQ8AvpHsSdlhtHpOHNQWy1efaNGGD89Nky9tVEgTyDMzU+Iu
er1IxMi/RSG2MuzQen3FFf+0M8HqArygzRrBD418cT1Fi4a7qoi2bGZFMqQaeCFO2QRO0m+o43yS
NxIUGKjNLO5IDE7Elb5fXWtSfqW9mJzgAvrTjdpWjaz8r6MoOqO1vNwkIibxeIrZ35PZMOgPNogd
Gl3U1j686MTBNhqctFXwSe9cBxQCS8qCHllI2iEm46i1W8nfVZAEtFFNMFZKqNwJwbZIQYUMCGJD
jdqPeQCJQa/nmScvffVdubHUfyyFgghRjdc34GDNgRWxEtybOTx9Kz1Cn2SKtZGiAysYZIvjLQM/
Pw0BEFp5RcGOmon4bhIj00kGBC/6xIsOKErp4+OzQa6OL23CyjHdQQPjOimNcVawRWHFR3frsOoE
dtc5HD3FbiEQYnJGAP0xGuxqhYMU5OIgtIrB8pwcHY6trAFXMNks02nlwNmLQ872kSFMpTqOCtJx
PS+Xb8w5JpycGHcDWr+fX6qWxezN7mSxG+62U+mHdu9nGQtvEFNA4N4q58Psi57ApsTJBzgOu336
O87QYUP2C+9tuYQpDMrE2lVbtm9OAGiPCSsVLdHcadXp95DOEert7cHeseU6/A6G3ZrHv10HjM1n
vR99XzzPx1T6wIdso2QzkRZG7bJjl8iuPE4TBNnR40nmSTbzonuSgIJ+lYfNB8AOBO9KowCEVZ1n
Sq4bqwGKbISQ4JSamiXPGKmubtbNL+a0x3R1vf9XZDNcQ22PLZRmQyJxvW7vI4771EFsZAtJ02dL
hWL61SuDyr78QmdJdLCAjir3DY2BbFJM4b6HA60pesYCdJdcxRo9ep4rBorgAXeTgJdWBS1XWWZs
AStje5e6ZKtbg91ifQgXQGAuMIWaHtX8vNHdwEUDe6KmtlK9nPHP57SyU244wpGCPtXLHNSOioS7
Rqp1rqpNM/lW6peRwtZ7xy5afaWdX0svzyRNXJuv0ELEL88EWIfuk27CQn6bP0qcc6yJ4PnOrteG
q4Wq4f+JwR+W8H0zYUcT8dvcZ9DL7IWmL+vYWCqweNsuxBClUzCSac/rHN1PqGSVmjoFtgbZdHcP
BcxLcHZ+0CvzyrlxwhjVuV6sEbZaFl4b5NfZ9cgcqXA0lOwKp28cmvfzDGkUEMuewcirZ8rTDP6/
TMwjrD+zlbxaqxO4lemNSqQVmLH9XId3YYLy3p46GN9/EaTJg4UmJMbHWh3zJz6JfI8V8RYbvffm
DxI+fqZsvH6niWNaCKpAQI8EIrZO8cqC2YtMbWKuFMvKsnflCQpXtcm330aPQ+tEGaLC+B5TZFbG
wRYCdIkVTMEO1Mmsivz9ndaZFM0aewN5F+nCQalWkXDM5LBKa4Wj9FZLKq9fKCYQGmesBQlOK7aj
5BYH56DLVTeCgB53Kh/4EouvVYTpqMMyxsU3n4M7IlyR7diFPk8TokpWlleWMhOS6L2J5kCy2vKf
njmxj5LZQbJE42JXODpbIuJiPAaEFdp+aq2mHsHi1hXJTXXOZCmaqAOZ7jvvOds1Kc1VjwZRHBBt
7F5Q0TB6mXs/WS++lfep9i0b1zNmzLtEQ/8Kyz7t/3lT3a6Yc0est1nRDM/NC4XLMWKJXs5Y93l+
kvVJ8DYtfXMdOrpogChYFVEHeSJ7Uh3msWGyazPehA1IzxtTmEal2KASbMxomhUzjadUVHkxxdoJ
zGtNltFlXnw/HXRyJkxGbTEUyn6nKcQNyu41bVGyW5BHQ/iHeE+6aMGFDHhFKnJPf/75kOYb7JB/
tTfCp01f3pW5Op1/UmfmuLV8l4QKXACgviSphtVCJc0alQaeapcW2I1Y9frG9eNxeWobnMe3G8bG
CMnSRN64tZSC++5IxKn/KDyG/+7Tj4Ha1cqhzkAQF0BwwHvnJOzbMLARFXQdHAhoxGH8FNcz/cQX
XEiKuM7/1K3x7+LkzI7cyUj0gMGNwOXLwVXvR2SCN6g4j6EK7LnG1FULqKU7wfojoiom0vDXpPto
sanRZ0JIAIh0fjuzlQoIA692oK07ZpdmtOdzT+5Ru60U5Qhc15lJnhbuer5oEPqUwWSTuHcInZn/
sGNDLXXj+gEhlaIcQRCl7QHP7Z4fmV06iuz/aCGSaDgJSgz7qgjcnEqWjISfY7pG9FPVaso1aJBV
XeCdA+HI+I2ejP5dpyurMmurBOFsrhIDZeUudqFWluphF5pAefJWT5WOO3wBrkTlPiROXhtCC6ze
Uw8whPfIcrP7pw4jW02B7wAXVwcsN5jM/aEiafC3gPq63egWxt0i/LqYCo5ujrFWnSksLFyghUoF
46wI/hiOnyXb+hcP9l9iJWuzRiANTHwmFtkFa+iDyA+0Rp8iQmJdlQhO7jnqQTVA7/cHO2i2kaSg
ARkpOBV1HcZdpyC+5l3zBEqtJDOTVkbwERkKoL87NLfPnlzrNU4myAFiROEPGLoDbjU7mkLsug4H
NDavP0XPGqPi3uARhXHNCcTfAD8Xx6JLpE0EVqs4aF34iHy7lNwArftWVzvi/vasVOOfB1Qi8gfs
72wAK8tO5wj8CcM+9DYYARmcVcP7s3Z/RKIyvgxFEHHDRnKcVpydPCINz9lWjb1sVTxTMDEjyQBG
kCdL/JhmFJU/gH4egvrIYsIq2KvmIrlA+fbdF3iMFaAHGSYYb/UMPE/H8tG0hxad3FCi2u2RKpDh
ubxajHRZynsb1zs9cgMsmQNWW3qEDcqd7qpP9/E9MSrIbW5+2vflo2mlPVaAFsYF1aq+Ak+y3Cng
gzbhMRoD++nD5ZRCNA4n1SGBdXdyCJdzi805C5PRpu19Ok+QMGjpCXZJ4Jfk7PJGKsIofi/Vlzu8
9HkQVH7EZV65D4sr87zrNI/bmV97v2mJDGUPR6nDkeniOhtBmbU0jSw0lOeRfQPFoENtAtJUPQNi
AO5CXuocsrTWSluqoFC2J70Bc0XOVXTAMoKLQaX04g/MsMLub52q1RzaDw9bPTRvaRVizYmbaX7j
vpuTMSVAmOxx7Mgf5xCBN29h7ms7ArTL/+BLuwEPxHSXoxPvTInC1HpT/BFOAcDuCNgzI2Z/4NH1
c77CEwVMjCNB7VNWwTSvbGfVdueguo943tO4Rm9hqBzq4AtIN2DcTMW5fLrNq/gLzJOBqK7xgOIL
ipxPY7mg3AbYo+mmz+uslHJLV4y33HUvB3LVTLdssJX029uFlZNdG+Pzzrtu4Fgebl8kHk1ZtPcr
73c/2W/YCo+s2Nm+rjtWy+DS2lmnh9pKja3L+oVbhXhoJfzcWCx5pBz7zti7slz2Z53XvKO+HH0v
/LODsdgdLm506jyl0WyQFqCf28pwgJ8wZEU6IpThOfScidsX2L3kRBfjr6q57AQgbpH9BbuBOA9h
x1ydHKtc27sdrMWuOF+7vvjoUacynJ0XLWLFe+YJgiM3V1iQ3x4Sdgd4+ZmyXxZaww7lGWtCeYt6
aFHbh31t2TVyZv3QkRZyGd8DanZok2C2luQz76FmRKXVwFhWkIs5Lu/GsVMwSWSemJIwOcGIGsiy
UJ9hK2iZXPUho2m87B3g1ztlR7/eoxV/2rT8BjnPnKuAMHxgFpniQXvQI/VPNo6Wq+RwCrvSwJG2
nu6m1SYgL1OtAzwBwJ88eoir7jppO4qHnv0uiylIlQmDLCOMZ+dqvP6gMNnmOgT2jkQupfS8Keh0
ZSVnk2BHZJ35mB8R6Lifgmq+sEmyZRqgKgCnKbN8M0YpH12p+sjJgbOxL+CzpYEZ35OZfykaPzYu
fGXzn2quP1PesqQFIvllgOnlxyI40aJPRNpbj7TrghHBVCmusRgEATNcVuNAESt6w95It5X+TH1X
e2YqPYg4sFnuJLu73Ax2ApEgjBaiMfuZa0UWcY7LlvodARbOZ+pUmQR350L3eEum7Sqz/S8LEQoa
1Zr5sypIJx7FoUKum3CrgyTwSRzOqpBXgtImX2Dh7mmM30I2aYUCF2GZ3NukF9WDLRivZ3T0B5Um
hEWgT18jDSLqKFVwTZuVXfosUcEOw98RC5Ja/iD7YITmkPIjXMqb4vf2XpCZNHwXObPTJm7wbzyH
w9UK4mnacvViGsFfkujFf2UdteRYiFQ4T376zqlCOw7TB/Zjaouist0bIWGZQUiT2EB7Nm5DszdK
+xeYjpGBAcJf+07IOq0aDZM7HAvrOzeZ0UA/jly4GeiOPviHLrxeBNBmBDlL2qqtfQFnPArLG8Ym
mrc9dbUAmmGVxLZRuEtYnt/nTmeoutNUXYb7PMs4Iw8dePaT+drIuIjEdes8JiEBj75JUQJHzNwZ
0djBXZx55rMmicXACPbWswPvpbjhudRTTfZfYZc435tPcIgaQYwauhCeCk4dw2dFi5Hudwvvc3K8
iG2m13+HQ7Ikgp2YR83mh9hsAIzVZkNMB1OWYHNqwMRGT3ZIOp5Ivf2lodz1mHYIcxmyVHEsG3wF
WEy/zmBEppHGtU411DhsFIcQJe5bVnGad1+fKXh0c/DeH7UpWIfabld9N6KVsdHv5WADGU+MTd48
2ODRODTQ+NUpbt/d9XhzUc1uk5oxgOtnadsJAeDNtTY4dSp1CVaOz3Ld77K54QNWjo+0BPqI/yvT
K1aPjqRtzwh80uolRenZIm9zg+roVGF5UppXFqIfGzELDNyyRptNBSwOC8J0l0Jm9hsFdzB35u3r
XXMr/r6ursTG43S063sbARQpQikfW9SY5UL/Z3s8O5m1oWm0DUIS6/osdP3H+ytBh5TrbypULM0O
38XUmsDdhsrKjUTEgm6hirPvsfsqream5h849q0AOEwMZR3NeOWvQKgOBTyj5DTrP3rXt6u1T4I5
7rU1UXDIG5Kr1vaZJbh4Zvhh/Rwqs1/BqpdXY0McpbkE20sF3YQwFQMOgNGMbL1CWginmqLzvWCP
Sn6LRIZKBvBnq25R/XtanGWpwdnTU0XADnhbMwc2c2a0vyTW6uE9p0FDMK03YsDRXSviWkEkUBVX
oScJnPTZQ2cQjcaALV9gqwQBbWqVjBzFk/aeEi8esiG6g8cBfrvrBVYDEOo3MM5kKlpaIH2+65WA
ICySthL78TS9WolBp0akNx2FwSnSfo0c7LBgkAjSoAz+CNyA2v/0F9l+FMOPJuDhP+vVM41BlPw+
nERAKwlHsgUPNBMSwJcdV76g7S018MHjvA+brVQAAuCEgHKyDm3fHW65QkZ+Ck5WWweRck2LyPO0
iAwEwa4I7yCv62ZhLd7FTVuPGvvadTOZuTnrYa1Ykuoqs36LOmLajBws77Fgb4hqzoqeLKeFQFnd
dvjc8Am+LW8yY3Y2p9pB5+dQx8GXjGodqDUWVowPUWvrKUvks+ZTvKP09Q+52msO3AmMoG2oUVVY
2pAoQvx+pLTDdicR+J5KnsbpNq4qZ/MhB8sdeEbDdjkCIMUYfLYUlZAOLMUUVWjk5XQPXRoa73Kp
vKponjeUYSND0xusyObVOd9RUjLN+dtQpbPNO0P+JADnfeEzO+vPdWHi267M4fWU/MhGhvTUCwdF
8OECn8n0ws2Ca1LigwL4Z2yOE8WG7vyTBNqq3yio2ACgQnu1gxO9DPJxeIpld/ch1XOEDeJBxWJQ
5TJg+UaFkBUqfhbldeUo9Tfsq7EuG/parxJiokOp+csvjnCGoq8JFmS+tJ9INrMVm+96SwCRWPQi
k3sWVLqqLfQL/LwKzDq5JXk1vfxGCF6zLqtrB4uYU93AgauPwrd1GUFNFx2YfsbcClhl11XH3Gkf
C+RlIeAgMYp+1tRrCw5LSrzA/kig3zcMd9nPptAocROmIDqJJn41X8PhNCaIOWe4bykPzVJM4bwc
H/IwG/w7k+tN4RNdzveHK/M5sJtQ8lyXVDS1iiYqMO7W7r9ViMaaOQKj8HEGfny4uJ8feLUlce/0
JvQwsn+29SxshAUaQvW75f5f+FQgTYvuEk0JFxRqg4Hm15d4OG0aCniY/1o/XGybB8x4QzEb9okK
wI+bZBWp5Bviz6ofy4aXiLM/oiZ/Me6+JCRc8lp2XA6l55YEl7Xoixc+lp8wAmJc2ON8uUGdnuNn
BqlegUwRmx1JI+eCyO+zLLsPsXFTCeL7bOwJj0j7M0saI2L47sZBvWvV+g4eqizeub3scX7eCV/L
mSCLUM4TVMD7rlrJAkVOwAdP7SV/qqoLjmW8tPBV5jt/q/tIXFeF1qlVMsq9eERw2i4yp57zepxc
HDITD0Hjov/qE3a8JtlnHJO+2I0g2Czkx+7Apsa1gezVzF+Dom4wcMUB8Xmo2OpKuqKtcPWkCthy
mKPRU3zcmgtL/WpGrX9Gfwls89MdAPTnyntlEj4Qj9Y5JC1BGsHS8xq6jdM1CCqFdMAu5axQQYAS
sz+QOP1pts1eKypsl0hfhhIEC23nY+ymjFZxebSvSs4GwA5H5/k09DX/s8amM5CuQEZaqIJmRPSF
yT1e4CYxMEnKcnHdlcuHixk9ns1Q892rnSiPrCHjmqCd2KvnDIX45Zt+sSsAz5qzN4eRY2U8tXBT
5Z+TDbYDpW6nYgj60WJLCNxUt4hocghB+ybNhDylKJocxjdfBlbAMT0r6Ak7ueiMm3sd5gbWez+H
Q3mdCd9cc7urIfE0wvbajWCB26gDBvVCQwR1OXxgSghp/4Jy5i27vdynGuZAVy7sUT4ka8KCMmsc
Y1AXC8KWBBHyI5J69sLw7dfs1f8VIKdY17bmi8GNhLmLOdlA1eKF1NdGsLYIvgspqlGPTOAllZj0
w+oSiB35OzvBEztUYMfYcsmq1cixjLkMk7gHPqcUdul4D+lDPU/SboHz0SYvUZnRqX9byt/HPVkj
MQwYgMlJoCisnkO27Hihlfdp3eBULu51YQqZDTtxbzkdMqAdcdQZO06urucZIlzb5fdlCFqzpK+I
xQPx+Rak40jin9iW363Hgss6m7xS8K33jUp/d9F7rjI2wZ5lGM34dJaaCCu1HztNF1uR7uCMGCMF
6sd7ThkFRXj+EWNZX40n0N+T+0Yl9j4VBnPxCDF6gtvvihOwqKQWVEbLIdYs0qV1wy11p6pT8Fqj
6N5qAdYKFZxg850qgr2grNznYg+dRx2Y9uNzml9d26cvvmeP69Kp7zqHxpcoluELeUrS2eVB2Y/t
914NjvIcwMzjHP8OxC+IKbUVeBYMeTscuNu9SUkULWoX/CmpMbqUJVqesH/2YWMYR3PyKnq/MhnX
7BC6dQ3d9C4F/y/herr8PjmBBP6jUBJkgKHhup96RPSXa02zCmZOWt4ofSbx0ARnQG8pUmFgx0R/
XfhE7tpiMQd/5Bu5hdcOQBvuiP4jhmi4j/7bZXd+yFUoftt2Sb+IGESOD6JGNrjy+4wPURqqXiwg
b3imxsFcFOaQypYfBF9L4ZRzdra48k7eRkmceXFx6kXx3hGDCwL20pcML46WbUzhSFKwqR3BomO3
uoIkA2rimfGmzl7qr8M+N9bCZbdB0ggQfjcwshRbQ2NAhgP0qX3S33tEgwhLIIIBMrZy7hXFnVLM
yvUVuodykrWJZVIUchPsJUkZ6EghgiqGKyy0XCiHrvllDYciW0pNXsixPVN3egQdHZDz/PJJBaSa
/ETNsiFwHS5Fz788e/YsYICHY3J+HGRVWy2gsGdScP1qKZmQOZxPccxGI7uvr/oFmHdvzDmgW6oO
z4n4GfmnGr52KIIfmhf27FDDQpp5USnOz1XFQy96MbhoNL9zW0fpDEOXiT9yTq3lB9442/SZWRlk
gxxkPQFWlRjyQJ81n9H4UrWGiVyEvWycRlIVMTMTTBWVtlXkMCu+IB+pNyz8rtG0QIaFT3gQJSCf
Q2fuhzckzSX9O0Xl0aymB5jLzjDEnWp8pbIWn9gW0mq2VwBHujKtECQ7bsDmGoS2WSb7OiXhrGRR
xiGi14+aNigGdsGbePN9NvotwEhn6CXgAr1YCAsdI2s8faRCwIpeisCTnBEAUAurkt9wdFiXuc3l
Ky2+XTqN9AkUT26VUvB6pvLRgfkztGfnDT1dhyi1F1jZvctDK1cgRx4im+MJhPBa1+d9qSWwSA8M
2cl+UIWcVq9mWNM8A4sx3JN2MQpMZtYBgaEdt0hytIwMxmDnxiHcYnIoabZ19xq9m6/X0rB0Omp/
VWqB4jUKOeoh23DP30VXWVFE0vTL/S2pEpcBkAb8xcH63CeKttgGgBrWbzCnwKNUO7DtZ7MQ+jVe
5Mk5Xj0vVifPUB16LwwF9xd3TjiEOykfnTeekE8cYE857HZubC1+GRef/7hRxObbXoUOaFc/mmJI
5HMuOR9TsObHUxx7km6LXgi9ckHvq7j87szlFzk/q8MK33wONUeoLRnTIg+cpnMNoanGx2kqh+d2
ghu1nMsFjtoUMA0ELl3gh8ExJH6uT0/Y3CusWw5hvvU1tn9WbBSADTqYUXXRKSynvJ1Yi5NiLmvk
ErJOOJ1md0c68bKx8syp9z2PRrjL2sd5uX7X0LA+2UKpPtc6M+YnvlH3KESwEvrpbqqmJEcDqCPr
iXb2VXqknVqhTpCJpozCYv422oeOJU+URjn9rmpNoMoy2Ecp0aQRFRtIpEQWx9xNWFQ2saV0Obkz
kvzU59p6tl7FernWD/2FbMkyfmxgwf2Gexi5DExU/Wn7Befe8CVbsA/ZhcDOtKunK+rq/VPIn1dR
NE3UQh8ei0PxiwyL110zBxV8xmsCOvKkFOdX1Eo4L6F04mLjJOOIGBIu99VEfs6bE7Kf4P2Zqbnd
Grr5HVoRm670zrBEioEBGaTIRiLGWEg38s8hDflVCXv+9LvwaN8QC185LAeb3VgViGUW+zxg5ZnX
QYHO522FCWRCVhDhNKERpl1rzUzApmZDE6nLUZlfozntgEkXh5L1+aRiITwoiPBV372JynNKS8bL
yLZCKJub6YMRq0kIxJ51orSsM62bJbIX6lGEWDR417M0jS1Fc+sbAFawiD0DV/DOJU96Dwla8/1A
e7OJZ60Cc2ZnFE67KUN4Z9uulW1slR0I/TTkfw6U4n215jKo1STN2EOuSnkMBNjThsIWalp6Q06l
jn9OofN46Ii8cZ27mr8YKTKj/CHAbQ4NR6JIHxbkWzXQIcMHVaYA4X/XZIn/0vsd1KWyyxAj507S
JkFjrD7AZCkjR+qTQKVV13VQdeq4Qxc7JsbrPubkOvsDttk6r/Ala+fO6Vii6E40LPMWwFYylgbk
K7a7KSOhXV/TJ+Z5hecCZ0FF6TeMkQlt5uU4mami5ZTgEoU6vCTeOn3w/EK/uJMJFUkrrrxvGCkd
Omyq9m6/DzSJtQEaYHxJQfKoEQjVwiNjAn8xPPr3AC507uQUQVcRCNPFZ5lMOjH/nB1udVVWKgtf
FwnE5eITVIU+2gkq59IjCEUZ9ixzR5PfaoF32+i7S9ngMWbb/QUNXy09AgmCk6P0LblslgY0V2b/
5MtI362vd6YzBi+bvA7i7FLd4y1eK3PVknyx1xAwTv0PLEzr8Y+BYS+TWBv9yu74Ouh0L30B29qq
fQDZq1LYkX3NV684KOOMjIokDhj58eaOxkKsGHyOz2MBPY9oGxe3fiXFpYrCGAuii9ibfn3mPlt9
QySqV1y1Na2ktJVlOm3E4FPCnuSdCfFhCDdcmCT3TWEh4LrdT0uuVaHFndwMbC6/HmJuo5CJ0rwZ
AI3GosVh2Bha7iZ6zZayE7g0fWeWVF+AQdi1eQOqAWdo/b9uBd12P+9lPxu/bS5XYpPRISHB9HNL
Ok1s5u1lMcU8hqvLuziG6DN98wyDzgbiagOZnsxjSjDkD2SO3bt+FXNqNcuJ1mBMqRLJceA6eimu
FaWMTQBsr3NHdmsfRPMQqqqf1k5H7oXSjLGSbCCczOANRCZHW3BNG2s+ECqZ3tX5UhBSu6BYdEF7
cQDbNMLryhrqFYr43dKiA+6o5Kh2zRuCf3cI3ZBmOVwRFamCE0XK7XRaN49lNlTHhZh5R5Pe9cJt
Ad1fgaQNdMkSKjQzlWWunszVa0yO6dJTMKFBgdlROw/+MBQ6RNjdJ9MvVgtu930Uos5En+a4BTTl
2Txq7bLqkxNeVKol8Q57rC/P2g74ytbh0/OjwLVztRbDKA4Cy+QJXz9gjnNvYYLp1CuQYPjG3rfF
of7XcHUdUwP9J1cciw36NE8k2MFtZk4oS0IHzpkS6H76K51/HUsXA68wvttA8diq+i/GJtDoLrRg
X47GV4hCd0VcQiJ1B+MCTp9zFkFRVRFghniNaoXCj/uQ70b5VcLADaZ3c3CHh1OVwJYRVqY6SfbX
PSNFeV7VHkUidtsI4izq3jDkbOE9IUand/rsoR9DlYjnHScPOskr4EUGeIKr8nF95H6nWvXpzUE2
LN94iZEbrOVOwHraxHjgZAIshZq50J2tiotFQrOTSt3KZ817ddbYAZzmv7deG6ovtcQMySNZu8ap
ChUZ2jBbMgRFkmx+8YeMZ5dPvTyTUKmU6JV//qCcQANb7vXTf8AIs7UMVl+qDAYuIBG4uvKpJARn
tknqyHTLnI1qCIcrgUHO5Ufb8L+0Db7dlbem40ghv7/Vx1Gwqy/XWfLrSkNc8TXLd1SqTXklGy59
uG+ONgNClsxAbptYEDxbjaGhoJxTskmWx3fMgJWgcT+tBya/o/SqWIMHGuIWy1mvQJmWAGRfiQZ+
kfH7BuPunVSaxI5knNQEmxwDUq3363jpHIIjJsQLiv41P9ycIB3nBSRMHeUI9ZuLtDzO0LCp70AH
SM7fnF3fGwHgh0UIBgfQMB+UZsyNDp7QiBSjAh8Ki8f9fCoq64AVonV1NjrUdhDSgehJhCEzEoxi
QBSpqa/OqmxlJyPXVGxMFg6YKWbY+1zz2vNtDBCAVEcAOS3NdU4wnnxUrzHU/fLP0VSCn1YH05m8
s9QTgE5UII/hmuT5cLHPcs378qprlhijovhlhFriqTZF3/ek3Vh8VbJDfBor22Oe8DUFsH7pi+hL
rSAsLw6Ccrx2wkwg6MRm1YSVQXMWzqIg4/zacmtwIIJCIiVyTjU3pAluhAlWkeRrHOVYtDZq+aJ4
NBaml6eqyymjZvV0NRei1wQRDTNTT9YxKFDnqr5YthVOrEuo+QCU06Xlskw/APVLtrcNTeZ7mMZr
y00vVF0ThoevSRBfVqfbGiDjMxbxSq10ntHeiYoHR4R1jx4ysbfuW5ouPcJah3J0Ne6OFLOgL4rS
v2MveFfXJuCJs5+zuBj2swZcXYPbtA4B5m4DwbdTAVprnN/W/p7SSS09w6otzMhKdFOrUXbfXZoQ
dNI9IDFOhkRKQb4YwPBXa6Vu/5iQJMrRbwBCWJgkb+XN1NvT4ZYXQEozUBgF4crh/snh5wwn3OJ6
yyogi/Hj/EhqHXbs/chenOzr0VyJwASMf2HIVs0FzVa3+yXLK6Wvs4E1nxhjZnodtFBjR526aBQt
UmTpFBHkSdzB1XWN2d5QuvpzYEjmDfeuxrhADXTPekcdXjYksTVdltRg1NMDdG6k03vX04Xyw9RJ
Abz0BIgiiQvx0O668B1P6spVMfVCmVwzedIATImac+cchkzSMa9Hp45931Upnpspz5cKDWOGpu2/
wpplXwLNchCZowjnmIjZ/FXq+12kB+NbdgXOMjh/4q/swb/jouJnc3xDLDfIlQLsMx0qBk+vIzuy
od1mj9gCJ4F0TRZ+W9bB7fZR2tklnOwPPj2Elb495hNVTNt2lz4ul9Hkav6hoB+p/9epCl6Zyoiz
Bc5I2q4FeGc/VZpbNLGzA+S/ksPmUSY8DrWaMe65TYvYaOAEW2zD+4775p5053CEfyLBMij66w81
/dHTu4QCbfDZiTcynjLV0lchqWv0aw1ZYcr50AXjNd+oso2WayXr6H/XwvNiYL/R/VI6QXiL/qtE
hM64bnGtEjXJg+qnLTZSXeBI9uS5AmRVnGgJYl6L4gxaeRWDpvZiygegKE6CCMk8Izdx3K4PHHXI
ShXq5oVfyGh3R9rShP7zxX4v2G7e7SmcaWW2I9ZnSzR9c5Q5Ohl9B0rxNj5+iDne8BL7yUXserWG
5LrIDEedEYvW1B3I0W8gN+MRitjiljV6ARTaO9ysEnfk383AHJ8LX+jnFz1prmILbpAk/Zv2RUEh
DYlluyh6ZzuambOYg1VjSqb7aZHrwgQb/DTi1tEf5wZ7lB6rG4YIvQaaIBQXE1KoFKgquZt7d7h1
toRWUQ9dDVpG/5iG7DyZ4Hu50+ixl4xUH9PwFhUFujsFaiZ0cjEE613mo66cai2wZyFMT2hQdleW
b6m+H0c5f2S03+OKPCwZHp4aFzz8sE48pP5tnLirRs5U3Okp557GxRH1RhxY5VRq5aV+Te9oPm6R
wdF3nuh2amCchMsrZwydPfOwEllxC8z44K1X3CH8+cRu3vgt55SRLQdtOBohH82NS6o1qBIHM6z2
d20HChVlZAMYuCscgsX864/dVHtKaOWWuIJ0w7cJbqT8+066l4NEp9ScmqrXRwSDUKyI7zcbE9/R
zOeRk4D6CnkEDxes4CwMcEi5eJJXqMOZG2H+xjwRk1pVa5sm4YcnPeo5ZSxV+Vg7f3wLyhCzR+Z2
uZtmxpggtZlsavF78/57zcfcTb/QLVQ9aPt0CNA+uVhjOtzc+a8IO66qV4ceRC54eBriFSgEvyQM
Cs6UOHce88jylfDfHy7Z0wNw03nLiP7IyIrAhDWy3H7bDkOTX1rq+G1pliVhKxxw96yqAQtKYV4z
cKC6ZGEHXzhjL4gNoga91Kz/Wr/fAHgtAqY9XALAtGunODkIb8bgZOTPFFBOldHkDRa/s7en/y4t
9jN0MDBWXquS14UofuBwq1RDWlUAlls5ojUEDZrAsu2U6QDIkDo3Kwwpih9jDjhIjumk4L9S8Yie
VhfEhJMFI2FUxexPn+V54I/LsQ+kNsJRiEIbv+oWFOkHuPy7E5nCmnCSWsFqqUUPybQ7towEhwMV
9roEGVlyp3F+f9MiajEwyx3NyblxxKfeXiNz+ShKLqmC/glePxnIRX6Bl3LRKxyQrwOvB7pB4eXC
IXhjUf5YT3cY8DQm2/1BBeQqaj/CAP6zh7WSgGtZoI9kSrEtv5mhFY9TZR7FWEpEvxYupjvynFNE
oqeoZyaYdad7AJ897kgCj9cdkMAn43ItrkzlI7N1xVcvkcusHGob1d4ovDB7pmKXKjs/DPuzcIJb
RUMvYBLmUNifd89JbauMzw004C81ODLXQ2OAtB/fV0OB1nXoUFUzBKb3X7J3w/mqiwiMDTSDp2H0
OXPaSZYyYJqVSid/MxtzaJo9phEDlBMbTQ+q1/vi3qv/IHiOEeIM/xdHP/TfpKpZQHsJAbPfef0u
VRZbxV5f21byD4nLQAQTHW+ZA3XhkVbnPpilo83TZnsInl6ymD6Y7ywEJR5U4fzWJc3wXupBnMxl
A4QuUAPSTHZQAzcCCmfLOefuL/zpwgduL9FbV03UpjU4y2hFavzJ659D1qQ9ukehSDSIFXoHBdWY
uw6W6x63YLAvTpuemoQ1XaBU7x25XwgHQLSdDvf18MY2sCcFh/LNeg+HIreZE1CulJJwp+IXQjo/
8/qmr56YOijDJwJZBY5CD4a8/FQd1KzLk12ISNWQ4UXnm9WTbBuqx1a0b6fPE1sWBRnD49WGNq/g
azF+QNP4aUjgOKux/LAeXxwUesleuwWTs2NujqkZwiwaNaGgPWezkiI2yYk3/y+8w2GDYvrwp0rT
3mKFqEmjkTEMvQMZQQtUfye7uP8ekhx6vTyIKpsZcjoTMnqGXwHSyuyXRRYiYejspLv/Xrlc5j/F
Nc5Ff7f7wNs4vyU3wp9pZlQUKl+DA0lDQUgrIysLE7hBvbRFvLoGBqNgCY3DmQg/pqIDIwmSclJc
DG8efw8lQENW0v4WRazrLhgnnSkqIYxrcm4HZmwAeA9UNxqI9iD5tfOQv7nM8kxHIg/w0ImNL+BA
Ib49yGlXXorDPaoExN1LsIeKOMhgJcyclXIgzxjk0T1j4/1EXOFSRPfz+B7ypNahpsYeS+Fw2IjS
oEpDwTi4zWKF8z+eJ3gTvkCSN1t+yznO8LAUo423dbY+UytWmNVxPMFJUHUSdxMdWrA8FOMC/T3z
RursSaf8+ZRG4sqDq20+C/UkbDhEikbzHsH0uknhlzlD1udYNsB0lBEL+mOncmf1vRdEUNeR5cd7
7u3CzKJlx6CKZJl5qBV3iqwLNomDGSDpmtmEFrwPaMdfFBn/uLW8QxP/2VZeXm6DXhaJNetZsHFJ
o+xuOlRM8ZTg31iV7PBXJZ5QbWNO8etYKgL/QQd/joL0C16FwlmlWjd3Fa835c9mpWYpKBikFP2S
BAAne0dtGJMohEmq+r9gb2ZjfDAgf4s+/CcqKW8r5oKf4YoZ4g4EjadyKr3/lfI+cUVvBLxM7RHV
zVK1daHFW12BV5tXXNzUGvJi7gbbf9hOZcrrrmDpbHC9vedeAWhuMMabGQQ4V0YI62f5YI5GbLgH
y5gupZDtL9aN3QBZbRc02ZbrmCmZFci8O8VUllUJ03eSIm43Y9/mXwYjalF/JYtSncsa1LAPxk4u
4FXfLRmrJDqXL2anXdsesz/p82TCpO62I4hq1+DFCHVbVTNNGkOv11+qjWPE+lyNjgKlIjJkqTqf
7kDR9ncE4cbvJct/+nuoRgoGdU8wBUD1LMg2VxasWkAlNyH88Lu8oIukH3j7SaIbQdTU50V9Ho2t
Smbp3Ah9c0fcvxHeQQoh27TIz1W6G6Q9DFJ0zH+Z+7iEPwbVgcgZpSLWXPh8Nn/4fosQ8FUl6t6T
iVenVAoPQItCBeaGoIYBytTrSg8sQqpuVpzhnRs8Q0tttusk5TW53OyOEBd1fCJez4+nzQLAJZk9
A0o7g9LybstCIqQUtM+FUw6Y7Eqtc5GECQkHK+dVizXcrCMNiRaVo7a2vQkhymOv/mxyk5w59lAC
1WTWeQWyLKFXfdfCZwBNhbVYgipuH1ORZRq3SIyCazDKf3nXn0Q+oYbcpOrnY6jnf4HBgl1n/jEl
fkL6Jyot/XO8jwiihDwdgJ6rLGKS3OWdzI7cMl9SijswmquHxPZ7vKuvCSyiP5PR23y6HjReGDS6
TVdRCPkas35LLTxcY2FjTi2NLiDJdSVRZ9T+tuJWijajxKbEpnO0InoeTX5JFny6BgOk1SyrzB84
/BbAkyUwsIdoRfdwyKz3iPy2wysdkyIVOpDrwA9FgW9NYMID2QaOk7Cfm5MysQqvwXMN6TkRcZbn
zSZQjMxSsvpuaO4ps6MKU+9e4P1hK/CFAygTZhRX/0iimr9+CfTWwSkY8bHZbweKzdXPhBLup9yA
To5QOfsQ5mWNBnsOzgxxUOXtfGyiwhmAPp0XzeSL8uWpvZe+rmOMRxCQnqVBcBHoWgrMz26PJg6N
cZX5F3IFgQP3J2FtLh+mibAYhRKKMtOWfu2AVv+Hh+impviIu26x2xNImfT7QUKL7hXskpG0LTGm
QSKfQynXZXPgPKmL8XZ557aDbPGMh3QEndyCeoo+/nY+034EaAAVvubQixlXkHdopnZKqS7UAKc7
DN3+FyhWJKtBEL4IX3Yd+DnDafGZ8ukAycp0xBTGV890eTm9yueZfyaM7pM0dMiESqCIDbfQDvBF
/Gkm5xfOkoiS7joUJ3k9IF1TUoo/grEdFXoX2I7xXdcQLLvggsTG/an3nGy5U8Fm7xlCEBxwgy9m
XD9dN0SQjzvypSanWMrL9aKQkLAXAStj2IkYwImphWPY9NBiNySSpUoRd8ovFhDKMkGKYmcMy9Xq
pX7iUfVLlABm8D76aqAaVjPTbg+nm599KowuqcdJT1PVIWgOsYlH/cdztRGl2LCD0czVvCYSnvWp
LtHsaJLhA0i+cHKo98jxDKPX+PKUAm7eViEZ+XqMETHT/hFxK3XWVCpjzjmMv1rNAscdrkuiP9+u
qYPcvikaBQoGaAbe+X+O/JbyTWfaSVp3t18Uax+BC4ntcS0PR45YBjcF4IfsLGV91zIin36IUhFD
rEAGkDzzZcQXrU7x28MLaOs5w88sIifSzZ0DfNrTkZSCKOsTC/J/aQavi3wJQlGCf3G0NiPtkyMe
Ho0x1ssmbExpCBg+asSX3UXpiD0vY5do0gn9EPszOK1UdGtzSAT7AXLiHhE1FVtRqXIdd9fdi/Xp
eABv/Z2NygwJlpZkN8NcyfXBidqpozXjFkNymWKxGGRgb8+kAQKhuXDvmj27CAm4HYaUevIRIX2c
DHNLtA+bP75HWayDkCWCt50H/WrGJ54LL+IMB+rwafoLbFoT5lkgmTlYimy27ThsDTwkhStE3Zag
x7N8DHn/tQpYidiZp9b07lXySG8mPIcsRwv/xqh1R94FvQSS5ICvQAF/H0BU5ube5K8ORn5LejGL
VL8txMKxLqnNOtd20ha2mnvR07AOfMzsa46VI28rvMaNFOWfPoU6LUr9sY50qup/UJiAY5fXotVp
yq5hNm0JRheOcS97o1skVJvhnL9Sd9vV3fQGKttgQXRsrbjeF5c+5mH0L4hASE7g93vSaVkQWByO
sdslyxrHgA6o7g8HA6IldgsivalcgvkOEvuF5l3wnELz1ZBPx8Dd1Hylpl0w4YgLcM9efVzIDwsC
SYV83DOsYBLz6pJTnWbU+U0xqAQONYOq0+TBpFEnuYPaPLu8swXdyliDCaU0EuXorvFRPMdg9mQJ
UnAWqjpWA7unESDj7r29uriYmwNHYTA8Y/KJA4XQauPwgD5VZGpPLVt+/rpZKQwF4AQVKxhK7B6I
DQRgUawZMb1safcE3ZrUZc+WN+9SnHDnAMOfT/aVFzYwzV7gaiYQp8EJX3Ipjiz7RwH4m8NGUO4t
HQCbK0u6h+94pC8nxZ5rLVBwVu+YvPC+e/QyZH4EkjshgIkejemf1uVYY/14OgV7u/Ps237uXOii
8q/iMlAmBp0M4BmBEHfT4V420Pp/bAHyKVe5FFjwIgjTGB09lG+tB7KCIQpcyJbxb0cxBKcycuhl
h4UJfXPlAgIFNZQwHitKIq8ok2CJRi5Lc4WToTmtMcTCgUydrk2NCDTw9SVMQsUlZaYbyFIGrNXi
HwAAqEZvN+rXhwl3B3g9QWv2iJoNTAK3rlB/bncXDrZXDaLmTdajtxWdHvYtQJ+SKIkpFRG5KY9m
+VSXu3E1EOs7KjdkERg6VnIGUz8cwJnelGkGaaxmPSaBLqBcTlSfeeWYY/bOaCauvgMx2QSqgHyq
lpnF1p92CxwSdFE38OfQRxLLSteb8mGJn3BbF/Vptx14syUBGoD8YNVSm5xmjeYbdCUZARy6r+wp
WF5E4h4i+rHT69K4YcL4WWo4kWrUKuw/6CB3qcxLZhqTlWUvvaWHbj5VlpRFqLcQSWeicuCwaFp8
SCRvZt40BFbnj8TVAojF+2OewSNUz1CQwM3bmC1BkAtrQYF4RhqPdni8bSyVTyhloohBIr0H7KFH
1NWJJQDVgt1463R8/z873/m7BxKeob9DfIXyG7oRhtQRtOadDedE+XSPX3t9iD+F2TB6PBsOIEKP
X7vVpEqKiRPy6hxPpmI5zx8mT04FJ5EdVpVFlgvukixlzQhoQXpv9OxscPlj0Po/VieOasb9skJR
s/zTSVQjgWHct9BdQxljwuhifYEkfxblull3dkrhtIX5W3ti2LHBFuMsuj2rwCXXFw7JIeXTZlai
ikSG8DvvHFq7YQ+5sqUyW65bI223hcoCwSQk6s1Ik21xXQUXRaKTh/+P88J6u6O/xVdTQyF30tAX
J8ZaVDOsYeVH0aKaxBrZe49+0lXOQ/m2PJypqSi4NzWjRkGiKY4zD8vKJXv3F9y4EUADkkOlXNWo
TzKdv/Ln0T6JTSqWGsX9AEtz8Ni2yTK/X52/Dz35k5AS7RYXlwnv6lkxpxZZm2AdShdC4UCUtu73
VRtlvjB5yI6IalSRjVDFvKZIjSILYafFg1OAf3qFQxuzJ1CxXTpalIQKVUIdwPrNEgT9gXMHf8Dg
TDIymoMVrhK4JBGyDSDsNaWdF7sEkuTWC0I3nO5CdqcNAjeBa6jMKWanLu+PLUiatXhl2Ii+YN31
RuhzZDmXAIrTOvW4C4pvbSafwoREpsQ1cyzMsKoECAjqmOlTg2AlN3NCEptX2Lm4s1qUFTh8gM9D
7uSoSGr+9WBjDLokTICYmP4U71Qdwz9ooBpBlUmAT8TUm2Q7nB4OE/TjwI/JviOukdc2qu6Y+PMx
j63b2frV+Ln3wBMOxM9NeDTZV75acW7l5jM+1ItsK2+/SUBPjHCzKEbsDrLAsI/kSXklabf84AIx
iVW2CpR13Jqldovg2WXwYy7d5DU9Ng3p/CpqG7+4/KqeO/zRIOsayskq40Qss6MDYP8+ixNGahSs
WXha1g/RONmR2paEHXTGZ7B41t5ss+9aoiyQQBKmdaH2FzWYb1YGi4MQ396VLuBLV1PruW5mY9wf
zJNFXK0bfv/pB67tGHFSRWCIaaStWu86kCn2gNM3lwDeZcu5lYO9bORobTS+0zmYwk4D2uWwTi1I
qu3DFyEQoUJk5xWqQb3BWxyKxf0FLvEmh6S0lYMekYp6zacPUNafIZQkbRcBP4Y1q2M/LhkAt0hg
HFLWWfpvffYo3aEo0Z5tUc0AJJuAhhPN3b3UpjeVqek4pV11w8sQoiBTFtTgIAzFz8QrVzQBJEri
FX880w4ljSXNo3u5ZAxyU+fuuivTP5rdNj1ZF5D59qRidPhRsWIL3aLtiX0enVvHoneGZdYiUzrs
en6PVlceoIPCvvhQYLmNjS/irCqrh3YignYOt2iVzzNbC+2Hrn4k93uI0L1GDR1rcdNkerDMJHdI
/240ynvt5gz1njzwY5oMXSOCiZoDm/Oisn1ZNbkDbfOjRcuwBG1t41qJfstTRYwedDgFMDJwgdyY
P+3B2mpPMcCLZrmG6iDvMj5nhgcrqLk21yTThOejiwvXxOpfPFiiKKvS/XOi1qJbKvb8EHap5y89
VEoSdb5KwZuawPtLXFAlW5wlkmd/gl0gHjnD5bQ+xcEwRWLHQmJyFCnZaVj/z0t8J6c0W5O5lSNK
zZjI0pzvsGT11Ey44uuwWHk/+w8gwm84cCD9HTxX2pdUaX/xRscZMy2QRXSXOFzFm8cOmZl0kj7F
PlhEsVAm7Oy+6ORb8cZJygUI5eF7zNTk+8f4UbzUVu1r0FN5vg0F+YLvTJcTKYBetdHZ4s4QaPKf
C/SjKdS3twrLbnLeKA5uushNgprx08+r++x4WKIVT/l650rPUr3ESITt0aHIbQWDAlgllIRIszuc
qFAzvAi6BSNqYV97GzWEfqdIi0/pOEYKGAw3c4aHcSElrh3JY7C0is12OMCw8VjYnqXgrorp946Y
bW83CvArU26YufSDyccWiiPftd1oRrogcqQcG5eAtv5JvtbpefJMyJCnIanWECA+O6m5ct+EHeCw
WoellXGKl0DPDPTnctnCct3IViljfjzSkGk9LgbCZBNkg7FHI0LtwNvw71CYa7ra2ktRt0ut2phM
VZt7oqCW7EQoBKsTwBeszU3v20wSkQrVu4Hq2yXopQmb5HKAFcTCYH2BDpd8gvz+u79JSYUDThAe
0aPjsfwmVUE2SQoowkDDKMHuP2UfR9tmUawClbOhld8c5GC3jcQJhmm8VWvc7mcENWZK+kqwPooW
VGlTyCslwbaglIyuW+o8FM7KQCH7ki+A/qMm2Ql/nhE/onA9vOLsVpni0iMechnCJO1N75aNO/Nj
B26BwmuNPW69C+F35fD6Yo6pxoId8PGQ9JdTcElsGDOEtScnkS0gWz8iDLiNimKkvyLzO8ivrMk2
E2DOmGIfOM5D1zBIHGL82oZeVj0fkAXhkzKL3fMWGJNuMNQ2XhFBXp7FWSCbFW9H2Hs9y2BXpUVU
pwPecIZml5hla6sk8/NQaWcz+PLPgMg7yneKOq/K4oWG8MEXLTDxH/URHS38d9TxhEWAZrCxIyE2
t9vdDO51LhueG18/hVsqgHlrLGGXuruQoYx7hrTA58yV9LSNAYQCSYOX6MF561hDi+PERIyzFjPe
wMUJypzwtzmtXMH4casM6A6THOHxwKg0bmmYKOd9w4ZQuVeGkvuQsb30PsZ2iQ9fiLkiqViDqOTw
Ywm7pjLGiB17duQlfbywmiB4ny79KX6yK7LdyMzORosLfDUTpnJxL3bQfS3xWwnI/yWUU/e3xfXR
rRpEHYdwU7eOvgDoq+DEVFHuw4JYxGsHTwlrZYV5nwVWdzYIQ2SW8Q6sneSDPIhcxbR9Lk5Y/egw
IMQKv+QqF6Tm+6SzZ3rp32ppbrCC27kb8MDY0TrjC9RB4f/hzyj6RjJRNPEAn3szM5myY5m57nuk
fMxZzPFWVW1uM00UjSh0kSe5Ccg0QUAsXcag7jqau7eenRJx9T3DtySvKWcrt74H3vckvLC+upoL
+e4J8UnPbv1MpCi4iLM5JDPypZYKe1eg54cavXpXVqN+0J2suwmnAPQ76FJP0vJNB7rW873Bf3Wi
3/EnRs1frphL3FQaULguR6wF+/FbWf2Yjj5uZowoOePs7sLkRq93p1868Id89brxGy/ALsN2tal4
/xenZzMNWy+3MiF51KlBOsU0tHyItfkThWcKxxYBi12zNzZW0HXZhTXpN+cBUgbr+dKr8+508HbU
90dm6YrVO36OG5w/AXXVJhbp2HoYtUlFiluodHFgsa2wKe0loV9VWHEbdHS7yoJPO6oi1uZ5JNGb
gW/yBUfsppBau+/JTvADPbqb1Af5mRke3hbpaFfLMOM4qeyqlC1aZjT9BeIdif0notO5zrmgjYIH
EkWURFxA3yVM2DLk4mZPeHQTshXTIblOe1eQ0VCLfy+9+RgngiS/FgghyXvDKVcU3l9x05BTKqiP
OR5/+Jqqhc5KnknRJqHzKbSLawU4s7dgrqNZNNdc1PRQ9e8PYW7myaBb+uENH93BGGKg4rTbrXy6
XIX0ATPA2iGbGHUuRXhJJ9lvnlIjws9LcoSnjVfg58q/Zi6ObMODwQEBjy93Nw1VvX2j0anFnH9+
QEzLC7O7UXjc7FZu6goN/XcaJnXb41V0kbAcAE6YgJOCFTXBqpbM8ebI/Rki0lUV+iIW01+rv0P6
syuFEp+2RQ5aCP+7imhoXOEGg7jULPlHrm2xfgsp4NpByL6RIGK3AoRRFHmkCbXKSWvemHaF7yVR
2uDIqhWGUFBMNsXsEQ456cHMmzligX/ttbIFbdf9+L2Lns0ViaGf85vf7q1uwFFaCupMsQgb2E60
yzQahMCPPNzvECsO0UNXPPrFNjbnsEN0mn5OvjBsE1EsO+myL0uNdpyQMxDm3HJ+NslLx2SEnOAn
4yFTvXWURaPyyauLIWetCvQ9RB4C1omeDiBfxAcu1BHo1vtnWbAVIpztpaXnF0c4jlDWgpI4+JnV
3nIMugRMQZxMz/7oLzrow6/rZzt3ysUW80L5BcS9q0uOWWGBEidiDUNdIfsOcSDO4LcavYOCguI6
oqdmBSQLB+eMXfK6L4O1gFDpwrC3QMR+ycy7EBRphAb2+ha25SfHQxMUxGugoS3fCG7PCJl1wVfc
T0pEGbReJKVVdTLjpAIlUuaO63+OtXnZLFygy7FGkQg8Wmuw5iPfnrZuFkBOCx28Li2I9oKVuG8R
jO0SX26QqNcUDRi1twYj+oiEP4AVUgSZmtv9z9CT/54W8Kta/56MWpDknLaOJI3h7vfxuMFaL+Xz
i1LhlZd3Tqq4xeunzLGLt4cPo3+3rKZP7NXuZPcMI3MMJm23MpzNakobaFN0TzcfVt//SeybcEzs
pEerBem69eGUuDUFB+H0RQDDfsYSiUZrWC+uoBabY/yFq0zQ5vs+bdHeXyn9ZwXt0D3H2grjvuAH
rW5l6kz4lBrAl1sULmeTg8ZOL50BMo5h5X84v39WCGhEsddWADPhp7fhesHDsrqBv5p9ES05QCgf
xe1CSA7m08JqzG68xfjK2ni1AhEYK0CjOtr7vEE7S21oFSbH1LTF1ng0nyqM4Oe9mqQztLEhSQn1
UyXHxQo/dUG6VopkUOu1KQC+AFYspAT4mMX7HFHxYXn83GU/QYQCI96vhEGRM7tahcBZqAd2zFBS
tU64lQ6sISTxswfty5+nroWar2XXPy3B82G/5a6BbCOVeFaHUZPm09WN+V4kGH97S5f02O0OQwSd
U9ObaBGjjHAoMCCiYLcB4Fck9Z4vHsGUNpsGOeB8MlJSm/VVMMQMaKIeZF15Bbj+eP7Dgma4cl2O
WtrbwwNdkNVkvbBdGUx/ZTeF6nKO3o+E1+3mSszO4AYx2kuh8wGwTtwWfgobQI5QoALFW/xDRNz8
fjbPKae9Z0jfdXetNVVgP9IRBr0Xhss0Qk6N//2W/lx8dCCC8K7T5j5ra4oDz7z9jOhqSeXAqTGL
DcAGI3t4dG5NM+1ex90dKYzd7Z+lGrkkYr7gNozO6P5KClvq8PsJV0ryobDBH9omAWefTLDRDIP0
WUg197qmMAmXc5+cC1cpt/k/4f/qkevYnEz798p9UWuk/8Clq61R1NxZWhZVT0TIYsOyLs6yd2W4
/6/ioIcAPM14GAMRYYXLeK8TgjUWurqWnlUH/QN6Z8w0mYNik323X1j0ZeWqZeeTFkfCIJSXmlMQ
HQkSqssFYtyCZ+xn4djTM/LXG8T1orFwYzpUTCT8aIFlpevDiD0Wxx1VkW8l3NV/Y9PNiLxx6C/W
dFAJl9tJ0J7nl1ajcfJDscXeI0IJU8vec14rMdjhmj3TO8YKlr+SVyAwQ5tHRB7HymUIxZWmmNk9
vbC4jF26ZRyv6D0VTPMjrKetrcK8gpAO4RqVeWSoHtoZEKKbpbgUad6VLrbTq4f34GQLEj2ht1dB
mBRgWIbQZ1ZWb5l3NRYohYbYfuDRIUBtgKllKJxZxJPXs6e7NspvJ9cNpCi1M0X/erSBUSp54zpL
zQTYTqEeeiNgD0N3LhhmiND6avpNBnKhpz7dbP/4yKBcS1u+GcOXjfOoQsZZQiBYlc39uUDXVvA8
cyvdAeJUuCpZyUecUK3Ng31jstvlWxr7fIk2447jBSUXbI+njzPNpzSx6THOZAKc4PwKnJOJl8PS
ftoBvd0jw883I0qqBYyCkdMKx7N8IWVkmU0KWHf66kyUEqSxyBWd+A4yj6TC5ppI2B9x7n+qGPBZ
OZwZbfFUIOOsdFOYkcAwV3RZ/JGD0F9kNvdEgd6q5d+dP34KY9m++VhgQbw8i3zjVpjNLmFpiqC+
ZIu+X2Atg/vJsx2v7olGQytZ9QozId41C1TeobSRo41x/4xXhPto21bYDYBqA+xkww0UUh1kGHrZ
vlwf1uh5AUnt/SJ6RvF3zC7EPkbkhSrbQ5uYG29WrZ4GbpmCY5CGGCz/z71Rwoc08ZYQZcZ1Syjw
rpHe+ezWgX7047IPRM77q20/jHBalIy4RKTJhZ9JGLRCeOapAqF9mmpmRcg7cpkiPyK3a6L9z+fb
bVGuIHWxQuTA1D1jKjrImd644oVC1QuD2eMOiuECYo9zGH3frM9FClKm+G3QPuRCJ/5r1Rt3tiQ5
3A9LWhUsBzppITWVhBipnnLMWFaX+0/t4FW0POFny+e25KVFdXI46eiS8eW7QnfwvBUJc+4hjYg+
RmeEuy/UyHrDtcTSGAIuBuWr8bsbrDemJCVVbNQCBBesaQu3GOv0DC5v6FlrDXljMYAMH+zqjYxz
W4cccKgHXJYCmQbhdj8vfXAQ0zrw4YMTHx2xYfeyxocQ0uGOGi7Q8N1m4X4THkxmdCFhD6xBbmpa
3ZLSp8ScP33WxmDm/cpCeLvvg6iQ5/q6o3cy4PgRF617uHA4CZL16DVSeUCZ9Q7j8YzJUqquuzvY
7vKaheaIGt1GYkZndfiN5zZixhamNn9SIFpiwNJvdN3KiorhBiPIS2ywdkOvaNr5Qr6qiATuN/Mk
Ijkw6yTA80XGQd33NxDIhRSIvxxxrZJuqqhwldcQadPQQ9WQZ/If922J3rcrztJdr1PirwAAlZFt
TyKCC++i1BHrP7gtFKNPnXiM/Vokb4NE/rhMBZ877UHQBTzeuqnEVlVUD4lOLmNf2wRxsW+h85vg
n6TV8RxCDFjk0umUkUtlqN2nd8uMCfBTAMV3ha/T3aT1hdOh0DlbIpoXcLp8nhjbXjz63u1x0RSP
ds2VU92Jt/pYBZHWCKpTiBV3OgoDabf2rH1byNKy3nG4ILk9210Hbl/DnmmwfpiOPDqHNdtv5nNj
ENRb6H0st/B7oZhsGkOdct00MHiuaXjxGFBBDxChsOdB22+zcG/BuwzV0Jwl0gwibol7wQFnHY/Q
blky4Ey0I9zvkjTSIua4ez+hc4ezTrJ7z0GXCYl6kgLjbYqqcZC/z3dXGd+O9KXT9eTnKh92xRRP
ydfSJZ+bIGaC1iNnDDuIsiyZ3QDTJl6eV2huhEE1hId8csCRX2D/3ycfMQlj60zLhCBcNMryxQG6
l6JgFVAKXrM7NAjIUhe07JDpfSwtAHWBoymuZB5AIdzcsBKkYjTEGIFQxA+D/rP2kADXg3/DGAhx
CpSNArgAZzG7KJRXNEeGSRKT7ZQlMRCZttWlwolb8MQoD9ZGyC8f7dmjGmEfG+HXHKzhv/ktP5dd
O1hiDT0cqHWIkaKC1PA+tVUa0AQWGe5GEdrC+wvVe8FvvBETtm+mznjyR13u+PuQ+ldtBkTgSUAo
Yu+S6YoO6a1X/XWSOhvteANXp4gIyK8T/IZVKpLC08MnwQlLwVCdsKwwOUWR+W0WdtbDX4EDVCz1
yVY0bswdKOVj/auepYA6m8TIwKZhvlG1K94mMfHdc5M4rjdu46w72PAYAB6PNSNQQlfXzHY8KzGH
evQduWEq+LmP8N1xeRTA1cxAKd4eqX0xL27c14i8p8L26PkFW5z9cbf8bJjXgh2lR8d2RON0xvbj
L1jAxq6BZDLL+aBjUQjjzOUAdnBXJWZ1Klb0bruCBmxAJBN4VNiUXwrpnGU4GVVfNPEtyzLm/eDw
nniLQWp6tog41hVqICQyMd4SR2+gQst0gei45MSpV7Fi4RXPeiUcXyP7WpGUfMh+5Odtq1tRYzDt
X98r6O5UUt1IMYsIN/k2vjrOI62EAgCnA57HnJYVuiBvU7mapsmRdEcsW6xwtL6vkFpQ0FBd+Ptw
zdidt+wsYwy0w/H9fhAVundsGlN1DUuDUfG9KatLfxe04r1gYBmO0D+IWyxDVbTSxVqlQMvnBkSK
Bbu8u1Jkm6jZQbyukUbNp9L0UwdNxATrUc5ehvLPGNbR3bLTZy/3Lb2h9SccfSp4lOOpniCOXiFf
65Gqm3jvn7ibOrLw/BqNK8GN7UsOPrDSUkwdHNavEtDWn/7XHVPvBeqhIDGg8wma6XS5D+ouBWeg
QMHz2OebDqAHqgY81JR3G20YJZtAdPEpxJJkQWEoivolnRo9lqKoUO3JwXeO2IeQW/ttAt1Jn8MG
k2TuY9+2PIHXJmeWTvYXYtSBAyoP0nqlT0wi+eOH6hsviCDHR7M9u6dGNtgX2P0PvJb480ZBxGDD
1Q/XWHqk0ybnE+7fbiLTjq5X4LgUbFOmXGsLy+z86QFAw+VDkEdlfJriavhADHgdZHuL8pW82blm
+DJSB66c2aq8nV8X6aRfWEZOW4fYGJIRcdOQO0GFOqRgnscAfHblPTPEWLnvJFrw+ouSL8M1IGLp
e1jyELONXNnSBUB765ZCVYVC4qH1BkEdH8uDw1dQdrR6AsavkpomB+QSNDkfEkkIeKHIEKSRDJRt
tgwQ8Pt67CiXh6gcwWl+IQAx6laCT0id5vdXyKU47ysjMVT3ScuMCjkHkN3pdSOtp31wm7e5JDp8
y6Tsa2RN0Mu0iz1WcT/iWacVBUMLvljEilVdoMaXtkCDC9CKs1g2s+/jq/rLK5/scoHnQCSfkEJU
I8lJa8InaMz4d+TsqCtDsrhWHfXaMe+vLZ/oEnvnsQrOKO3c0FFlbDRiaHfnfKdg9iKVy82xQwk1
Yowl+a/esI2SLrNGqCztbglWEBoZHUoPfE6qOdtqS5D2rsVJd+B1Yx6VQ7TilL6irTAtmPLnaXk5
UkqDXRiwY2CmfcAbIt77R0tL5sUiXNDjYrP5bgdZn8brAeZyDoBnhfhTmBq+whdLqSKx18TMVH42
NPn41SaSYynnoKQt7AY1ad9VdmmNXo/K401t9xR+enVxmDg3sjd0J434pQ+ih4tWdzKM1a9lYdFg
4u9LnPNrn7+0QHlOytpDOkZSRJ5R1KB5wkNIRPaKhw/FXArVJf7tbF7fvEgVt6Wr0mcjlxq3l+uq
9AiP21k9iph9HwprQs8/smgx2ZTLbmYr48ZPH7+eUs+6VFvBUmtiiVOO74sqm6Oc3h2IoE0CU7vn
RFDWldi91jxlRTqDQr/m69GCHxoF+n9YH/JhPAojJEKHYuG4iqWO9gDNL/CPrl6L33wYiMTmiSOT
F7hNzGpFctHUuoG9cvN6/X/ClhossdcNTuGAOAWLm1OFFUHFmJTF40PSogcWTR9kaMKOjn7Rc1vn
15DRr51o4W4dhcmVT28sN1HdQd1zafHI9KZE7yYo2BFscOSKy1ASWUMPbmFUC3pVHRvVIcnp7eEw
3M99DjzqbRSR5nEEj5ks887HQTfoJDu32Ct5dt2ioUknnlCcwf974P/1Sg7YeeF1DQOklIMaIWAQ
mCj0aOWPCOL8TOT8oDlUsIS/I74VNKIPYCNlDzGYwbRn0SCnTQz/1TDRoa+FlyyzDTyxNKKxXquD
Yf5pPCOxE+ABEbkMgNk5hVS6ykpJ10O+SXMQdiQtloNziKlapj+zrE102Z5WcbOjTtvtW6ysFT+d
Yyd+ipnDTLgd5QwIc6l9ULTeZM8sz/iSwhjS1hzgq/XYTrDeQZMVpQHN91Yibo4lyI1ZSWNN8rNe
w1acLlvcH+oda3syNkMgkNjMJY1eSJuFmd+/ZhaHrsaOH1F0a1d57ZoDPhaOXSqSOXwLmA171mF1
5tdIFMEzrxOSSCBokqGO87jS9dPc/c8jVF5PHjyU4WyLGzD9Vbv2PJNBwuxG8aB50g+rFqMQ/mJO
WouXsGiK25LlngXLoz3DsC2olJnUV1suWyoPMBMN8p5kmEOu7mCbfNyw+Q8OA8Y0TmaF32CA8fgB
/QGN84PSZtUCt8GxLziNgUK3NvxXc3apuk23j05RpcXZV36A03iubRj0jIra3Vk3t68xXW2+ers0
zlXl+CBbKVTfoszyfQ1Fpflv9fvo9sTyp3t2SUgY+9LZIU4onaBXRndHr8PC2fgozSQGJSDORcZ/
gdVXTnPrHEd1FFlxIR57xynsk1y8p9zgZqDWQXXdW3zCvwy+hgX05z3p0bpJM5p6XW2bCGr5gI0P
DwNCt31qHsOVd9h10Noi3UyPWlipyRqgumCAs01dv49+0QHglgA5nCMy24SzISPxTCzT7fJKCMJ+
N/BSYJAK+GrLPWw5N1hG14NebqFiqQMcewQxZwzEsofJdKA2vuT1dI4zZr+4U0+b9E1lfy1qiniU
8tcY8sis8vp/FvKA/ou20V0J+lOAObv+/wgMET9ESXF0fJ42oejltszWoh4/ECEG3KRi/Y2R6EXn
8+EkCZidI44NcU25tMUBHMPzryRo8ksoejdP2uv3X9sz/Thw4J93aKB66mWRRAijhTu6tqAgjC/D
1sZIKOXARpGgNdAlSWNWlooAxj6BV4P5oSnMo7i3audFCGsX/VnlAC984bbfWzUe6wcH581095qa
UM5a0WtKSlcVhkQHwUjV7aCJiX9ETDe1UwRwzfBm40zlz6/8pwkbHFwnX3zjMYkOewtTXFaCgHy6
ls6/YHAk/d3/Dz3xxAX5ZJZ+F5k3NrUNXr43DzbWDJrxI1pmOAkMzDUl/1KYhQLlh4X/DYRucLjB
oW8lGx3/y0G7XhnvlysEjLbdLcScCsdbT3gRYKIETD3dMJ/47yUCYwp0xOiixwSFQDy5Tnm7zRf9
uo6XIOqxux25VOG8bKD/JQ0Vo8mZ5tqCrakzl7hmUG5ZRVTJM15FzKu6amG1yBR1yWaB3WTW4AuW
wmrEcxbMm1viVhPrgZtXBNV3kzFqHCZ5Jrh63XnwogGyflKlcHwRc9IOBvgEgO8QeB24B2nhAot3
JLXwJqVySIXgiB+YoBKbMXvQKOKJv+S9c//7B9sBm2LWVVYtr3rrSd6enCGLGNOecLf4LNtF5kJ9
f011QQSqBRURHucOFcZN5n8xtr/0zxc5OSgjF6HyoEhKxJnZ/lTs2+Npf+7ClHC7GWvsxvQHVVFL
MwBvHVrdDHxAPFdCA+R0IcyzWxD7cLtKTnuwbv6QXvE95O9pp/WjjUzG1V9L/7IadfcagDGLfzpM
4OXZmdsY0qsYYDh8UXo4+b5SZbgCG3bYQpokgXNK9AYrq5mAnej/bL6bg26iE5zROX8ibx+d2GnB
o+TtdnJOQi9gUr+L/wAi0BwsgLGE+ozYWk0264InLbOSzVznuq4WlhhaWrbiNaURaMltgN46l/2u
dC1zveq/SU6L8h+3iq7VJ195HmpOd+siY9rY73UoAov5tSSjN47XdIYTJKmD+xsS82FpSNmRYT+K
u6oDJgs7ppnQZSuJp2xyRnJfsoNOnDxuZ3aHZfMe6vvFQnx6vq/cV8KsFBYwGdvpPGm19Y2bYJOa
2yh3wt+972rH956mtbvh3zA2tuhN+WSLwwOxhYAt8XCRvhoEF4XB2RvDuMJUxaz5q0aHkg7jNf03
mhw4AeI8J46Pz2Oh9+3D4Mr+jdBv+SRrIvAr0rhLbAgRnrjnFSCsvqLSi5rbkvdThkr6OwWs7KfB
nK60abzpVd7tPr29M6ARi2ljYOXvowsDT2IzbOxRPJ1T9QCQQL36A7TUxCbXKPfPzhLAwdoLLaFW
6GeSZmWFHtX3arv3zPNetxAEThdkWVt9GIDh4sE6jBaCF0Bg9G0ihNF4TiaI9K9ectUMh82O/Cp1
XGcpQPbzczFcY6fn1vqiVo08ORLyTXGqg8HHvks7MUlv8M9BfnFFxnTCnQuaRRwnkymxZ1uJrxhj
2dQhYb6I8wGnITqUAShfi8BJV/DZR5HdSP/dIikngvUzQDoBHHlaEar2+sM9uxiVcdz1j0Lt5ASc
f9DrQ4k8uVCWbSRdic8ZH/Dzj7tvTYRTW5gRXXFDa1lOLFKQeKtL8O2695QziASpmQUFRADrtDKs
lT0IWWreuqqqEGq86oblAB+SnMrM1Bdt4pkG83aFmZrfQdcMKgXRf34VW0hzja0WrMKLNXwqVX5U
p5oMetjF4jZ+aYYt+GIvUPXVvsY/JU090dtYO8Q9Buw57JkrEpwNS63mv0cBjLmMpDLEXDfCahY+
BHWVl7eJC0x44ES0xCyg1HsYu1JPMCs4RWl2BgwXQF2WTj0dbALdFqx9S3hfk27B7bQwA92gBXLq
0XKI2woBbNPhyKnqjFaXk1SaiMEX7J/mdGNIEjPFEeSlmbTpmjA9pLpk8sD2nmrIa6sif/KA66Eg
HsSbG/9SticHC8zsAnkEhnUHzg5B1pYf+/+4LUJGwSQ0xxB6tdKrGTiujXG86w4aYU99RvIKR1IV
fSIkIB0ciqfXX7F0kgS0ijEqbDnHqCLf7uiMqpNz9Ug9KH0dX6R8qUpt2+bGfBCOR0NVrekzQZge
CLwU/lUe8VhVh/gZbW69PS0lbVfgNu5YhXN4xVLYz3AnynwJNII1XHVxNmUBVjM8L6BwVPwg+aSk
H1aRvWue7sHAEZurBfsiiiB2wjMxMKfgFOHSbo8ptsq05/xsk9STsRmhIyGdQ2/Iyapx+6maGmJB
S2D8Dy1Fh+kKt6VmnlXlrpv/vkZrsnXZu/37ph+hZbcQvXKleSYhxJ3wv4EyRE9AByXBC9XONkFF
/QLy1EaCSlNygkdzxg/It0oWqN0DHpPNn6caxGTGC72xTFyncwDfDyRG1smmaOsz8Fy/p2C/3XvC
d94Iz5yEiAYzb+BnqNFxTnEpemhYqYh2XZcPYa3RjtKdclf/8xDBzfzq/myNTg18SqNCJBmYrasO
988f0Cdvh1PMgNkWjv7EOCcdZ/Vk63iFfT+PhbOxfejkV0Q9hjcPpHaq8iPEbuDAOxcwS1rWOJgi
2qV41u94uwQ7QW1wlOtMh6mzKEKv1QCfRvXVUdSgEYGNMRnNv/go1RwRo2mPBmnSr6geWQsmcEuQ
p/O+U3HP5xnT5PQHV5wgnNBvpqeFMZ+jPXWF2NDct6H/6OusN8A/wjp8zaReYvPztGvBp95fOfaN
LhWzuRwmr8RDoNU0rhRjnFXBKZ2xilc+eeujKKCaoWfnyNhUEDtZPtbspfQzNTGvBr00hMmwLWhR
u+99h/nhS2oy6YlEXfzeN+5mSPGGXqQcUcxvVM2VoT8brYVkpqcNsdRkM07kN6DyFglgr6NP8T3G
SIrhn4mA3IuiIv0i9CkCmyYewT/Bbdka+XfejNsSvEMqVUVtHeg0mU/bdY6GoiR0bl0odp58KOdx
sN3+o+GEIOcpaMwRQbcUPdXe/A9IpB3hZP5Zf3H3bOS7tDbKgvrNF2jM/68o1t+LG7Ja8dbKIa1t
ZxieJ7ivLwH33xxebZUmkL8/UYH5iHZaWUIoZQ5njaiz4+Af6uImsJh9wcUuTWHDYUWrcvfZJO3v
UlNgKBZcDc6lRY7Md3MNNyWCgMirNwbw3S/iNmM0ez1EuGOSmyr9PxAk4WWEdbcCB7S49pBIOPHe
PBni1MS8M/APRfC53uj6C8BQohehYr1f/HjOwuj8nh/024PSvZmr6u+aNygq0xg408to8/SoUpxu
Agqo0tmolqR5PxElQOCidrhBX19VMYZANL9HEh72/+9dUoclOwWSn9yWVT3QfXLZ8uFowANUxsOJ
5ben/egF4CurSgNfEKIrzjx49Rq6FgHYE9z7q0yRDeE/4LOt9xVwrrLyYXCb4xw93/QxwtnkWqLc
LbZCYbpV2LCKue5oKVifLLu2QQ9wuMpx/lV2iSx5YMwLq/cDGrX9ppne6c1fml/t3Qf8AEizgFMa
XKMGYrExarpdGwUzA5KMpiUyupoxyCrXc0cQcH0e7cxg5wn7/LwPE88RFPqTwJ6+5p8e69tEvo6d
wLC4b+U1BI2NVf80QWWWhXZPCG4/WJe//e8IhctnFgk2XtriJ/WBV2jjRwto/TFfJEdXPJiC0kSu
TWU/CGq5MZn/iO/YtgWvrKSx6Ye5y/wwR1rsnDoSxHGCBeyO3uFvDUgDZ6fSJ8CqO0T5WueYD246
Be1AMhIELQz8Z5XSIn0Hd/tzq3pmMgxI+hXi7rIn7WsnV875EqPK+ihNwlvS26RN5sLIUQt2B8qf
ZaO/LHxgnrZPxm6tleGuVwNzBgP7Gx3l4qs0I7PBBNuUIGMDawlNKa1OwJgr8V71BzUzYuR2OcpV
AGigy2LHHYKaKL11ge9txpP0Kjhuz2pbv8EuBUwih/B9OzPEe6N7+JcmtsmQF5Yw3GY0RAy4ibQI
nAsHKH4oPc5YFrvZbNGgJwO/TVRp4VehVXyfyU0cnYLBqhiHtzWetODUqeyi+7tr0KZ1rJ3x/sOv
Wmf6FXkRZHHPW4UzXJERoB0PE99TGp/sufdu4fN4IMeFPO0UAQAvq8gtSoAAEv7TNb7dHfdHnaXa
7zXF9rb/96LFJCC/fo+2sO/HQJMOpkt6rhWGY1i5jTpIa5r3s8BPJLm8d/+bv4HkGJN9b5sbK9QU
mzggHe6pTMXXicaB+fGl3Ky9c9yrTSL1l6WRNlSTHBnX386/5nCbSiR5Bg7nnF3Sq9QFVs6LfhI5
6PMLGNthd0amQRr6Gc6bbotgmrY+ePKu4OwdjU8Wgr+YZaHVXk9TkFANx42/+3Br75t4xZrmWmsP
0ozU7Kl6ByPveA69bONl9Zg3LVcqJtoBI8V8IVWg+NAuhsdpR4O2LYDHP5ZYDwbEWfZc9I3qlsIo
dRex0sNkeT5+z6ou7LMDYE02VDO9ZLEtJSqKGgw023rJ1q9Z5sySdI85Uy3XOZ99VIhW6S03RZKB
7GnlrnsNnryuof9JX7Px0AseGP2RIVuOKKOZlP3KSsBTJPEHQUj4oSh8M2NnceuMNhllJ0qkU0bI
CMOl0vgE5N5QD7Bmh6tg1h2Ek6aV6ubnCWEK3ofRtJp5M+lngeI1bwNs0PPaVYnoyc4t9zyStOka
bhFxq5LLVG/PfkMyD14nq1W2FCIRpzxPFOpTwWa4NpP9U5nQnbWQfa97PdEcBN0slsNAdfbPhe5F
38droS5ilqc2Vz92OFWUCq+5ecNRQ/QwPkH1bk+hgBEN4OuIFDmbeEvWat58ac41bEk+IVZV2v8x
/axS6pLrAsuq1V8AtvSvfSGu899VFbvf8injx+tGC0/6ofr5ztSM3cMu6a5F+f+MxfP4w0VT3V62
3ErOXY2SoIzGmXQGbZyM82VqZ4EIDuU35kBgQbRCUtVaNAhtehlcXCCzWsXwvoCmdgrK55RRItLF
WnnMxjZmnr1blwBIvGmOYdzckyu3lg5kspvitJOBjJUSFe/vV/tLHjBSIc2SJGD7Upy5eefRFqQC
NVZvP9Pidmlq6EcdSf/kRDvzGK2graOwD7FpGEiMqsXzBGrDvqLlhRhy1eU/2jVCFhIRVOcXhVLy
RY4L+9J0HFStA6Wx3mXTyMhnGYghxS/OcZaIcGVe1NnL/CYPUfhtqYpa48Rblzx7wCl145hI1gom
32lT3jiBxS55U52d4PslaXZKb6NcF4dRgSW3QV1HA7NI5VsZy1WoodYXhurDuSaNtYMlxD5wTv92
F1TkD4WESq6qDOpXjwcoIyogX0KQlT0H2KNoc9Z2Pym53mafNIfG6Q3E4TBtwXUuoe2NK2uL/yJC
hbIPpT0A+uz8Jonwq0kUmmwZsknYRQpKYL5MM/9eWwQhyAmJ1A0v2jXNiha+btQ4yxYnxxyJaKv5
cE8o/TADWbDH5EQZj4F+Ovm0MewsAnjBHjzs86AkRlhACr50Z2kiSFuYPS1GE+81A+yl7Xz8z9aK
0OpISFHNIAjGCOhN086InzCJgOjClCuAVf3/bh94hLc5ali8FaBX3r7aYdBsgwmg+8iH1bHr7M4y
Nvfq+UJFP0JostFX9zyNE3L+rbAxKe9JpVqmqYqSzuE5LLnIQ8MjqPqk3WBoCDO3srIwYyk9m4Pe
I+YNqomr08LViMMhUhaAxg0FodnyrFyFUpI9cbHbCyWkGyPPqt/dq6908cXJq+d9UOdMOARdZ1yp
HUcEZYsEW19itLSBSJ3+6UcM4Z2Teziv7wGAeQ5bkRLg+qb0CaGwwgKzPxI/HHCS9/5OAW2HwLcd
7P8BDu28IzJW58kFETOEMaw0dKdrillB94/LJD5/XCaeZ+A9UlcOxXjILcPRg2DJYngZarkjdEc6
6X9fZul4s0RXcKQOI5Wv/U8V4OSWQRRPqXMX+lxQ4YFyTYn6gya1tX9TmLiVe7PRMCUYcdj71Wbz
qgfyEmQn+6ExJbNFA8WlCVk08D/s6DK8uzJUP0ayiTh8X1hZ7+Ebumuz/bDyiqmdCST4geAK9XLu
8waDVFDip9IQ+A9qTxQmIzuoXW2hlLEeuBmb3+ehPaGBj/CWgnfaCJO7ABGl2ykO0Uto9MCedt15
oODbsESs16n1QE2hPKhD32Ky+Crz5raVdiioCjHQbdxbGaGdmtI3U3GuBtfZGdSmDesmDKsUpsgV
eWRDHQlxcDtwZmCaM0IfZJ5q/w2Gw2KyisXBwFlROrrnmNCz1vQFsF5U+OzTNqdcEvMPmuKjKj0J
1xQmiMf03uXSfridM+c7/TjbEpOIal+gnoTtb0cYj8ieGTGOGAnElDpg2ENXjtAtQktYt7s4mn0d
DGRqdEpllr4NcSkGNaGMF06jEA81S+2Rg/VTp1DxuHkJOjMCA10bOLwG+xHSj+EKN96jYfG98Tby
yPYEMqr9sdc0yFiN/u6hKUaOdRaWnsSRODKGtYhon0HaESjuXEMsYLvcmTdY2YiJ2KFYrcyyCfQ8
LFx+ipvLFeq+q5IyoYpJcH2fRr3tVKHZe9n5gNN1BbRgOHco4S0EFSz6tChNvhiXUsxdkx1GQhIh
MThNllyOU8xgY/lOKCbZ8Lp6Qs9rt7jvhzCYwQe+SHWX7DezEBAB9AVR2PpXkuJ9bBxJGpaX/ylX
Y5Ww3CFo5LMldx4qGxaqjoew2z3QA7SkUopSZweqRmR10TNZz2JH7ax18EjBRVIo435EOktvoHZ+
+1ejGNf2lwwqLeXCKv+PPqo0TSwrZb/NPXvAy0q0usnUh5NfTVQ496Zt7Byn/r7ldL0wgZmLxzo+
ghNfmKMXT6wI49OyZZksrObWjT5XA4slwjjmAcqw7tsxNPrud59/E8/eWuzH4Nb8sPdlrwaFGMGa
apGJ7vdfbmy+zIsi0k1M0WqjcRNHokcDgx2JuHUymS7r+AfyKyp08rIt7X1Y+ukBTf+sDinkdZ/x
AzJrmwAxD+ZITpfesSKqc82HA2EkB9C1fHjE2osenU/DxPcA/hfFWbp0+yFiHz47TwiCwQju9QC9
UPNNET7Z+kYzok10LFZSgzZTlQp2m1XPOxJBUZFHx7smNPp1ce9Oym+Pr2Av6BVgEbLlQtrz2mrg
oRWlml0gf/TL6yvO5w6KarKDfUq/LyX4q9YYF9Vkj7ri8vvgYkeKVRBs4vrHMvOSE5HnFoPUE64n
pD/Sl8m6PWoYpjrLQuQyr+7m/RofSfJdZGGQd5q8NKj+Q29uwncd6eP49Ftoi0oTWyFgygk+oa3M
ZM2+xl9oj3/9WZpvOZxByQ0F3d+pKb6cL2p39X+mXOIKRjwZ/ddA9GUSXf0rj+AE+/6MzlR2lS8r
bN6/1tn399EVnx1csr4f++k01LOcGhh0nw4/wZNGR9SnmnOA3eTRjX5SHvA0c1Y2TETSIvKRQnXo
F0cjRTX6UfPhAkmYO8SVvxKjhQW0i86nYYVudDq2EN8R7vuS4M1yz+xyrYFEm/3bk9XzVUpxJSmK
l48co4WwUU8Y2WFpcIfloEpsPrGGYzUOE0bXwsbxdiLgbqV/24CXBevRWVeU1KL09amHndhwWfxR
svKDcR8KyE9YqZk8wWBt9z83mWpnQMNzW+FO6edsiD4dkkyyHu27WXzalWZXCexL/mHEcYYAi/Ua
Ggr2SiolCQFn94B5p/qraPmGCJY27kaIXQnsk35xeW+ltKuo741PPyo7ob3lRfN+dwT2yMicHUc3
5NsZxs6D7NTnii5wXmm3oNTvCtGdPJ1WqgqQx01K05O5nOuMlaREj7HjyPOSBTog1hUMOupauP+l
TdrMlj5R0Y5Hvi9yZD23DNcyTdZ0fxtZWcttuidZT190puR6rgP9d+CfsqR8E8uhOXyCAb2Cn2mU
5BmAxJWBT0mmCi4eFmB6TdEOkbE2+QruS/AGPsc94ynBCAiEDfE1bPKreRdJ5ASr8pyvAzc83OER
WVe8Ss5UP0egEh/MpTJwA+rvNksCCe8q61xH+Te5vJUqj+vLxP6xeiTH92g5unfsvyISxOe8d53A
Yh3zytfw1KNtNMjUXXw7mUGdTQUBn483LZBRI9UFr3l0sOS7Iqr3ItUUI0S4zspNFK550ZcZAeue
MdXBoqkPVWB/y3IcPh6ckg1NpscOSxN0mCpZw3Qhq7mcFqsSna+WhYPFNsqKiD5i9t1ypyg+QQlK
cmu5zkogsiRClNNETb0thVQ8nuzI0RWCIUI97j1b5K3jTrVKgPYTkQj63DntzB454ej0aWe8SuEr
g+oOflwTlB+DEM3JnG7LDq7yU1TZxAvc9dBJr9YFdzN1wx0lTBjofesZx0+9nyeiluuS0XfDVH2n
p5DnA+CgmlfHjA4cVo49of8DaCkk8lM+dHIZuDxMlRGwtSVGNOiiOqaYqrLIXnjv2Yy8Y4hE+U8+
XkFSD0SNxs28ldDutaCiHPIe6ypKAl3OnoyJ2/aaugGxhL8o22hZzVXAL7mQD2hQwwKpl62HF3A/
xg2qYq6v3QUPBWjJbiWggcQROqDKLy9Qa9IL1/8SdeUqwAyUxBoREW/pnqPxcxoyN/aiWvCe2vzA
gQiSI1AVbMp4m9EHrxNdfcsLEPUhkeEajR5HBPGKxh/PxkM3wkvTWY+euPR/ZWaRkn/8C9cQ294W
9Jh+zH9WodA2EohSup895c7W3osTXk1jdJjBJowDifI99eXId4P/Y2eb4A6I7kcbj39WXHXSig3w
egbA5pFWL+iuqAuHvHOajreRhekTvPeJZDFtJUOLrv0O2KMpM1DKrplGtq2j3YBG55NpaDeXDC/Y
dPb7wJADmMVMP+Sp0lZjxzfrlan2Mk2NZo4sRiRZ8aQStzBYMtN9GT/pIyzOIAtosC3d4gUV1GJk
9Xf6z4y8m/eoZWBslVum7pJtr0NyMN6iccqg8pKb4fjFBxMZkP2SeAJc3kO3L5bo32A36R0geFhE
9uPiwYl1/JVLx14CYWGuRV6PkDhQCNaZxWZVVOfuMYZw2rRFThAx4YGpfioZw+/mXT4NOnC8/bWw
m7kirgeI8inyqp5uCwDkX7Evu1b1sEHGN3ZSTJlWpfzG1/WpnuZEjGqoQXgs1b50JLF3TfuE+8mp
FKdGYfyyPyynuJUPrM4GIo9i9tzy/aPGgBgSbf4IW4VxzUlQiJKVdF00VkX47+a0xLM5mFNtZA4J
aA+3dLEpySE4uPlCd96vemJYcAb1I0zzooZlhYjPJm27ehjb/ctKNU/wSGqu4n/EB9QCIn2lJeg3
l1dpKPDipujx3PMUhwTLD+m/TdVMuerk29Mn4pwcIQEXdJJn2v6+HzAhJ7DLBSl/LfaJ9PQ3+Ln3
CJU2NUThGZBjoBD2lRKCIJgQzUQPTeNP5K29XtLOxqJGKbsPq4cmslnzQp+d93vyweXAq/+U5jeS
/bmwnPbUp4PBtEIK3haFAlu2pfweaIUdMRwfuXzwbsWdpvWIXKPxJQ3WGaJ80h+FHI4S60c0GIdA
5eD5hqBZ1FFBT09xjG+iLfVW0n4Zgn/z9aJXAYW0vfFYIxmGr6YHfpzQ9sPQJclg3YxjxclwRdf2
wwch2qt7r8KQcSNBFDvvFdQH09c3kppcktK3b/aculUrQ3VKrrVucQMOvpawiIQXEjkYe5oSSWSu
goyy3F0jH886tiE2AB7L6ivrUrtlwSbmg0ZqLfaFwgH9JW8lLtaTaqU4llBSOgPDrUKb58tpYSAi
PoYGT5XO/BYpxNtppNeHqcFG9gqfBxjNvwMFh/QP2MPlpv5i13trwrWsPfUqXyJW1vx99cfgR159
mmYUcSwlEost6hSTKfPpoyqb7QGb0cbI9XcA29fvJ5soqSdATIYBLfJm7/sybSvqPYlCOvPkoXs2
GKppbyDhP7pjHXY8Q9rzWIwU1diBg0F4eDSUAjWcRdit6aqu9YoZ0PddU50BqxgUJn7U445y1pQJ
H01fMdUtukFpN/lNXigvpq0CSszdsZUb6y0ULHm4wgoGD109seMxOLmbdHTNe6WVfBbHL3BlWt4I
FWTDDzWljveuhTX9/wtJzcCrsW34A87j9qcbCQSr/8e4zJ4uHDBqVPxCiAHUbwbKX6U2tTjJjNK5
9+1vbu498c6RZBdpZsW+DYaLGtZ3VBfh5r21awLpCAxKf0faRNaDG4ovhwt9Rp+HJfMKdHz72zG+
eyDz5+In1ywG0pPl7OKVOuX8PtsNuDPaPRkyIqO6h3u7btbeMIO6yccZng4oDrVznlUI71042z7P
mPxRcjRpC8LqQxrLlIrlMhRtO8Naj6182R6RWJ3KXShFaUATv0Pll45dkcWo6ABsrsep98jF06f6
Y5xt9JpwEjh1XC17JSMwfwIialhJ9HFqGpmmMeaKVw2R2J0at2nlRYtfXI9TCD9QOWjEtj+720mt
MRtLaUhK9tlVull8pLtwnquaH+T+cg4EY/NgvKe2Bs/zUgVbbpLc1uLeAeWgs34xMCvWeV1pMbKu
vfMpox7LueS+v56VeVK2HiKmbC9p9ol90EszACjev1wRutmtAPO3xol86hjuF9sEWSKQ9PT7HVn7
oKc3Fm2gcUABOjsH1jmNdE0EEA/6xwC8+Rq/lmVChSBX+7JcM603k6HqNQe8EKTFyOxlesZlFKxs
0/nIGciknv0P2zdmPslpeC7wUrx4OMdRJ9Df6VDvxUB/Xuf3A9uzwexAH5E5M4rvCKxOx69tLNuS
ygk7AI6xuEiFgPMlgglU80yi+OUvvKKNPPj0fGbE/4+Lwij/RBbcxZnqI7CZV4veBv5d6dg853Li
STTB2KqHXQbk6WtXEUN4IuQts6N+zMTaO3xqGU3Tyk/gbqQcZQ1orH8PcT5G6dsbAhTJ8JZQayGR
8Mqa0Dy3alf5Bxv00pqMlyyZ8IBQGCQ+0TGN+YK1VjzKUuxGlUCRJU/fXjAU+jMJR+cjW9RB58pM
3JNB1BdDyYvq0sYQth6QA+2kwmqg7O0MSWgiyVNzBVHf7INEwRsmCkfr4vrcVfWWGgBN5Ku43/Lq
cH5l1Z1rJ1910QmT9XizYJs9Og3WTYDNHvgKsVsWbx8ZknArGtQvv0BBtftVO/1NCYtRcKJgbMMA
jUsNbTJqChVdsTeWluBeBDL262cWbyX9YklKdjQgOFZXpqUsTjI9UUMv8QaMwCGp3FLcFhWNUiwk
MOOe66FAmxOw9odfSyVWPiwJ156vuFtO7jPm2ksWU3X7JqZAWKz1wB0hA2ncQolrVueFaKC2KzBn
IuwtEWApxpTLICtX7BItVJVSC9d79K/DbvLF1b8G0mIlshwWFAr7Dh+NBOsqPn5mLUIrRhGBe3Q2
3peLj/E2N8rJkNTQeZXMqpseItIfMqOrrxtdFYttAaoVG8qMOJX6tenN1afq/Gv2DEDZRv/AN3G4
XhobRBoCjgPO4UXmMErozH9SOuoTJZTxd8m958gGZqRqxv6n06DFlYkPSkXUdhnqt/2LypiJdKDt
ODVYiZHyljoZmqYOlU3+5G+7KWOzT8hFddB8qbWpnjLZ8bsP5lrphxjAcpoh+1xS3Ith2f2npDzX
rJJ2jAM0YICW2vHbj7y400ymXxhXVwPcHxpU8XaHKgaWcId6diaVSiiULlr3gVQCLjvvgu/eePcN
5Q6bqKkPf2vnsl8odxotBPdWn6RUUKLwglucyZ4+e46C74Ix6LHgV7k/hQFlnvPsTWjYV+YTbeCq
ZniaSvxnTLX3XGpruey1Fk8KPtDwvYwNnjlrcUn7dbHjNHYKpZOWg+ti+z/Bc0mS1+M8Iw4qgBVn
ouUdvOyp9Oni39yImWzveZwcf5Z8TyKq+c/6eB/cOvoMsRhnSmurqEPz898pAdpfcvO+nqSmuAmz
IS/pfq2it2f7J/4/ctoY6Y2YxgJPQF3H43TmJUDcY0dmy9ZHobwsCokzFIUpdE4U/4I8v83TNXAH
O1Y4aS0v5M80gdyW8RGSwZB0z+i5kDV7eWSTeRgC0MhLQW4J33bQXt6Y3EaseiEphwCUo3B9WDXT
pkT3dmD/e9Fislxa8v45JCJq6O9DcLsdwxcsBaz6Z1j38WmNkv+6iu2V1Zr2KURmIAb/c4ubBJ3o
tBvLHM8wHr0laerU3o5Gxir1Rwh8q1SWkQQVfXe5ExBuZ7NaJayxsJ9Holvq8wAkjs33b4ASG2g9
ypf3Wi5GEr1lru/8CyJWOxoU4AiYr7ozIHV+6bsiSzwP9XYficDE/5huSwKWU0dF8Hfws5AqYJ6i
nobeJwBgklXVWwfpIGwOhQoLFbI88DL+C/4dRsHNJKLAwe/iiHICCmw9ixBOCpZT2Bu+q45jyO+i
AU7/R1lIxsDBQiM6DPFlvoHXhJnpdXX2csfQL2liJ4KbFwR1WjaxGXG3KL/amrWem7VRkd7EUUwm
FeEvv3sNSm8NFaXT9edvAG9HeKfIC1rSb12l/d3g99dYQa6tdj/jN2ztScZqh9EvSTxTbC1OSmEE
7TqphhTG8T2YRLMjRSCDjNtoYYCojcrNdXXvammBLnZ4VDOjIo3VzLTaIFr1SYI4WBesuNGFwsMS
hD25fiIJaCcMZldI1tnkSwNyo4CyM0xavsG6cj9+VbeLtUr9Y+TEZ/IOXT760Vu6uGmPm3du/X3t
ShWU/hkNo9E0OA48th59v8LUSe2P4OcTdPDs/gYcL0wFnAC1btHYyfgnWhTC43UWeSlCLWIaynWj
sefY9Y6sOoB8RPjn+kjiXsvqtcu3fanxesEFOB9T5fpeUvbYcYT40ifrL4UvMBLYBfidyNBHyyjn
6tDFzcx0zAAD8IR7vKxHA9NfVG1CgK5pQp9QNk77TlJvPgKsYkf6Uv899PgSveiA90qeD/OeJaXD
SOVfdoExSZkUL+G8nKrAP4vZQS87qPZzA5ungvd52tbwjzPDAmbZoKDeKrLfWjKpE+fOJKx6YTks
wz8OYO8DfKLB7kq4s4UKwNKqvPFITtw4E1mOD2bRGdvv750A4+qbhScTJTxQfzo+Pr2X9iOXXwpR
WKWRJG1GN+5xxabTC+XVieeLJdRpyj9tEdFa1IqAtlV9Z0LvfVZcdjHDSnWmi5zgGPcYfgit9302
4hYQ2Kby10JWGMu7GKk9h7Nc3TkCJFqEYDQDXTBbkCompjvMppMoB6oKMBGJ9tOiR2NUsA+9sW/a
Qyu9W0gWStDTRu10VSu+tssauooQaFbpDc1DFGMVZSTp7PszHAN6H0H48rC3dV+BZQH8Uzfm/EqS
utopVXbMP/3KO3JXfIm+bE/qv/4qEha9JLG6YALzrFajGSrYN1keJKmJAdgnjFKvWaHaQaXxy81C
4XUqaCGzWNX1ezzlTtskFXUalnnpJpHsZGAYL02DNeT6AT5bB2WPfwJ39kNyOUaeDGfJW9Q1E7aV
VDUizRiJBrF7jyi6rmjillxBrb//r5eQAP6odyWUBpJsFNiIVA6Ntw/F0G2IrvwkHhsZneqK2pkt
ysPD2jsCsE01a/1NgO2z7oiNf7ps+b5547OO2IaaVd9M4c9oQ/adBxVeuiNcr+H44yPy/qNJzdgk
PMvo14VEFlNxdeUR0ztoyMV1vbZgn18AmVdR+Scv5dmKqVJwd4kDS5wC/ECBnHWZx1L6kSgmR5ZJ
oghXMc/QnWA6Z6Xfs7EgU4BYd4FpSaXY8qOMf46kT9462pXdlCGgywpfqaua70n1FQ9Lj+FcZzTA
FKkjB1sEWryqEwG+KLIq224FW/croYYI90Fmdo41UoCYKkR/e4pTf8ySUUhSZItVlkt0pzcaYvCV
Hw535E4uA7F3SxYFtHrKZDLmPN5P7p1//bSBHVndzYdcGh+moB7PYlBdad9aH9cEQPlFTRUBGVWx
4kKFN37l3sULRpATeCPgv4BSz2yHbLcZdW6NDC3U2wwl4rsME5cVoAxFcEd/haeBp4M1YpGvqsXf
sQpcuQHq/OXZzIpTHRA/uujPLXfH/N/OfGjKS3KSsao2TyRj77qh4wCdILVyS2M/yxBNG5Dq4eUa
YAKRnj16xVjxsj264D0qvZq+jU9W6GfN9sAHkeVmKFI0leR8UFNaUfurXsPqSxjf7cIibbTnUpsD
oP/Qv8ya4KEKufJiLshlxOGTwS8875DKlr6qMws1rX/3qOlyyEzlV9Akrpkod64mVcdVnycdpvrQ
HlSpF/pgwhCkU610Hx9p+shc7IF889F+5iF8gNz7TBr8jEEtGZE9zdXTnQS1HUkFJ/nRFHgBli/t
E+C4oG00f0z3ysCl5708c3KfN49s3sO1k1xXnVu9YcghP1pB8F/x12Lip1RY2N/hUty4MEFO8njX
DDC24ikf1og5BtVjKM7NSIfcU73oxx4e2gnAOpKAEpDEpnTGZQQR+dRXgiRK2vptmzKkQan0Xm27
+jkS0hlSZgk6bZdy9Tu2UeThzDjrEIp2hz1NikxM+4jJqD61cJz7CTU1EtJcpni/7koW6rH89NZc
ucANUPhKw5q/iBTSQT754p3LqCj2QlKu3Fs0/LJVeybN2VvLMHUPzsDTloXpadeFREC6CxwQAYWr
0Jf7IrY/qUTVfdlsFjUFvYxOOks6qBLOFd1/BAphqybi2CdCanPnykcoY/tDTr7STgEYxitwmQsB
HJtVTOK8GT9xkau545aCB8b7N8kQ+vFotcxLm0sLY8UdAbKam0DR7P4dfKRmYh8ZAsIMbOsN+AI6
GiCQf3nEY260HVV6lHp5WlS10uP5jRy2QFSwM1H1ASpb4J3GRs4TuYljpN81eta9gIJl9yTtQdtO
l1zUt0GDrD60VPEe2OJy2vwGln01EW/4xOamwEGoosUHjwCPyw6XNXV0tR/sxry13Cbg53Safqhc
tSIQ4TnRcDfUocnbQ2Eh3wLtz+4pqfWnuxlZj3YhH8BU7Hhy8F9SwkNbXFShTHAwMwER4R/61A5B
hTJjhKq41bxN1r0xeTx1J1bROj5am6+O1AGf9WQKR2CPfs+4Wu96SI+mvsD9r5buoXjrfFWKqCqB
oClvlyvw2YwOwDd5TPR3LL1I/cYuLtPJXNz9a9gQOgIZc+Egng8ITlygPk896+FXt1so6i55K9Wa
MNS2+d2qSz0i7CppLMcxclWUR6mQaJA7HNrOuFpsxqDkgwqgthXrsdXS/4caB9sXWDxb+vIbVaMn
aMHVPb81qszTqjvNI+c6WgP9u9DEvohcneTtCNR4MncVgWcq4g9BM8jIxNiu7srSudVdRKxE4lM5
m3BQxXAMoCJhbT0omYCUnWJ67rRzTh1pJ1CaXfq0mdbWGKFgm2l6LuKi9cr6k70yH7zgdswwe51H
kQzGsEBYcL3xSk8jD0iDpFHumCeHIOwRFkMX3aJPUaIDeB6DwPMJNBp1SKMNdw2UClaW5V6fmxjk
f2q5jld/GmgsAxSOxBkewtEQ5elcV/l/JwxJnWvjuDj5jDNIQ+pySIsRqr0OfLJL0aj3dQ1a+XXf
qad/UHdcev1LFMxy1WAZSs8hXUczXmwXRQ0bhAue3AFf/HBrTTxlwLa+lhLOrzNbcGrrbqvapADg
diWraeF+uGIJOPBV43ZsncRsPmT4fRoEtzmorl4+01/kldmxWdE+oWND4J7lgbLmVLHwbXH5cTCV
d9axbi8qftPQvs2fAqZxoBHxU/ZcXlc+L4LqWHnyU5UQhwc7VLAkneC3Jksd+zKhOCE4Uq4N6nuG
yP5WeRz4Uzx1YCIdoRWC/XY+J1lI7X5rLruIsy7lz7ikZg0US9yLKNYtJruwgkpckEsDUtXeKVtf
bnSfh+XzyOU84rsEC55HhfKK7yyksq3VxGYkMIz1O0nsuQUwdQGB1laALz6XjAEYV65LqODVD7OW
G+Zlbsa8AMJw5UxxEg+XZRAGo4hhgsRirHNL0D2RzCTHOzwqtJ+8OokIyNhmIs6iXul758YPjRxh
olzcP8NUHk1OYMyMAX5SSrqqU+VHDNCUzWYkcD+ZcsIW4CuxxqjI0woAzulkHYW2dmS7QdIflqK1
UB6xfZCnoTpNVNgfNWeAwT7pG/U1nNmTj8/tAucQt0PxXHOS+Qh01zcGyTOTxfmFJaHjXMPr3D0t
sKCuOiWO6laK3HfgNi7UuQXSFHI03zjLKjx8+iBqp8ZJGgLEO+vyMQovzgkzwLofNCwdSvDsIyCg
jrDLF3yu+5dzVAVFUQwBwtPE09cCQVbCff4RK+kMRpAUFg4atymsw2R0QtvljFWWkJ1kF2faSYxc
YUs8SLyhbed1aIlvhpzCx6ZizqSx1s/0S4r66yO13ZpCPO55WRxbgIXFkoxjtpkYfG8Vab6B3EEc
8Oq1Pnsz4aG5AdkxVhvujDCpVJfoBEf/fsqHUKoCNkSsTM8FnH6uogisUxENlPewENm2/yZc1RWY
eaIQyIPhdIwbnW9IM6iJxe9/Ucj9St5QO03BgPFgGRxTqHtvMxuKt/skEE269+IWvDb+R72WzWmx
hVdZ2HQD3c2I+v9yjECmpCLjMsvJDlUnH3xcr7RXO2dtDk8H1sAlA+nmlEMbmuOqZxatTkx6QzHF
h/pK1JP4K0lz4kmP+0sHZ2VuRsoKqW8N762jqkeemG2sucyfqW65W2Nds9fGLz8KNAig+1nW9Zi/
WS5RRxYxF5gW4c2b5Nkb4AvMOkBqvWWAzl674WhW7Zk/snF/5bDL+R0zk4zuDTxUsa8ZgZyX9bF2
NnyKsIBVZ1Oh0f1iIyKPwaaHlr1AXEOM/4RtTd2YLopLSuIK/efuYM+ysPukbHVUoxsOrr+d2nSQ
6tsptmyGHZPaZJsTeQZeaKJCuPLIp1oOCYHSKj9TUC8WJ/EM5j23RocDYEe6t2Ccg4MPWHZ8Ltyg
pVh+BPZRreJHLMg3DOB0PEwdXVY+y1QHl7vomklPkO0+hBwAbSJ+N18VmEtzThzjv9rBOHIOUUYr
MFK1o3t/iIQPtVvkFAl5lZq9t+Kqs9kbZ9/gxFwv9d2580/PH+YqIe4IsHCddmvT3dJ+oh35z/di
islRNL51jcuLkynm5BlLj1PXj0w0q3UT5jJbp59TMLZZI/lGrmSAujW5AlQX7KJDdCeoSuQeIydO
TalFgadTrpCT4TT9/s38WkVqOQ2JcxP7ufzP0HmSbE1cX/clmPZy9TsTQmU31rC4SkcDAJKLNhYt
USWIqgICiZIKx/UD0QHKadWwGYVfXX3xiUb1KHMiMv2Rt4UAbFuhi1vNygPLRxJ+YLSYGw2wEErc
u01yPxNu6CjWojrfYAEZwRPgS2eNH+cksNWxdU6DHqRo2lcvqXDEgek/P1Qbuh2MseXyQcMIMSdd
hk5CF993eQ6Y+1C8Y/b1Rwa86C2vTLyUg6mZFimBLQ2M8lQQ3i/er4l1/dzn1urIvH6G9MJdLx4G
PIte4U2HZkYwNKJeyUb/HsEQMDDN6TWu4xfjKFgvzB0Lc+1fo6sJMmVnJkikdsL+XPTsepgqBoGM
RvI0HRVLUTXhmhhYDSTbh2P1csJr+8hMBMkj4a6CHLZIPdz6Y3kRMnvlpaMvewgpdBfAgBOudBZt
e7Ve1rFO99V+SqRc4qNPV0xQy7zjdLqekxgBBgy6EaUXIbukTnT35dm5qQ5T3Kb9ojkh4bOaJ0va
wTSqt+zvAv5bdiZm3fhI59v4e4j+/aoLEEua/HG4rsQiHUlyJw6zUEcV+ZPl/33IBl7fst+wEv//
5eVjVcMnzq56iqTNhgNQkzokIOZKq1mUqV7MoN4UWq5hqWl2js6Q9Ac+ZAlZ2IqIsre2LD1CkvXr
N21QkVCXA+x3D/6OOO+tvXPXLSczh8wVzdvQouA0jmkVSeJjxZWJhTKbPEl+Y7AnoYee4WVl4wTV
5SuHGTRcm5+WwBXeSgDJ+7YYLf/5kAjTuFaC209iw/qvIbFoUtuw2lLbC8yHPi0xwGgP7/9bBouN
kMLhKtv20KexYuZidG8AF5S8XmHxaXneQ4UX85GCrbVRlpomTEoP7Yqw4y5GgXNKPptAeNl9sUCz
hAGav1KxP0Pul34U0lHJz0McOwudb0lleSsSzOhmO9KsujVfqQUWHHZaJSyloO/chPFxvVQB28hV
akVe+S1pTNpD3oVoJfMpQchhdnfRw+qQlLIXrVS7uwI5LcuX76UIGCApeqoquoZbmtPO2mYVqPkQ
osONGwID9uRSLoppq7+6DS9rntlw2vkRgvy9e6f9fN1RFDiwkvulyzgelhXXxeP8RVLpKe/d61jE
J6mZCSjNwvt0wAubE/QKU145sy6043XSdw6Dg27K+eWHYKYIRIukNFIhn+Lw/3R7igGYmpAmrC9n
3dMIjFGd0iONOwNfLMeqJAghCHPiKwA9DdRlu7M7woQhtk4GngWcEK9Y6HVDdf4/g20WSRRkXpE1
JNOJRgf8A57w9DPnWfe/0ZliPUBL/mHf26YjAkxWjNCvBRJiwlgRxARoNvL7jzZlQ/piaoAka4pk
N/U2gLxfmpJwVXZv4pJO8bBCT5XcSD9AbMvHp5ep/KlDUNNm+2/EfrpN3j8vaIcyERCAc9Pfhm14
7uzmP1vpFsgMkkCiUhd70otcBTRB4joKvxUSxbD9JrU0dOiEI0wym72wZVF2LDjp5/6lFqw2CBlO
E/a/dNCZxCnNRCPUO+tegltetxhyo7EYjLjnGYGTJFgEWgt6JyWmtPttyfkNPQOr3KXdP2smhafA
3SB32oBrv5Cyk3ePTlVDl6rwnc/Ahl66T3/fFJhzGwEKYgIhppF2CcB5fT/pzvBAZSQY43lcxk2z
yyxjQ2RXqI1y5S3gdcZXQ1vzaGwsqp+v5mmGd4Z2xv6T5PJNU1Ajx+IduB9v6hB0IRzdfbqi4kaa
vptW2Oz65vhRaIBdpf6H1T1prO/DT/ryg/pCrzNyRbAnmBrwKBt3pEKbJQH1MLVZ/JuzD57xXqSe
nLiReu0oNFsWMQY+h1MZ0EVuX2+Nfq1cAa//Inbwbx+RA6IGdO3KmC0/vbDLnYNRqPKvJE9VAvDl
N3YsRNo3NV12j7wO0drUqxTmg69AZ3Yhhb1zL742O5wzSBX9peOMKihMlBhW69iQngdRx9/BpE1Q
lxKYfGEEbj6HnQl47QXv3n5AeTAKMet2h+Sy7m4vf/bRfyRa1THF84rcS1AuTLdzYWn7dJ9R7McW
45TVJN6/ERX1K/yxb9994f1iLKHzJjOcDFqIZvMqJk7y6Uy/JV6AGxDkyjVqtS328OpAWAC5JPLP
oIKJciIUqjq2KmV0CkM/vJqwEeapTRyprSOoaKLhw+Ppyylw3uFCNssaUsQxSGgQOoRSE9+nDK/m
Kp2zFiS1j7HX0wwr5II00FjjGPuvyMjYhZhPO3FQiqhwyvDB3Zh6H+S77dVpOGgnrs+RQKKTPVIQ
wYUvLXgmg6zmS58N/WzgmbHkq4C7Ct3ydP5fcpPHi42XS3B1/JewvYLeyscLQTP66dS1/BdRiphC
KjGw0Md8lnvEPMKacV2mpnPfitVb7/Jl7TxjZkG8JT+F6vlznUdkCHCZRgE6kRElCJF/THcDuvzH
+wzAj9FWr1AeA3y5OJf+rlslU11Ghg4EiE0wuCGaO0IQTeJ6si1L0dzTKSAM4Xy5xaCuAyVcXcAz
xpMd6NKDhm2ztXjc3iE0EmNjeBDzGqrjZfNJmssvZ/IT5Qh7cqA5VhKWz8FwY/7pht1V9eaD04dV
w/jyi2NvROKljp5WszSh9etcghI5j2gkVa74i4q6fQjJBDqN18CRItsVNtb5jkORfm0Umr+22qYY
8taG0Pxy8IneIcqJfrdG6QAjMqUAeKH9QFP+TkcJL8wPqJ5OS2hcXHbspDAfUHDaxvM1UmeWE3gb
u52wlRmt1rBu+c9BBufSQERiBwCmXte2CuL+tiQIhU5ljxca00JNOcFJo1kpLVdH8MLjug7xDZA7
wYs+4OLyGYgaoizpVEHOaJxGRrkfbhFNT+XDmQmOIJoBVoQYKIIn/fNQA06vA71AWGNr57ERBCNN
7VvZ5zIFyrHuXpGxTpeYm1MLeEVahtKWBhXg+7mg3m0ZATm3Mg0jGw5AL3982dCv+G5pa5pbupKb
myN+Jw25nDhrULcSjkQuA+hqwrMy3/o0I0mMPKQYtMsfhF0AAp1jVnsZSCTTulja73eB2Nocf19c
DAz5Tj+rj2CfH6v0T44cd/Zi7X45xPMFXu60Ajsl3+geOrTZytHNYqO1VUGO/mzifA8sTm9ttp5u
WkiQC6JhEoUfsJi4GDE69EHWYwFPoQ63Jsk5/h4OBSLIFEmhr1FVJ75xQF5wgHYQIdB5pScgc7A0
ZVkPTIJ4dLiPu08QBlWY4xXZfXH4NM4FpelG6RahB0f3U0/rRoE6rcQit9CPy5JliqVGF4WEuExE
d4A5jK3YZaP/xAfEr3fJkQWoYgBd/3mHPpf3rkW2XhdO4HUuYYd+SibcNvTTIxfrKO2TKP4lQDaB
n6DfGU6D9invj2BxYLYEaTWrAkL43zUzIbIKITom/IKTuy5+h2fHwFnLaUAUZ5kqlLk6eWtaMmkE
DeTjm5E7kP/WaO9I7ZCZRhQhomzSlNYK8RMbtLynu0i/lOcInoRVnLFt4dvqviMY2FN+OktOu8Py
1n+3T2rGCkh/3oj5PLtV0AlAiziOZ+U3KnVsbwUZ5O6zYIFtHzONQVc0blQuGsUkzFGP9oTl8OAN
14NAXJQmQXtwUGBLmCLOOA55x3ufAgVnhj7ZaIYpXjSv8E/8Z/7c8RBu8/Xk7HfuRxBWBECyOVYH
Z1sqE/u/uUKMH3J2favCoczDlOKEcveQqaXedFh+YAP+dYXIKx3oGUdoWDTHcXwEoBLZiIsZ03cJ
OusILHOUmSv0bS+rBg/llQn/2HwLbAJsqvLIVzTrZWRdrJKIXpUuXJXDV26mb023ORAXN3dIc6Zh
ldhtmgl7qwnDRgrwBI1yUggv6vHWA6K13lEhmXTHG678iv2lL6noRZ1Ct/VqDeltURSvRx3kmMf/
MbEFhzTCwWYwu066VjL/dXaV7Qiy05RVEAz1ufG2v7rA7Zno32cKhyc1xb6smH/AWLm/vFUobQjL
ziWfBUBhiCinWA68yowHzJEsL2N0nW7uj0hdF2YKDajPugYaBbFIo2aTS4sXXEVPiea+5ecKDYnP
PtVp7eohwz2rMc6ZWT+mQCik1/8ZEiTNC0P60netwNZE5oMuS4F9tgF2jLOWBHHC2tGWws0RuNuX
iKtnxwVzOSb4hhL/zXWDbnekLOMSHORNM25IgVlxCXk+n2h5KxrUaiMXVSKLf8j91nXtpQvZFOju
V7VJOxhi40Z0GJ+dmAkM/p/yo77I8B6hVtg6krMHFz3rCe5AZ57FGKD5HJdzF6lcX2fnNBupkMh1
sdBh96+N+DsvgNF31MGC/AOOxNke2sK2vRz7EPsZP8+uEdBdoYCzR6HaWpUuXkFOrN+BjG1E7hDX
J97FpoRRd7qqb0gPwOq0hU1mXgZpYSrNV1No681w8LOQ2FKDGRvKvfDEZ5m0X3c7AkmthkgXJ6UQ
+WH7fp6bYqp/nR0lfJWDGsy9BKH11YpzWXZ1txDmGdanD2BxHW4hl0FvHVEUK/yHJD9w0PrvJKzq
YX4UDHNGTLTmvNQ9BkF3g+VKlW3JDNnVrVaoAneMyg4NLqnJMd6Mp8CUvMWQWpqPsa2pzmU+hdgt
xd+VsQp3U7mqPtkp4KH9g3jb62/ByxGsbT4sRun4v4D8WeghfPjpJ4JKECMT6WkQIF9X5qxrw3mo
UI+voxz2heeqV9/1dccgXpKDnJht0OX3ubzQWpQ3FqyzeuUs3/cPQBS6SBiV8C7QQr8HyRFfoYJz
kfvGXrXrtjjV/aDcKM6o909KNyMhV2nXG2/YN1AWFH3b+Won6WnbArtmnvM1X8+t4w4A8Qd/7mDc
+5f9X6PrYEHv+UXUEa7qCHUhkdFYkyrnrSty2Camq3Nyxy6nbebrBDpjbF6USGs7s8XwkN1NVT57
pj6nxWVxj6XfqIIHohr0CfJip+9K6h/+M5W1jxWqnP0yBx4FDtBmNaIJeTdZsWcrguAYAYqTwfPM
+8wDP6c+i8U5NmkkHUDGFw4nWnzZagq654XG4iqyyS39YeTZVDxulUQZ7jv5Uf4e463JBmGkI3c4
EQRCKgcE3H4Lhn70Dt5ulN8etfKROh37qrFR7apg0hKognOEw/88q55blPfTalZB6d+YjcCcHN9O
P63f5Y3dxsmb/7AGPNr3k5WfHZkC6fSl3Wq6nwpzR9RXLqOiSNjJ3qgoYJywhJxB/Wb2+3djRQjL
f6PUFCdXTjMhZbRQS9Ou8O+8lwO0pR6uAdJVXoytwNstrbj2mel01jgBr1i9LDkddL/TXMjs/nx1
02RSb/9j/xnH6XXO2p6Ai4JvYncyA5R8qJ5Zy7U0/4qSRWrdYFIb9gySrgWcHhqWPdipfgmcpVNP
9QT1sbX2FLU8jNNgJ38JxffU6xtv8YXHhJf2USd/7M9rNPNDMmicBXD6B2V9s5l9TSrZyG61OnnB
iHr3YLKMg106EFyo4fy4O+1xiSDwrZk2RU/uDRTrHcVrrnuXRbQlgnCg0TkzVh1k7HRumgNfFkdk
kdQ9ZmADiTzXiP5WW7llVrtTduev5vadb0hBjo4Xqv5l6yw+nOxQEv70kYaP7xzz8364ug8goPzC
57ELAewKx9KbyWt+NcJ3dSrLFKsVqLPtBjtV/SA+KPGiXZZQOHcDmqTS5yF/a0PX6U3Z6jqjKKPS
yHyRpqCoHAkftMEkLvUc9V3I210uH5bH/mdkTpKfWgeU3Z8tbhiT0kInvT+FlElZFVgFkveoZc/2
33C/KjJGT1PvEP4J/8Y/AeBIx3B6noZdLYBIBtWds/UwXzQArweWIbVE0fngdIyakE0mfr4FTO+4
roh9PQwDxOKGUSV54VTuS0ZXq8GO0hNOAsmT9eY0OGzRIuoHDZcnl73oOka14qHgDcwSo4xsmdWH
WBG0j9LN9CvgevNLO9x0OoY/e3JF79zNpIZJ8OhtKge4EGmliOGfX3Lyy3lc2hu/NChGJHBEhVaQ
jhFQH4+iLZhVG/BH2Q2Obl32VYRwbqaOlTKqe60sP98jiS9GgWvzLrMTEvFM0SqgH/xU5YB9jV6a
DSCYPHknIlXJdo0Ai4YEPmb9iEHg4eKWvkW8KBmKI3Qz3i/SYpc4NPq5DwxfldohfmzNmM8u+tAv
RuOx+hqD8XzCA/c+sBrArkHeExK6cN6ByS3fJGHZYrJnehlZxUgDmzV9Gbh+7X3QxbxXkh6G6t5F
honppdf63meiWqA2FlQEaXeUSLnjbNJ+TzwMU5LoiDvznuoSUYtMVtkswURTz+p7MxCW1D4EAAJv
gx3KJLaPV89ZDWmgJRgbKy3CG16ciU0FtdvimmW6l8Fc11bywAsKfIKzXUe+HJqKfW3MajeWbgad
auDTC9XZ/GFzHnt89BIiS7VV7tNXNFXaVmMb0Sg7KCJerzNrj7tCzTK6ZQujWX8TPuGkcGfncHeR
bKxPJlIhqohXntxCB0KtXYnjGXyd6mfGqXVTXE65jVetNyMY8ya5ruNkDsx+c1cqNuGOS/xNChgI
n1SUe6W/fTTLFBcmVpnBt9O464O81jYELTpVAntbGgm5qTHsg9FpsegKdZpK3d9tY5o+KhKl0pQ9
IjeV4Xf/5uDcvgu/KWlzrPNgLI9TnrxNatFWAD4DCgGBrxv3vylJchbpb3c/42tHAmeSnO0QJp4Y
RB8WvUQC4f+3g7iquKlEQmI77vj3SY91YNge14sohN7SrGtj7kUdSelibceuU/1Oqqge/2gns7yb
tsudxUH2D7oEqv7ZC2rM4xwA3HFDBL140WnGjUD1H6saidEQb5T7X0awcnFvv6BI1DcTkz9eb3Gj
azjVeYiizb7ie2cGN6ezYuV1W2hQaHsARk1dhlOEy38YmHg4b/sCcflE2c1yqhjRO6WV61wuQ0kM
qSeVuxr8F7Gs7Osrtegd6bpzNMEtKbQ0tjqNdQuNrEt1sg8faxMp0tZ5JiTTj42WiPZ8V+xAUQoU
apHJorHOAUJTVFiXnqwIz/iUZtI9tirqCNZAa5TUy4KmIyC5kJWOgXVC0BnikN+dg9cyKPlayz7X
BR0IogZOGP6W2VP2H+ylJ15HCoWW+U7LOJYC0DHo9IpSCRze5+VuqRj8J+RvhyJ6W6atvX+4BNrL
IrD8kovP1vsErlr5RoC3ys8UbdHKIM6f/2J8q+PUGWdf0Hdv+fTd5SjU1Zap+XCDtI8DXMOcZ3qx
qydUoCTJKSZxF/j5/mWbTHSjW12hdZl9sx1pZbfSGCkDBAP50AL0hWBvPOyeak0fkpKKxJQ8o5Oi
7isfvzo0oOB+DdTzNfExBPJOFljsrBJvs4JF2hsVHT51stD8SQfrBad5CeUTkS/a3bI88exOOJ97
Ua85D42ZAadd9yxZigRF7ywmBgG8lXzuPAcRF6DKHNTt1yrw6KFPbEm1JAVDMOFQ0tI/ioWNqhjO
njhuKEcqJDyQraJhhQuGP6H/EFvyEL4ORhxtXaXyH1ja3SlnOyEk3tH948tzM+sxHFDMoRPWgZbD
lf7axI6MMMiCbIFUDn+5lpBbCu9mkkYGUmgb5AchxsvmuKMfUOYPV+wxxMpUsa27ob5C5VYcGxQg
XVp7mwdkGNqk/IO9+LwtuIXonf7BXfH71T+VdGBm8tGW101tzKCoiGN7yUh4ThjMrcY9vak2pZ+t
K/2NROjCFnV7niWqp5YaDetljB/OTILeCRZuHn1mMX1f0ixFPIAKMil95zMwvcRvrGCxNbob/Q+Y
5/jZaiRAvp3271tPf5xkMwdy0vQU3iqJcAv4BEzD8mo68fgb0kCnzaQ/LJ7QqNnA5Cj/67tBlgx0
DwzOF6rLOEHh2cBb69JbCZtXdjrRJfyWVhbX0K/4oDKydpDClzWPc3lmMXAC5Lb+lB8AoqCgF4Ci
ydxFXq+qi++3yyWT68XeDVUttfxnFAf62HZPl13Hyr6G2icJzS2A3IVAU+D9pEQv3tsU3krEJ1zU
426grVyXmwGqYTLSOrp0lsahRydxxLl/5sBCmigB01slEaovBrhgNZN/ObCJIZ9/DKapusllbEdD
RtML6EytiTII8lDLZ+qD42un7bMM4oGOtexsIFdqHOZgE7HtLei1ImNbBb4pYpo4K+hOVPCzWL0+
GBPJysX+hbvYne/RbmsLx/3yJeqRkQ4m4Mf6CNm3TnHIXGaHLHHFF/qxisiAPhbB6YkDoMrw9ztO
vh5jGjCGAERmR62se6QVqPCfBwjMddEElqXqAAYrrfF47L3zdlink1Er0e52YpTP7Ax8kN6MY+HM
VM20AfcOq3g7zd+1GPYsoxq9j2BoEn6Gp/KjLwwXdCkLnE//iTQ/UCcbwgklcyyCiaDA1wbS2TK5
IoPI9pC2Q12+ShakOrlZVfWaTzfNskWwF83k+/YfejPhATFuPH15H9WcnoZa7ZpCJriiZgMTTa5h
xmxzaetEhDJ1q8x1kD/upPVunRWO1ArQM6AAlIQkOVM821I27cfT3HU3jItLg7T2Rr9iHm7GoHn7
Q4BdtxVJGc5cVWIuwPwS6RPYg4HXmKb9CCMet49IJO4sX5PXyIaHIrwzpewL/x58BcrK9sEOrtLl
FkJX3EHsoBifsMnGOF+t0tMfqXRlljUzh3X2DruAHXaLxNiU+VHzYM6xWVgYHAu+2CAkK78PO1Ce
whSAdqR04yfnxGU38H16clLLstwYt0wNtLxVAB+l8zNCARSqHZAR2i/hJj4D91EJ0ZmGI3iE9IOa
zTJ6Z75zXdhrqgHtBquUCuJmWpG5gVoe9g1Otz2lFbVnnR4Or7l+JKR2FGbDf1e2RKHNcCsramkN
YERVq2NHOi6dcmXC8KnQmLJcQ/zrIC0MmU9nD6//BnTpQUTgcwi+v8DKKCkBnEr0UiJZ1d9gmG70
fYrj+OqnpF4TT+5MTCLkuaDr05snVdmB/Us6nZPhPZCkHkcZWrCN6SKFCR2xiq8J+xGx9NCHNF+W
d3rMpa/VbGqUuhylZV7hqwkfYlvYbpD5EIpBJpl3U/SCPg1FZgBoZjnH9TiCn9y3RD45RUgUbQ02
6t/Sj+1Hv8ry72BwZ5dpCURypu6QUw3pw7RDY/T2ljLzTeFkarHNBy3Wvi+XU9hNjQnxHHBUEUVn
Y+SY+ktlNl0upVYH/laf+41AxwBTtSWAqeIEi67PPNBu2u668xf6pYy0j6dHmnXqSh+IlYgQUpnf
lneuAebkMB1ypfXS8cQ5R3c+P9MuTgxU6BiwwdJYx+w+JjIiHS+9zpHPlAyYlsNKyCNTUEDyAoBc
j/5OvCEJYF0VU5L30PeNN+lgkKgoA+AkyO2PlGb7YJj3B06gmrFgNfZnaj2X6eN4kaIX10M0cIZQ
s4kbH1U0dFpnjrFZA50v62cF8Y+TEe9vS8JqUITDbHVc9pNjtNpikaBCABsqBhgZzeGmC1wshWMy
vo220U50vAEuoaGUdsM7QQboNy03VsgoFNOYWfVeYUu6MyYOdFiCcN8SzAAxtSnD7ugyI7rsch6t
v2l459jvzKXqhCYazz50hM4NllE3MhNaDGK5C9lJNO6qWJs0ggXcivAhkY0KS4Rz4H2BFBnnauLy
0PRvGkIVE1nPJ19A/NM/eFTWLjcoTNOCjg+w1lQhpUFynRb8KE8RpRzJS2cinnvhQSaf7X1DUtKJ
KByytTT/M8T01WcDj63iv+oM0KFxLt4n+pRzkl72nktJDAtq0P3B1M0taB4m3g4JGg44bOtv8LU6
iIQkRKPAoUAsXYe7oAWVvaKIzpXX/TcUNlvV+D/AoxEXGBiWP7d3iZGM6RJrcGGMdNsUrPvVjJyG
Wn1Rphj7Fx/LcGX+XRawywb2BKBWKXhndkqgneF9f+xF3cLi3yX9A9ACOmltl0QxHqma7AbFpTTD
1OtIA1JAZZBxV1JOnC1lPBrxIH59WAdqbrJpMN9Qzj5Gf7YJdZsEptq7IOmK3MeuLgbGBBdg9/MO
NrcxsdeSN8c9p1WlZwvJigGhVS5tcfXMioHVj5Ju03t/otPlGUU1u1PSvI/HxxoHPn/QzPu9rB+P
RMF0ZDVKaHnwK6aBhYk2hUjFXDtzg/CGEiF//G7gN2AnP70QnmIT0QSa8DDRk6sSDAKbr/n6IJkS
N8RV1mqqB+jspI4Cl9TfbXXQMgBpLwkxdn1FrOn0StlRWCCdzo4NUOECnbyKSGaqUr5kMhU3/BYP
uU5GZJGSXlUic+CnVTGcaCA98BCbG0SD/3jpZr/2xn2fUg10kUeSUHvb/3vxm/TXqjKv9+ZoEsge
vng2I8ftBq4ZbuS8x7BOlrNeLW9rthdaoFYGDnWym+fbL2gkemKcEa5jIobRmETZ5qe1xZh651QO
OBkXJPC5BO1jYCG+dofQJ71b7fDDkCwy45frwvNxmoXY6HYaG9p+pk5ygYD1omJPquCZwBm94pF3
PYUGaHdSRF8S25rmq6NiPO/Glk3UBjnXXEZin27WLxfBCsbHeSPsp5sEnUdrUXetIrFrAe5OgJs3
zUpwXWk2AG5IKfWuSK5ABCvC1/BuAhspj0AwzDNgm1LhbTP727ZLSup4SZbzZpVcy1EryiLKR8mr
d5/bgakTPqIVLYccY5ViAN7J9c6UGPrlvNSlWD+NbhOPXqaZy/SiLuvAbJ0gxAEYq7s6e17mEA/N
cm9vvjvzm3k7RXq1m/eGvTqkunxPVLCfiPMfzun6wrSjyNdEh4jtKEpY3Wzo6kpRDrcfjcFoEAD3
xIKU7AnVNjetbMVSfK43Xsq/DElc7KNKBCBfBfY4+8iE9m7U5dgEllcN96rDtaEIfl8SaJ5srj8S
aAWPJ7JZvKoJZutfK9FXj0tG2rXU7mzS6Qq/MRSHExisgprsXLfdz8768uOblHZ/fbH2V+6AXuvK
e4IhToQsOEht+eMvEKDb9yiynmFCgwf1yEpwwHMUY/4dQx14XgcveWAK9YyyUVpHso370zqcMqZF
t8o/x+hY5nYQNfLGQD9/EvzVgxWy2XU8oupvKZCypU547aCfGSI/vvsNOSDM6zs/E9z5khwUltJf
sbl/P5ddWr2NcAQfb3obWoiKQ71GYC0YgbCswYiHBfrkLsxcsb/SSF01XlpUwjpKgYxotS3vPZnW
taW6Pj8yRJpFZyGcScLv+iGbeddM0HqqX7pS+WqLeLEBYsn6wWoQA2qxN4i9XZS5vwSHg/8VjRFw
RfF51lCMKhk+5mSB90X9FF8j4R5BfsP8BHE/y1CEWRwi74IAIkoY25jn8ODrGsm/kX9qj3o0WZ6t
V8XfUyg1IsLfO+nNSLPzhly83Q5KHdTrBmEiaTPBYf9lX6NCZ+EXu0prNwzwPbfB4hwuxyOQM1S6
L5FVS/x0/7hpK+sjlUAQvGS+JMhRRCI+l0mJfeGI8/AB9zsWg+MjqtaI9cvp4jIomOioQXEC3aAb
Ix8XOYbKQlLoP7XW0D52mvpBsVkvVEQiyvGbI231yr72JNek9oEauAtTYnKoI/f2jWoYTJTq9b41
J8vRvep5pZCAN7W9MV0aDMoxQbSP/GXzoo3Ki8/zQ1CTYt8LLgji59PYMdCZdrP6gqC5Sz5W/sks
yHfIJxAxrOYN1Ucjqnbr5a0jvWFjJwMLA+h5A+CrBOJDv9TdlzOINupF/yCpuRGegwiQoSi7Maob
sUL+CvBgzODbYOcfJooGF9OvzG2X+IDFlP4cfRGE58ns2sYyBey0NCwXY5RBdgT4kC6vVkpyeqos
gvhPgt3CEK1UyGStpU9FfgAet+3DJv00g+R+qcnC9kDNIZ5M/3zJ+uIdl1hhRrqQpr3P8sJSPNoF
Su080u3sHICBWvd7HXztPt6RPOn9jAnJhbA/jmkhcdw+Aby5xNP4iSslYitnDqF/lt4l/TVp23av
3I7y+L8BWVSBMytEHrOX/NtxQ5PnFeSyI+7JgWY0xtFSHy+5VZBOlpVLVL9KtMMDHlm/Q6Ud+4kQ
jvD7jlZ6M32vnQquix4/MpTAjSI7nJWbvr9L/oHaBUGxwsR1c6UbSTHJ6AedmLUSJlCXP4fnU/RN
A2foqygbUTViNwVeVT+XHHDSF1F5ofuPl60RyMgYt4gWbD1IlWDovHDe77T9BPxNvqVM6N4Tt4uq
uyZmKX4mPIqmxge4xK5MgVaxZaFK67FIRx2JjbUMMIofxqclX/IeIk+TZDvkiJc/4L9P4w8n6ysK
WL6Nn7oDGxNy22qq28i+uSLN3EOJWTVaB5/ava6qjCmVX5bL1OKzBibduyEaix7YdMocl+8NNccU
Ca/dkvCB3uvC0rVTBV2ZrC0suQyCH/XWTr5OWQi6JZO8KDkmyLYZxyrEC+8P/XxDI8EtOxQ40Vf9
AVQczAsoDEm39WnkaPJbvhkaMYS9bmeNYEQWiw7xAzHcjOKeHoevsWglwnLihvZfCLuqFDcU7AW2
v9ekBfBjub0xIMqrY9v7bCFZF588ErhiyejOwK6doiFhJ8NOev2b33I7eGpXcDGdmzfCMCoXtqyA
chvJXGoIyb5FjwyDwsg0TzjHBefZNoRfMtC3MOjgW9BLQApfK+ArIsm92XkAmSbQZz3b7q/DXG+Q
lnN3FjwNBWQykiVl3TV6Rkhoi54yoIOKLgGDXyItNKJ7KlQOe3b6syByz9OjjriyCSQ/t+Hyym+I
B5ehSNWGuwq0oo3n0tEgek+7UzQ65/kTg8IyZiASKwBeVg5/OC8z4DWaewHgQrxYOa82je5mpCP1
ehNXIGm9M/svE7RH32CZw6xBd/hP+apAYgaqOFVPHQR4w9EGNXdnooxIjt2mqNvahI9JyJAsfZsy
1FSsOy418tbRkYH1r3JRlAyzj5VC/BIMl/jPZeyeX0yvNrM+lmxwFN8IQrYr+rvpEeu4P+/Hdo1y
LiJcKn+2LKPWEcd2vQ7AVCJWfTyraM12y7VGbJfjKCQnnf90i8JFtgamoreivphG/3KghGjt5Pa/
xhpcm+kk56TREI6FsTAWg2KiyBu+CTTYJwuiOZC7ickShUeWie3FxotfePo3VRZWjquhVxDTVbJB
NhCBtwDkW2sW1DhQ5VjFJA6PrklMaspqcuNfNynMq0RUWTif6wYo9oyW3wajQjTUZIa6Adhs+++d
u3gMePJAdUZORRczfeXrUqf/HYhSKw9kQd449tAR1iGDefDM95KLRhrBDX54vODwK1Df6QkfsHRS
Pzq2tQIGl6JTWOATJPhoRtrYuhruquFn7isppCLkdmtiyC+jx+ds1grpm3C2CXZUMzB9mv3536P0
ClDFj3+PIHiW2H4EYOEAqo5I17/EP8xy6g5xhUgLoZ9ewo/h3LdrLrGEuPRYtCR3GTXT6+ksdcaV
KevOa8+A1DKo2xb0jVOcibexUUjvOqMZqvd1az4JT7z6XLmTwMhx6zIBoUYdflZBgtLzI2Hnd3HY
85uMBoCZS//Nt3FaZ2PdUqxp5rTgb1U0bjhD60ufgyRspx8YuqwZS201s/aTicczyRkCF75S3Coe
DgD9eOFS6JLTIfpYjDmd9hqR+WOBV7+TOiDaeui63HcR8FCZ1VNcAjcjKHuyUu2nEh6RbRHegc+F
En0oURzSz4qxcnM+WB9Zlg6WCPkkcuc7TnY6GVSnh6ncomMF/sAq0P3ZWkixd8O6W46mIicHwz/T
QaKAZnjZQ5C0G5V+xVI1nJRyXmUUrt6TRTb73qX7G+1QnkegcQq2LTz/ooGaCWnITetjX1b824RR
nUs7zxxgDjQx/cfcExCIksUzd/VboBnR/STqAeNm/z/qPEAqyKXfT15MolvIsEF0dYyRTKtXLW/9
ao0hYu9KZXW6IlJN2+dra7XOzPQ40ARsksXItubQktvYZlZympt0a6OdEEfeDRVZx3mS6lBuZP0b
YlqKT5fWdf2DHJKGQIhZc1WLagkNTz7VArXiJtvWi4fYJ1UZWBG8L8qPIYHrU+LCz+/94whgAYIY
4HfB0MAaQ18+RSMJ1B/sPclNRZsgjY+qF9MVXzfzpf+1hqlNLapmiDD7l50lrurcwgivPRUDTGRI
aem0c8OG1A1QciJnLoLiAGDvoAInYkwiWonT7r52UTkmENOkxiCANLVb4BROjDYpzfezfXORdIUH
/Z84WVxRSMJ8PpcXNk7j7CgqOR0SvX+64D/xGlo1AUG/THhPH/bZWm22aPBpUNQMvRnU4oUzywoh
OLPsQNCS8H4rWZZJecCEVFJRveX52TTwHIrjJoLy2d+erCDOpywhpZEnl+FwXEn4z42+7AYylcbY
R5j+6SRapOKIruKDcaLSczPAtqEKynpP5THSDqaf6HbqCpBjI4owngyHhR5d1sbuyyNlizJJ2nQX
pFS8K82pkrJsZ/gc2NtHAGWSr4Vb2IEXWJFIOppJbSVFkuQafhbr5oMnKtsRcpEDbAKJrgflDgNv
0uVTUuNdjM6chDDFb4bLCJt2C2kt0lQQIS4ZmFJfCiEMD/RfTuU/6BCiyFkX73LXMHb5OlIRHYeF
mbHVkHr2l8R3g1pH4w3VrSCPypwLtQ9SKVFTC/BMJRAWt1QCCMLsscuO0VSge9madgXrik4EEXx9
UEbuubWHjdfhumBBsa5Fm7o/GnmZs3xErQ1bGOax/eMXqRr/J3I70CIMOY4ATLrEbE2RVKWy898O
5uJmw3zQTcN/05+kwfn0h3DP1tMJm/R2mBEfwEpB21mMJch947C8LNaPkylRlxndtz8FQACXvjvi
fnBSc5PHOpzKaSU4TeSuYKx0akCV5V6axqOsIOEpUUY+CC8BPoAI9VdnMQ0aqrk7xi1X6wYEVVHc
1QSmRIDpjJYKcepfCY05bllxD84Nnic+bK8zYfJkUzWH5R4xssrKsIsOJ6BTrpC4sI0f66byMqEb
fyExQP1uIhu/yLf7tKz24uqNnbT3VYrE81baCjsA8Dz2NvAkF6lZogutLWJhNZ5dwB0UuRCqqEPu
rOwqeOBeP561g6RK0UE43lRTKPdYk1WBITuMhyWR4240M/joyU8dOv+//W2K/CkShBQgebMtZWPy
1EsunXdFgCKSai4HhgPTjoOBpZEn2mqSCHjhrR4vjKVCAoj3LYnj2cVdnq6+ptvzKrM3H0zyrHhz
WmrxpyOafocH/nQMqOHjrFD4uZ4d3JH88t0AbvzPnY8xsYpdl78CcXpUYbjebqDE/jdebc7W7NgL
UkC+kAvlHqokcScj5ErQymtqGYv/8MMdFPpl168t2BIiaijX5wBY4wrhRhT3iBOBA09oVfuy1fTv
9vz5kxtVv9EXgQYGjZ3Tn0ArWsvgV5139ucxhErFk7VEFWPB6p7r9UNgljWZzOcxmOrQ16lvxDaV
+npM92JdrP5/6JrYUJuzbMxy1NR7dtUArih96p34IC7xHxHymR4dPrkrOWYTb2O8x+QdgvxelDgS
ok0oGE8S4h2zRmi8d4s3x+QcePBA3l8LBh3MHreVC+bEn1U/ZZ0rfksh+Zj6ysleCp2grlN+Q8Ok
XaP1IaVm0566cQB4yDe6qE99YKrpc5UZDNYexDNnn+I6vzux4nf61HDNzvbuJ9HCORLk3Ik17J6D
p2hZhfVxkRgZZn/EPvZzKz1cffiqYH55h6GG33UmB2ulUmTbPgHyOZVHzZdNZm7/1PcLL8e3jOr9
OaNddloZGq34PO5ooQcCNOZYyxw/f+gKpsuWnQOB0I5PdKCQibFMvahxB/qaaAfcZrXVrysr1fSF
0ehzTSQqo8DeuOMKm1EgFucowfi8BVB6pj/xchx3b+gvaqSuO1IzaQ67pIq2ZskcrxJkQkUdmG/V
pRUnnpKSRB2OXfUlzNbEqlRb5XY2V1VMYCbgkmGWoroXFsLvyxaLzSSk7XadGbbYxqhL5NGXQwNe
f38C9JWIj3qnhJY551IPo16VLn5Ga83184q/JavFvoHn7fikVvlVJ2ESth563fGTh5JTPuqYVZsh
T8ox+UqCUoDW73WpIQyaSwDYNiFicC8CowrgrNG3IqrtTqHIsYphS0MkaWtjHKvRx40JarJh5cbP
C51CWMh0QLWuKhStcxa33tUi7/CMXCT/2AsVrVypaPxUj4X2PfZGFFUEmVtgFgv3dDtpkctI+jj3
RunmI9unCrtTC0CWcdgItamFva73fKI2D1szllkPWWYOWvenYVF8TgFU0YW/KuArwxQnDK6Rk0kB
CAfWx8zB+HNA+7mau6t0oRkd8uHKFJTBBPpogyd4D6JbBBq4udQ2NWpuacojsZtWOGVbd2V7EM9c
n9OxzT1Q5bdYj7yBAMbdzxO2rLZT/BKRwvwMzdOXS8a/EFG4cub0SrQp3fVYLN6GMgxSCSlf/qlg
R12VASl888GwrAxTvn1uGbuSTMvSvheiaJQsakNbuDw/0dmiIYHFMLUNpJxIRrpk30qPZgf2nSWv
tnRYtpI2C1PZ6zTlWv+abdKA1OOtPpMDgEaEeIfTSXQ2bAAiKMFq3U2i0+O1bVnbdUvvwGi6Z3Gt
Nrp/8CxO+N3VCGMVfTCTBnDYZthCp04Mgvdf2Xed4fx+hiXdWtD7IocewFEk7SZcNWAyROQO8Q1Z
VT4hKOF4oZ+ripoQLO3iACqj6oH9R7LKbNP2KwKnq1klOFL7h2+cbC7FmfAwztiTZlPfuX3KUe9a
FGWYZOL129o+tRGrZfbqbz4klZI2u/hUK2eBOm2rJNGfnlCEzGYZGIZsDIKA7W72IwpUa8NYYzpg
3/Xhlk/osiR25vxcWKMGBggWKJaCItOita9hxF1qIGBvV2DzQc3UmT3yxBFbN/TADauKPJ1pYkTF
wZCfHuM8xdOAJ/SFNXA4Yi7ifXWLGY8MXUTSs75H6e4TY192YCt7rg2zm05nDQ6iSRUvQgav9yf4
ReaxKpGf2Tq9GSIuNu9KTtPVS55zfPtZ4zzEB3nPIvdMGCkXallLmmyyEQHioO85ReL7Gwqqd5Cb
Ts2tOXOmohPxVhKRVeXJsnStTeBUUhyUUzrz64xc9PwphrPSacop4EKskyEcLdQQRJ6WCP3wNG0F
SC6m0+ytue49/sc8nRuMdESoOp5y2AyLSzPdGD0Rm6PZxe4GVgLWj8DHii72RiJzTBtqRbPqEFDx
RuALC5n33jEDORxI2Ri6RNYzYQM9YydE+XtkHE0tuvJLJ6+i29SQkQT9QCWiP3IRVda0+V04aMs5
vbHCu6OBDqOXcofwfeTOExlm7i3ipo9/015riTd0kN2LDRKmpPJISGNLF8p2VgncYqugC/btFPGE
ov5ik3MIgWidxEqGeu37Dnq2WPu8kP8tEyf43XBzbwSWRiVVuzL40EfLIFE6LkewMweVqq7C4eRP
ONm6x3v0xM1ZgjN1bV6rYOlex1qyy7kr6eDK4zNeGpS8YneMZ6hMN9SrEK+nsaMUeMpqmLnouUJG
kmJV57RjEEyV2ccqc8fSm8JptI2HUGOb+LJPie+Yb8HWFA0ukCYbhAf0sLmvZ4K5iPIG8E8cjDhD
6PAKLqGDBsOmfzb1q5FrVBDq8e5DM/MR5DvQr7+SNDMArQVv1xbkGTBuJe+xFpofpT3nZ1pgdHcw
avO3XV1o0QoZiwayhw8P4covVLt6UgDeQ3JUayziRy1tKaySJHrTrLxQMUZyAqcJyjnNh8NBMvUa
eC1E1jXj9K7aGuHYkuZJB+IRe02LdxMwKsfQZKqDK8G0/NTX9e8ITY8O5t1udFPMfyzomyGzYBEZ
411fG/ta4rUD9ypcv2jvtTemGNXz9kCfwkG8W9fOy3vRDN373IZhJPmy3BI1H5ucPedVBGm/E1SZ
tHNHnytqx8hjDuL9426E8qGPH0VZV4fHwIkph8kxN/XbGpsXs3MpbqAn3ELixWYiboOsGYl0jFmg
4JK1hYggAcXlHnZriuKAep16oC7xWQdIWJngSIkh3+vAdVh8FtbgNMpnTC3dA1rjFI+07wfOCrYt
R9f1eEw2/io83cGPKPPH3eKm0vlsa5wmy7kPY8gMDPF97JNIU40tGFN88iGWt9lFykZ7T4Co7hVb
ghZtTiMMJkKyEsEw9jxaMrIQXlSW0FSZxrf8JGYjYbTlZLZAUoma18fkhgipXjtfxFbIRltKH1tL
A0FDMzg9S0TJUXfMIK/k0u7bq3RhH2dgJ60HwyHhRwNGLuBnAynX7Hyyev+li8Qz+UhREni6EvX/
E4RSUVRcdbQ9INreyFB5442TUPI+Yzn/39f1vxbKKHOLT0R5EHxQDa8VbplqrNsHwUKSbTTcyFOr
4RO+XgnyTT7bTXW2yTOMM+8LHwXKNrm2WrpSZ7EEIYUaTIeBhJ3WMpnWOGRvUE26PBhjYMn+jomi
c7uXGP2epOk8LK46Qlw65ZR4yroHmWK4JzqASeWfBSVVsZAfZHbCRSw8Dy/BM1aUFEZPZJenUF46
H5MyI+ZW2o/GuGVoK3ZVyMApiZ6zTd4yT8krznFvKJKg/+aZzp2ZpuyUeN6SM/3sMp0Jn6mHkKtO
SAdXWvxPgBIRzeAh4HQNtOo2bbL5V2xgmQlLelWc6kgr4KGbRokUfVc6kbjkfRA61wxUyQTEEx+C
HvsPnJiGhRX/l+lEuRsw72I5LVKh9SWwI53FqynUEyNGA34XOoUXAdH3MMTAtiv/JgYZWnLZuM3h
PnjmWDe13NsxAu9wQ2wgac5GNFDmKxmu7kpFrwoCzVdK8Gpz2zoEQ37go/re6TgRh0wDkjNj2hDF
V8B5+eaDtqQXhQDZfi/NayPuW8yJzXb78VLg+93xkGu8LDdZZiiaYh4XUTpGvZvq2Z6aF01MilGU
uW90g+qZRlEww3qIZM0LvcuLsg0aNDHE2NJzGRp3vtjS2mMBnmB3j8m+ExOU0tRiXWpy0YCjCQMn
P58/HlhJGlYrFG6oaxUKXsPrz7SZrcaIUjqGcqXml2hygRIx/knqNKJuzkvIGZRgzlwgCGAAo7nk
gmcrPJRAZ5JWbCqmMJkyhoV3shMxDgU8MJKoj7EQWQqKbI7fOENaMtI3Qtv4eynmRou8YsEzyoQl
hWW00nSluRfF3lqiwvLKhk3+vrENJfcvRQHXZv1orThwdjM0+xpR/bNChDK986iqj+X+MLKWq6wX
U2v6P/VeArqfMaUOAFn4Xnj1v+hBPA047JyeBPjUw/Q3HexQGLY0bwDidFVDGwG+9bb57HaIUiN5
r2UuUK/SrRm7ho0sfFfm++fmLq40nMi4kWqm4Ybu2lvolZcoDGPvsG0G9zp6iwF7PuB5HspvHIeM
l45lT7OXPPexBqQPJJfs4LHj1cl00w0Co7Bx1hnS6KeVJ1r0GXTUuDeNfkXAlbXMVHfrp/3EUOjm
rCCyRJE8CO8vzh6ANuENX2fQtsxokDbJhY+OaTx4pUdJEuGuqdRj3hEqLvZmxtjpGKlHR86sfMG2
59JISQdTcARFF14FCgCF0bEaCsCSjR68hrJ1Nj4XsUSSHiikqgU5FjmcIPVi/Okx4AakdCrvkh13
wksBf/qyMCwjbecW94f0BsExsRt+JYLZPagI/eLetmFvX7uB3PP3BXbObwA+NlvHeo3+BqfW20jb
XVD9qnjj6QVLKpCDUCIax5DLT1d34R+DWORBjoiRMKPaGSo6tGr4PfmrK/7gx3eSTaNaJOq49SiU
pZYNxyY38dyP46ZQDnyDp8SqKxCKNM+/EuH0o0xIRUuK1mSMdH6zoHL2CBbk0N/JkLeX+hSU9PrB
T1WPqx7ckDEGInx8tTtWmBAyTNFoRbSym3hhfStI2jJcqPlKc4haFEmSvEZYOxlR3FIJFJw6QxUy
NvDFCsS85GNay+OWl3N2UQaLJi3/2ZH3y8KOFgzPcYY/KyOhOOBU4OzlQCf3AfpUUn595QAdocST
0/r0k7tOv4YW3tKq4SDEUmSexgrVEXVO+klEmHUQk4ITz0lVq1C7G7fPyNMNi/Dscwe24biID44D
KPUQZw++qD0VEEWxn8LL+LdRzx4f9gl3sZLWKJJo4m2mcKQNOiUI3MxnBdKkYA8Bi2W1qx11USqf
zgyIcxzbGbHwky8IxewXeeaIb6NFecTVUxzA2D0o47ogMC9iCOBHV5dPjqu/jzmjmypypVRJmqH4
gUAkNWm9ViL2p1acBfYprOsUVIlHD7+A6VEyMQc/2vgdl2WUgKtyaAdlQLjfu2mxQ6zY7lu7Jvw5
sYqR+aCbe2ZfOHUtXYvTU0CHTzBLULDLAugvrNNTaCSPaCMejXzAJ+sJHxUyU9lBIhCbfvfDSsG5
ltruOfKrCsLbFobBSwnuWBYis/0MSFDihDke68AR5xdlvFsM+489YqeP61oTSsQqYG6c1Do4ikuS
GB57qh2fhD4jf3IhG41viuFP8yVi2AlRPg7VmdFp82aDYo5igVzUqP1JKVMVwS/iIsNRFKK5DyoS
RYTzLYrYVZZ07S18roCQIF09c172h2Otf9aov5JHRUC9LJGKVU+LXXVUIBOke/EK3ptQHQUTr8Er
r0+d1vq3o4FsoXF5Y/GuwCLRBV6lbhVe5j73eW+KKlLJ5jS8bEZteQHITRP/QSvU6NQMgV32lVyY
eZr13/mx2LCX1L7mqbOGgWLRnYM2hWNodB3YzWexgOrFGCW4qgMHrhMsjgjzpQVPwtS1Yns0j9DO
ndiEfpIQrj+P5aVU9lrc+BslRysPv2/3JanHpZBtlcVPdsQysx1fwnDvF/UH6fvuIwcQDUSsrEis
UEOZVN9dlu/V8s1y24+phkZGStpihW6AWbDLI8/KSn3Sh4QqNLsrXld2V+8dHWNwl7LZbhH/twAC
471K5h6xXOXSx0LAvzGhUesRGNxHnpfUgMItQEBe6loF7MA4m2Pvr+FaggBDqHNjDKzi7nTf8wNu
ETlLSHm4KTowC+pX4/XTROF1/zHxAYfdm86AXzOQ6CuZX/eY11p/DoDNaoXXdUzibiS1vfqy4qsO
FiVXrxrHN8IlrSvcqyjzwPXW7lF2o4MiR4KmIYZlNMbyoqDnwoiDl8R/SVo2yr9uukSiUqDO2J40
dHe4WX0P4Uyjj/oGvo9/u0p1bw++4L1GQ7pnx10zbykxoLiWvJVf1TY4oxsHloZp6feUOhLWpkT7
cn/6m85uQBB7OkxM4v7b4sIzgSVULMWOC6tApMMYnDTVQgWlHom0YL+s7LSi+RGMb7WJkWQJ4pLR
oPsWwGqDs/oPU2MnPqhk+KxCBJVfFXb3iU5rAqvlsC9/XofuSOPwfJjyHsW17gZ6RTSLKoATnNDJ
q1enJK3nbmtO86v9SFJrkUQ9V3ohEBwFO8Ekz4LDfcwjmLe9L58GxGIoeC71J37dVgXOd1RfBnwF
nsEYc1y7PMnLKg1Vs9CE5k7guPoERjI8Jbz+Dgnt2FCsYVsXlDC98SISg8Cbuyj7zM93dOwvw/RX
+M3vQ/gGGedkJAR0X5j1pwtG5waRkJSEeQcP+6Or1tv1DV5yi2Qmor7XrtdXBG4h4ZuTr/FTYS9j
K6cTuq44CyB4EovC5QLs+PwLClVEZKh+e5Zq0MkU4dXtXjJVWll14Pbhl073rHCSfxJrT0Wp0Vi2
SpfUhdXCV+d5J/qSOBhKLaJwEOvrr7ohxy8BIXbkaa5PDDUbvfUkFVMthmVYUI+LU2ECzd9oD9Vc
Y8jLQdq7hSwRXg5S5Gzjz9Li9fTdrpqU2qhAxR1IgBrPmlO9u6bdqk2AvcQlo4CVR92AVzUPhyUy
f7VRkpWT0jsLcMB9aGkDxCqVBaStPCIiJKOdOtaTqPDGwTiMS1ZMF+3+yDLUcuoJlAcqBRVkaQTk
hsoyBTCesmYDs1hHrguTnJArWkII2zQ6wlqCQOPHOlgHKOrC9IO607O/vbYvau5pguRCFCHgWLot
cGYlzW2Rtsi4jj+0gRsxf/51WdggPX4cyhx4SzkPTQVHPsXXPf1DPJ8lQnwY0RuIiUP7wu1Og1+/
AQ+o/iyo6ve+EatGJZRDYKZfGNpBnmZwaoUZ3pNwBkMXDaHMCrhCz5oLg9TT0SJQWUlSRa6k36vF
bWSrXrJiRGlkKCkPQ5Ca5WpUj34yYeEtqUaFmN2agScAy6ZgiNn+GwuN7fnTOqS6oXIZsNWj4Ax6
B9VQfxMFO+MKMPiRS7/a/Gh2INkSD9rTE5Z7zu6SxfWPdEEXhXKo/Z/9QK7pAp1+RPbSQ2BIw2i9
62+X+iiqG2MN4V6sdAAerSKXwwZDF5DQHpmPQfE6sEA4O8fvPH+XxQ3mdl221uYi+h6ADKrybhNC
oInXhubcJaIRzLZGPOH5trppuuh6u4rNCjt08jUifJyN0TtkXKtyvQCnizWyqRs2SnlockJnjXlR
baWYCK3ucRVjrxrdISZ/xPAdDf278df7fJ4eaOQ1V3rME9Jq+10JabeTVP7BB3X35E3/8iWWn5nB
a/JfprQ18S41Op79CsSCDZQYrWbnWmyAVMcgdYSnvUhlks7kZGw072Y02eMKmYLis0RscAs+M2f2
lqlNW1rx0A3VHZa8Te3LQlX4bvrohFWRIHPgbalsZV1zeBaQ8cYz3QBlHKmgjinT5ElufyN19Jdw
/b+bavU+sbftKStteR/VDWO5u2uneApYdL6pE7QusmdY36ECUdOc2Yd4JR38tmhjAegtO65EiCj2
2qsGEcgov+yT4/d3WlavelmOeL2WaSxkJsHYJTBuCiAGJcMNPzx6rcJo30zSC9s/UtJEn7VGJPkZ
wTC+jpwC1c2H6Uz4R2PVSbdXrzb8Cg/wgz0lQL6oOKsm80Tv3lfnDxHva6J16VeFEjGFZHYJ3pyA
xDj8k6C8hunCLRVFI1+uDwmiszJB0i/T7fi8GnTXXaglWtXG+DD8SFkBtR72ZRUZBzOLWPI7fJoO
Jiawj2ZOzl25PPf6Js/dKgKs9tEfhls4+YFpF3pb8NOwtFHV2Ev5+5QMZp/nwuwGQRcumMuqCpVE
Ucf52GJ+PIr2GEE3xnCd3VuChLJ0ZgR2gkepcpxVF+7o7wjosCDXylTSA/rRpK3AjXojvHWtTOW+
mKcPlF29u9xkLzKYjYkglUB3A7KpYldRyd1GU3FLqhaJ0Iv9LZaXKhLT8dPD35t5rinvR36PCk9F
DWmtJiojH/9MDkupccnXu5bUtMFb6bdPPrWn/UM9xikCmwM5Y/dyJFzoHz6UsUqiILSfc59z1W+W
80OQuIzHl7hhazWkK+U5n2xhpDu1rtE/A3tI8D6BF3Lv+TxfyvZYY4BiAg/+0KoLbqJWdFoYf3ac
mZvQrKhbtLjul5qyCt8d+bLzTAxVJe+xVyJ58Uo1alFhGfyJn4oQEo3r7k2tNQ7Of/cciuYn/T6q
vbQXnEkHDf72JhPkpNqgsvCFsMQoYgLwpObKvMRkyCmPHOysDhU7G4VC1+UkIpz69KryYpE5YQJO
ig+0/MeLCRAuxcf/TCql6egBZHOaMY26YT198Zpyo75BRpQC4oRUpmKNxQnn4QYYe7PCc4JlGAe1
7lEUj7SNobqRSevV6Q4r7Vg+4NqIuCK4AiWo8nnzpih2n6HD3qKkdssrC8gysyeZbhszmrHkUvba
cJrxTtFJRQ8rXXRU38ebCgKFDwIL8BRtj1s479csCkIVY8zNAMslevId4F6L3ENGznz6KWI5krDi
Vn+EG8RLMYYPK3bex+NMQyrlz9oIX4XiBNSAJYrgCA4L/mJ+LdU7f4X3LU2AMgXRlOtd0UVYGTIo
VZD1J/wT8lYgHnj/34yTWwHPgjDBp2Y2dhJ8FzQivNVdmJdUSdHxsal6ZMvbws7F7elLOaWGu51i
nIFm0esyUtDs5HS5cBR9nxjVIBYJfwvTUbciJnnQiYhgKu71vgG++CxwWjCvc6Cyz9xaZ7S2G+X+
UshLWtkltPrv/oJyf69PGTT+4NKn1G36Mq8ZdDVNrcm5Gbjnn/7rdqlRm2BZtna+PV82A1V19FWZ
QfSHypqpFpd01a70XJ9GRa2Y3z38LsD3/9v2bbDMPQeZpWnG1AcODsvypDTMKckpYxocUTZ6nlXl
ApgKGRfHpvHdjcTCwoMEjrnOz8gJ92ceXebqGZHMdI/4uOk463TUGiJcdhKeblfN+CFkH8MJOrFD
rrSgrxNn48oqV+biewFgwJ6p5PajH8h6ckIeEOeAVbdSEnmx4dvJ+sBaGo/QGepmVxIKALHwkcJJ
qpifpVzAR9FZ9mxFBJXel++6fh+i/pTbQqXPx8k88iGdI0UczNqRPptdM4WqSKdDP2/UktSYMllr
axAL05EnxPIOufg7bz+dD14XEdF0VLr0bLMPt7G6auUd/Vjxo+CBbxOoQOnMAV8vPfKriQbCQTuF
tO/T4aECd3AkjdNUkIf+4A4GmbIc7Wzf+dsLv/6ibhdW+vxxPB/3rghnAVRqCO89nBNhabz6+GzA
CwA88bYCMdG32rAipVcq10xhht8WXGAz5OUCTgY/wTnF1h37A3hWRQoCkiFuXv64ZL6sSqqtAylw
fTcW9UE23gQafQRm/2mbnUABnumkqiqLXMa/lTa7aDnnBsyQcR2lXAXPjD+ueZQVhNTvKzEowd99
UaO67GZRC2JJ1Z1wcK40Tl24tTgbyrO3FI5yA87JsX9Elxc/uuLNrY8EBp6SvrOj0coJsf2Okzvo
BqQmyZ1VYzmnD8kRWjUz4JAS45I3URBv7KSpUxFxt9xT260+1z6VNBsRKKFN7JD9wroWjjhEY3pD
HODup3o2Wyjo3jHlv0AGMdi1WPCO13Qw0OGFJgxv29k+xyuebt0EMlC/+o6SCBUyMoViVdLilh+x
TYYHLjEyQ1HNJMA8jzl5hs5TddkdhOuRkyaWj7CwMzbz4TKsNAPkwMgSv01M868kmDvUnG/8wdmJ
GyznuIBDH4t/G1Becskq+a82dLR/KTTg6hRP2P7HKZrsdWkHPc7dDwqmqeNjcnT2O27+6f4Jlfkx
miprpilr84mHUHO37sJuQOXiT9bp7pSOsct8CRA2YoW83pkYD3jsnDNotsIsCUFTP12uzC5kuvkk
zUw0mqnq+9jTcLaFv5VGrMasoIYhk/0XHTwcxjarHe7L36Rpp4sNzMkcJ+be/dZVSX0uv3zx+fPA
3IV8KA8itTv9SgIgZbN/+7GPwepPjKB6h2xxSFsXuRZKAkS9/MAilIc/iirMB87YJpYWVhaIvjwQ
lkigcWNr5YqpmzjpUBYSp/9PbUoXLrB/WEOQv0PgOEnp//bo+CktCMy5HZMLr3kN2scOz6+ov3sv
5xKv89I5Y9BEtSB6jttGLmduGQQgjj2jEQ9RRD4lZpEyYXYku76E8//+FMCaXSYPKeX6qgDdn1Fm
dmmC/1an1hE5ubfSDfDOQ5/VmcYw4VY0VHXjJk5GvQF/BRlbVHuuVThaoCoElEAvOApyNjdyzmIv
yQavmVvU2/tHjtQa4FFOppz78aa2SUTYqXo/7KEj72tq9tbMQTuv0dDtNvoThU9T9UyiYW1Mm5oK
mYF4EyF6d7Knimj7Cg+rO5OKNFs2/1GEHZjPMUjCxkSpeIp1ezXN2nl0zBl7hotyOXvmuUgM1taT
rdPPGA5owv+6JAB/lmOKt+pJvFhVWF6/Ow3Q7xERVOChDQpooWN9PZqPkOIyGO/qlNntqVbA158l
rQfmlqNJfG8Sf9/Ry0e0K/iUJGDL+xkn3rk6DFyxTCHtfgchbdcj0M9tNvgIss9gh+IBt54Nk4Ne
saPwKs/pZPwgHaQXn1Mquiwxfi4emIAio2p3xTYh2KeCnFZZS3HC4Jbae7BsRZ+agYv3W+HhvHWS
n0/xCEgIjWiAgeKcSI37rg3rwLycVO2AcfJfWlVO1KxWbS82uqLRAoY7C8y+8p39hn2Xca5ADV9T
9z4hbuSoHM+Ri7QzTuCjyVt87xsExKfGanu1lu2fQZxU2Ykv9AhAi9GS+V7hl09Sv6h5L02CHsJQ
k2kdqlD/CIhB3f3nQBa/ZFbSmg0y0zFXekhaMIdicw7BE6ESEaxOEYgwhmkCOUQcpPHLKyM/uJlB
T7dldgsj6u7IoKowJn1m5vxvyGaPX65gwaSq3/8brfKZ+HySvLYULfYDx7DA1q0+F8BvQHsijDq4
3oHnH4v+zHtiAvQA0wEVw2hgc0gtoIYtQBH71esWMs0h/UW1lq/sxHkoC164qIGNcKh/Lxx9ynYs
KEmlkLApqH+7k2nhCd7FP3YEixWLbJhXSiwBjmLl/29hpkYKegKuEB2zKdkOuuifJqUjzcovHhZR
ZDX9mH/rs+4GQN3TFKWxhAcgaGRlw7WD97Qk/CFlWlSOcDGaJBuS3TuT7iAYCHELwQpBSnxTRWby
a1rc2ne400l1G4WiuGmoznCXejsU6+OokkVWL4CGaKXKpbpYBrR53S2CXae07QIa9/xkcyn3wgd5
QqxU3tA++pK1/pQUdk0ogArVVdz+WXWdKNpyzSP/mXnRsfQvReSW0vJZaMuiImWXNncwuMEVrN85
zJc6ZGhOFWnr0qe87Beo8hiX12cPBUM3yY1sqQHmiYyCRmjlDqWbErY7kjVLgZtOaXzmcQOUgUhy
5RXmxbyg4XZIeyIOuBAbmJSThYhVQGhpdehBwt/UC9vrDF9k10p+yE/s33rEMn0ERQNV5NkHLNZy
lVLHRH9LLrysCq4v6PQmYJsvZMI1Tc0Z1ZghI1g+9iTsZaFk6/qSsQIo2JtCrCDpddDd2ldOWgN9
OtLsrz7oIBOCu52Ov2l2Zi4BZilWSIqgT1A9yWtiNkgh/XEAmGQfPbO0QEUwKNfW+NRBWs+PG/D2
BXggrkNW208Z+WY/QLSPPinBHv5M8bUPvAB6JdDl2THXiHqOGbiCva/rZLWublDlEBVXU4WXw6NG
NeE90raprACFnrG8epQU1W6gAQe0PibslNItIvD+kWWWPJuNJu8IEHwTxQ7teCQt+FxnDZasOFjO
1CNJwaa88udTONShmzoviShzV2TVhrhW+FTkEdUGfD96EDeXzwDjRcaQW9og72aS13/yQZm3Ph6n
1Mvrbwb5Xt0ZD+EDj3jVpwNnZYuAtzdLeSJ1UOVFKoGu2Avz/WTeVEEQzWj3UFdDcQt0/ATEqSpv
7Y9k5+g2dOdB6XA3EzR8T3uiR2T74TLfCbqWr0Qt4W4DOdLCotiLRWXuygzb55kXXET6pm8nRAPP
7zK3nGpAZGMwaL5smXl9vEYDH2VEPJUi+FT9uXuF3BskHnphJZpv7YJe6+BfxgHsY5/ma3o44Fdi
gJWVC+2EbFn471zotzCyX7War6FNhqiiwKET76VDB3sYnREYnVhYD7XC2Nd+y7w9AUA7hmWJrG0W
0uXlI9xvGfa7tjE2YJdGtZwcfSRoST9vdcErfMYRG+LRp2/kg6zr2YYtaqT7lbnb0BqeIqQfWMRE
EN7eMQcmriFkUB2QsIRxfHJCsZiuvDHSpOhuSjrHErmsCoEZ0f23uCNXAWxyvfXTo5FGsg9K8zUL
/w7APvPb0BNCVKUOJ8eTGqzr9e9lybH0zH1lKawaUoI0h3jg5LcgHCE312MG1HMywnjKYih1s3g/
fgu2hxYoSdSrhbC77sBOK3k9PPHao833rNJdyTQimm+sJ6z08h9gAnHrj9E6V7FPfPE0swZYfPJn
G2nZLCWApSIBOMUip64jT/M3R6AX7cKw7eh39VIrIrP2WyOLj2qRrFHjzKtNZp+TDIqAMTux7HzM
PGUjQDVqxCtd0hVVdMrpGQW4cVPtwhV9Qb7Tee8X3y4Jbhj9JQycfflONmMCMjqPWHDfOWmCv2Te
J6TmTX787ZiHUccdeiHWsk8CMKvAs04fN72ECejcKKV1oxEI+AdwdqVsOQSkIG/ADSodyiIwPt4j
EyOos1b+/gsWCrU2J9TI2tpszt59wW1gg+H72/Nv9tpZV20zunJd0S041e+kQxp50Sdcxn+VQTNa
DDH8PAd9cgC7GXx4WStaxFRBSuA049Ogd8ukOTO89km1UDMTCT9PKSpUXnlid2h2oyt6qYMWI9hl
c1Sb+y5Wg9bcvudf1IDVi6J75RatBdHkMxfMh26WdJ8612Z5QVApiFO1vRKr75gpnq/J4lzduP8w
DmdIElTk7Oxx+ZoZk26ljY0f9AV+UXgeXaU4BobYIcPGDGmQksmDyO7RjjKGpPaT+fu4ErQvsHI4
cVA46lDreaLQknNzTTfscp/oyb0npuXWR6aq5JchJmKnabhVhK4U+JGwZG79ECkfDuMzQTmcLjrI
tHRExxWPOpHgS8Mutg85fzz3gbukIv12cEncnrRaPQfKjVYaUQK6Lh1lBMpmukAlFm1SepjvWyE3
+OBg1M2ZBYzE/CjpQPQJnPU6s05gu9I2KVZABPywv01607hsbkclBQBuJazy1rozG5lOwUdUg1OJ
1x1s4pZZTH1do1miY5cKPzCAPBO6qWY3Ar8hIJEFJI3oV5yaMnuPxjExZfwLX4OmmVRKgan/548T
/n44EOf2j6oUiZqs+x4cDKKDTny6dmr0OwRNyOiePqSSCRKqkwFsVa4+EzENLHMPVMc3stjg6464
2S3+PJ9pfd8gWm7PSoRqafRC24Qkq1cBeHXUCmT+ywp+hC4kTCf6OKhorMvzfEEM8kkBGxbEvjvy
9+K2W1aqUSE7QRdWGKJqfUispvVXscL7vs8ScAxzEyuDi4mGLgwZuPkZ8mccdbhiCl8WBjFoO+V/
IJ4sjjzlCOllKt7n+ubPTHVNfPZsxc4y1YaR84lQFG6q6NJpxPLXNB/jw5Izik3i0QspHRlYaQAU
HDLl5/GdQQq04N1iIRJFP9wt5pyD6dbb3I4BiE0rm/v25C+UQDaQmo66w9uXjSex/CV5e5cXxQCJ
0WZRj0qx6HLiBNagr8+I/Ths3YhlS+ZRDwYzEtH6K9iSL/PiRbTe8iQ8n6VIwACPuvZb9ylypHBc
Ar2F9ypn7FYSiGLeM0cM7pK5mmkEoghrATp5fwD6YrPgutKQePYzMIuejGn8WjBFyHKuy2iONCUx
iA9BDuqCjdLUyHaSZvJcy1Fugi7vydo4M+tClTcyey+Eby+y0YWetGQicw0EU39JBQZ4Lj+F9RyT
O0hEFkPrtk+mbzr/3dGyRDyChExJRXJwoq2ODa3JYa5cz2KfLDhcnXh2UPiVfwE3jU/rprrrGZi/
TDkBTddHQgFjf1xVLFNVaei43d2i2Dq1OmuGpYBFv5pXOblch6SwPYaOFHTL4ljoxgH4X5cRgOjn
/QOpBY0Rdn8rR+H/ZZkM1NxIXWF8bhvwmXo9oBitxFMAIz3PAuZpTcQqY0SBzb0bDMGCcKWOMxD6
nQko0uPyIzMGDELEA+43ACkUW1llLxRo8nznUEpTi3RDBcgHOGG4UJqKhDBDhlqbqW0vPsOBgxhe
u2hawtiSblSBVnrmtbVDD8CxWgIirw3bXH5JOfobOsBF+f+wYK+dPDBYRqR754util2ZyaycnOJs
IWtX9zDe4vuAcrXGPM61HSswLbJ9hA9iru+UOaXhaqvj9DS7A/g00G3Mc13eTzACBIqvkFMszGOc
wgypTyR6bmJXDoRxjWiXfDZgEPooYUCbOj7aIJ0XEf2TeQRQcTwS5QoRli29xVdGO3J1vvaN7GB9
DwbtcE2ZAlW2QsZqnoi/sly14pHOz3cq00oGX0PvLvfcPa+RW5zb3NhkBFnHb4+2dCwlbNKYz/q+
GEBKXYuN58utRmuB5kyXICPNfRDVn7odfJMgQ0P3pXFC2CwED3z8Pws3fzuDrJcSg8pPmRklRrjw
18Non9e0LfuzX91weZZYPQ84ov+qsnoD1XAUB12kj6JO15DfQjRaC0i/kc0519vIqYssesF1bmjF
eYa2zMnML9RDWnLgI5XOd7nNdV9/ABRM6YmvSX2AB5vOTeWBtmFtLIEm2Shtqk5khLa1UKVcSQp3
TdcwbKj0kknNO1KfzmY34nk/zuVm8BfiAAm7dekF3ec1Uy8UbTPsGINY0clpHbXjjZG5lYUdLCIp
GbJ3lWWa0Ntsg8vN+PJcCknjnwPFpDM4STwqtxqzeO7mcaivhD0h35atxot44nTScuZCuAH1sxlZ
BmpdHyUQKYHWTDRAaJPk8aNADSNedRzUMpApQnK/rfUKecsVzCoq+xx1NAQ6yxMXGKslzFMGL4so
m9g7rtEtLMdI58uLqZJX2jw5Bg0Y3RfQ+h5FAZowWg/IQ5lAGIhlIkuBfow/kR9Fc0D26cj+OciH
1YmQhRv5MIRgBCR3+QbZ54sF+RMsKkBZmn4aIJ6fcUEd0myl1LbBFxqWMpQ+F0zELWgIJyDRAx09
v5eGbHMmCLf9MkgPDRaifiqhef3AkPvHSYdf1dNFc1MlrVaO+HlBq9of55LFzldqQEtQg1iajDvr
OUX5wXYYXZ7hvrvBYYCA2B6VP+dzco/2sXZGqj6ngupTU4sla8KwT4p72StBAsfrv/4E7sRh7bsk
z5fICW46QGQT4OtIEnr4noPcC1OPfJdTpZmAFfdCdw65efs6hVzuBrIjjt6hcqBfC160bTVtvuK6
8wOi+MEmrUFnVwh3Witv/8Fl/xs4xc0nyRmcD4Q5Sisfkl3q3CNAvq+3NPZjxgHt/ED2A4RiIbgy
lToQtC4GxOMi8I2hITJciIe9MFn59qYdQ+YLiucfX2v/rYVudmb5567sOe4hqf6FWT2Scs84gRQu
JXFs9fWTCYXstUUawgF/zaatLTO+/4EMXGiFcbO7N/gwUzi0LucqMvPy+2DkGiULZqSKl6VvQ5Yg
tC4+l38M5dRXIifRyVlsTcpxRyjxE09RT33gjzDilE2tBcrfSmWdFnYrZX2bPnan/9A031QEBl6l
qPDR+jJv4/DoxITc40GtNK4pSyLe7NlKIAD+JAXh5y4JR2/6ADXb5XPqVfzlmHdEzu3Si9cCJxii
TjQ6UxbejKKad/DeUkrKlgfJIJNzCNEiKsz3L8QKfiDaMEKClWfUtyhoZA/VsCJvHi7vuQsLt/5C
QijhP/nX1aXoq3t5BpeMc0nvJXqhDfAWkPem4g/rZx8/+QvIcKjpYAL6dr+Rgb8SZ3LoHIHIzjHm
fTkdxDMC/kjL12YeazNHyx1hx21s3rF6dD0XUBZod8f19MJ+D2NT6ea6nhEdMsy81TAOsFE1fJhx
tGgbfoOUtwYftSGLMTDKURCxZPJxBqqku5gMjGOM3hXElWGH9wu9Ac1o4hVMgsvagEMac7r3DHrr
37vMkABiCazyDV5kEm3P6qS14myaBjnhnLmg4jFq2WlXGb4ppZdhIcKpW8ntxcONDvyIf9QoXsyS
BDCXb8X+Yb34ZA0QeGl3pxKgu7ZdWClmkYyyJPk8Gs4Ei6ES1lmm+Ydhl98ZsuZKb5AYa+Hf6k8i
6RtljXc5ykxWPR/JiS8ppRPLQUyKocx8vAT2eGi9xXCI2gusK71pLnmC9rinBOIY9oIrrNZfO0bK
F9QMy2TGFn664dPL4ebxsgUU3MinQIqPNZA+RoKaFYoPTjfRrHRS1nttVtvj6CV5UjiGLvJecSLA
vq+xSNjN1Z8DbIxjc/3CMHOoqQ5yhKYz6ebeK8iWJR5Hf6UA7wgsaKgJ/2sJm5pGbvFd6VkFBZ/Q
BZlRtUsuyxKA3PpnrCjEJfDrp0nue80/M67Oy8qnklwTspahTvt6tEYG9PqA4i6imJx5EmUlq6jb
oWY4Kifq+QDdkuI78LACawAI7pvGUV7ADJ+qJLhQ1RykXNubS1mzhUEgGRWuMEh7mnJmLf7Pr9tw
fSoV5dgsjjhJMFEZuY/9qjjyFlyrRE7OqLsdUwY9IBpsTti3qsKHFGmEY2YN18FOxLhRnEQM0tTy
gONNMVt5IrIzf4n7jbuAkPZHZ5CjSDDT0c+iTjGduN+abXfXpXfeAxJ3Mgig4yodOXvIWPSWALXL
sD0E79s13qzceZzhfy8OwwFfrRKFyo+QyeWsuKkWaVS/Z246dg/RpNtYEGBCTV8s6tesj8xEqeD6
ADbn0skryxnMess61JTCRkxBdVyUk1B0RT/xE9HmR8xTYmjCnywjzxgw2FIru/GAat3whMUSxU6v
Qoc6CiRFswHSTa8R9GoDHzfxe/O+GLyi0RkMzqvevIbB3nZyrIbgcbsdE4r7PEUYid0v1Y4k2yUq
JsnPQ36IRYf2whN9pT0+PvwCDG+IBM0c8ptkJxaU1sLrudzUTMyc4Whm+aX75rm1SgOUVgj7QC+z
C+/wyjHB/D3HVH+3Ee16m01LcSmxk2q/BrDZox37605tD5uO8kW0nHN292AxO60LZkt7HSS0yu7o
MvQ6TGKG6V/OZtjsmeua5rOX5up5/hO45R/OhndqetkmadBlYsf4H+1p4354pF4vLQ/GOaZNFyIY
O00YVDbPqNrVDS23GCjNW3M1PnCz5PeWrtXZOOKSyMcaXuvtjtESNUSaGJom+wmWU0+jRAS+dYjy
kr3YqTjx59eldvx1e1jk1ihAfr1479SwZpx06hcYFgce7mkwm++VzqWK72X+ye8kFQsk/bSgcYQk
5F9UpGpKgGOBV1p8+vIKEoOMWwzcvxXGHBVmHavMzUE0DyCsSFm6xC9Wgo7nJl4b88xNJxl9Xmv0
agzjQLJK7FBPY9yOXGKiyqfmodqglCMb/1DTg1K1e6U0JZnu4Wh7X6skRVERZCQru+z7jn3kkrNL
fmD5lRoPlYwC3qk8S2GV+M5yX8icO8az1OodRe0YHSEya1+JSQYGpGTn9lhuHadiNn9BY83Nzaqc
T5wYqwtwFNsTA7UmGmdVdXBKZP7GC0o733fAf7IEVlyXDYSxbco8OLPMKxO5zHPMrVbLWnw2sO2L
rR4VXWVvBk8p7aWUAEr4DZyrF0cZl1NgodDuen3SHcGnu0oBYDdiCbE31fNa7FxtZRM/H2Hnf8Bi
ggwQ44Ac5TFNcJwxIr4mKUCqpWfsVZV9EtmHkn+yCqSf7DvUUdjiiH1TrBZ4X+CNle6WAO4JxNHZ
6WpkYGfGWPFu02BbePJ4eLiko14vmhVUT8wp+RT1dC4fqWzpSkvgJNumwNOXkecwqWN/cjN3qJwh
mgJd+FFV6dfaNih+V9m8PZ5CVtqxNW6r7pBLAzTFTBR/5lOXhe/waGYlYGIN1l4ps5NBHoGH7Cvp
wi16RGMnV6Qfn7bzGQfruZYNPgxKu5RbihJngs03JQLuGs8EuviHkNzSvNGsMucP7sjrzUH7BlR3
EdjeLpee/R0Pxg7cDM2p+Om4WxloUSbQNGiiPmPuXPpeEdaoL2MJPAsTSeQYBAxQSagdhtx5uL+k
To/spUtaPK6Lwc+1Pa3bL7AQZL3Ozhi6O/lh3i3o9mL23nsi9mR/C60KLeu1Lc5gL111qmiu4mnH
+ivJnR8sFk0nkuvd7uq0WY4x0gAuvhWl2CymcQRcS+J8L6aGGIgme+hrMQRdKrjwcI6qiyFQUtsh
uBfpgM6TXd2q4vRDsBpK3Oj05XxC+tFZT3vrKQOdKseRFTbCI93Per+QvN74VlGipKYxLUGQ2o90
lEAIdd3a4J+UjE7g4f16z8Nvg4fVwi5cdoehJRxroF+HBl1zQAAD7Xw56paiOwbJ/CApxBCh9j+R
pP2g4XjdkWFXrgwQ2F/+kWwTwIFstMsClmn7YH5ucw/A/EJcFHda2yWCxrjYhGFdEOjLZgTkHHKl
RstGK9dVLKcir9Pbjos7gZH2yZMTqNhV0pRRvmFMbqM6xySU53iq9JBlfvFjmOT2jwAVWu6OUUbK
zWkFL/pS8OxRDudOBBTB+h2tSuRsgm7/BzMv5zYVPFBl+5NtuJ7FGRYEOkJdiMDTir04koTNfN29
C1SJfolp5wDlGJastEyhHBPsz8YIDhxSZa/1ZWVdIg82Wy9VbWH+jtZeUEP4p1PXslK1TQKNgMy6
auWARovQ8+OP/TOhoqKV252bm9BRflhhYQ6L+kWxAhf6jLrFVeimgK8VWNDJmKYGbbb/9WnFYL+n
c4tN5jDY0JPw6aQlWx2+0+8XEChaR23NbPZ4ApgXLWr0vW7FLMq62y5Bsa4Pu3FC3k+1uQW4XIaM
J7ZYAKCt5l9PdHgNOtT22sOFDVxoUVPlvdIfK09TtQRnQ44yI282+JvuDLTINFlemNkixvVVd567
2SXwHH8lPjAXHo6xszJqaiKNsJNykvCVyziCmLbPy92+4WpRJPkVTl7DsHRr4mO5wQvXAqqamCOU
wbF/4cekcur8AAtaIyBMmaWKQF/4SNAHEl/LJP3+y2a+UMb8lOPxyQpiJakhqJsH1D+NTMu43eY2
0YgADcrt0eSdcC93Q8ZzwhmoMerx4hgN3cjtB4/QXYWpNnGA7IltiWVuC39IMa8fu95mXGb2mQT2
A45LcXuzJ54a3/iam+F3wC8CgXTdJ7x/7iKwozm0lhd0wfLQmUVsIytkZAwh0JUJyX+0jzsaO2Dt
Q8GrCTJ4K+8ugmwZnw8qoXCtYTNyKThURxwxgelbCC8qhpIdWgUs1otHAB4fJKau6UId6ijmNbIa
Wri2xKNEf6ttNHT17q7CRgZ9RLk0m2cZ8Qq0XkkEuBMeJIHZ11RVGqX/R+eWe1Et2Cg+Pfj3cTTv
bxDlSWMYvYYquFyQ9+zNsOCQqGmNBGKcq1uBTbyn0xG/zyl6VNU02cDd/gx28FdbwkWC+cKvEnOQ
PgdRg9GmFCbq1qgJe2FZ1OOeX8rEVF3pz7t3j6t0KpdG+/sDbXuL5d0OyMvE3U2m7YSDOaNRn8cY
q5DI694exdf4Xy4fTW4CGJScVnDX7tKj1K++rSGYxlzOJoxH4Cz2+kF6lAwSS2ZDdUOy/NVUQp90
YPWg8iqp6VzhWiySxDvg3DDAgukJjXd7N7D1CVzUW4OZPv4RZrlU6oKB6Ltq7D73ARPH741p1cMi
sbQKxHjJqY9vHR2+ZSv4MuUbK52QsmiWHZQ8b+oDF+DbhvkGlixLJ3Iibj9OhML8wwo/in0vIVV2
jHi67Ey0V6rweAsAk5AvagrrKksqQ7tpYczJ6uLXbTg+K880/TiioaMxQK6UtYKkqq23gPSgToul
lFX7KqVMQOZ9qLOZIUh6dH5/M2HLyqhfKnbIfceRSh50af7dF3bRzRq32vtq5TnvgGOwxLxLHp5A
oWP7mY/MU9teRtB8ZFNDzTzwXSq5iZxQGljWkMDhOgFXccg0eO/R7emAb9CazELNimCVluMn2b/Q
q5TYBg6XhNqfCwxyvU8ZoUa0MnOf8eOP4/WRapf+P9169lEk9NBevOrsj0Dp99RUL4AcfI0eb96C
tvrrYjVNPxK03H8vL3uCNX9WsjrBA6+h+9LV3FWPWJ20NlEGW54NhDomCXPquvma7Za1eR4JGd/Q
fTIzfFV76dmtZowwHU+fepa3huo+UoY3rMNuwVvYzE0NYwPgM0YD0M1+Asnz7vedB8ykM7cWK3g/
7A6Dbme475l8lSn8gMDef3rU+BXRKstWn2dgqQ0dsK2adDJ0Uw8KNvMhx0ANxFpu63QNvPjcHn/B
Ck2EwI4KC2sbJyQEUifVm5lpuJU+WkTXEFLgsghRMizj/Kt2ovKAo0Rk+Syj094EYGd0C9QtRSDV
2eKSj/apzfUINscaMA1MvsGKbCruxNLuKDyCiuLq9BO9VPnKBF94vcugFOxhWBNFVmFEqQCwNJVk
SnL64APe0c9Xmu3+hnRq1K6eVN3AP9cduud9Bilo8xhGX3x/P9CGbx69P8FJeemrd5uAKh7CKKgm
XASgzKG7m7q/lURjnbxhTmSB/UK94LHLDVC+Nl5AJgiU/ITmvL8K3brjyU5xOaA1u61TwQ4bxxBQ
DHSmGo69to/LTbgE/592SuSiopWSTGVnnz0MXCGSSV3aC92Y7IILU+LIGgXpaVGV5+GbPk+cgZx5
u/ihHf+4kcH2xQ9FAp5WxlktPJ29c69d9LZHTx9ENY3JQnV8ryYzBIJCZW7UDWN7OfzhY2oLjfga
gqx3vG2Ue423pARMUelouoIaKuxl4CLfLKUwjf0h5XBojEXa5VwynPL3jA+PohHFgK0YvABe6mK5
v55dAq8W4MxwF3dDATaFfa/nQWlImyzF1XiPh1lFthCLoThUAU9+wlouKA+NfhLZnvxcRxwTXcZj
QljefLaC79f/49Ynzjr2PpA8/MLKGysIWXWmLBITzNkwny3hurG0mg/uLthJMaTAhH4h0qphRQt+
yEbuLI/eUqA1bQIYYjaOi9GMR7jYOmPkc9JKsuQ/WSl8M7XjqGf3Hg1gZLQqn8BhBodLCNjcETsd
nk2aG6VgL6xeMJyOJ3CaKPhXqOgkF8vjpNa87+i8gtULaRN+R+yqssmGWUF9Xt0IeXFhOklCQcKx
ZRdTWNIQf64KPME3Q3/bSdv5SoThC+aVl1uHGFS1Jw8NFsmQUCCqJ5azqvGl+vxyohsccSjDKG43
8DmeuepC4R+H1PbM9+IH80If7ZktrWQ2WGio2tgykoZElAhhK2H5xFscq7AsR2ouKUeOlH5Lh25H
hq9RNuF1HMmgWbgxC1dZe+hgYdvorUjmf9/cZ9+9zPPm1wm0WoJtyx9gq9trgVK6h1prRexuQIAF
iRGHrqpXKC4fW4M2+3A6+M5A5V/6Q5U31FLTCZ7yd8mRP5lZcx8CAUlZ/Cw53zrIW78wjypWsB8z
iotP44f5/S3lkopBeNkB2zAgthyZlJIjnmtRE3zqtaV/rSx3v/HciNTXicY0RlYp/kIm2I2Cn37w
iHB0C1M64EATUDWoIstx5ox401QUxUfWuhYfXnYkwToEzjFAoAtLSWHJ5oGpXkcYGpA6Mgs++/Uf
rsmMzzK+m9u/u7nNKcDqI7VclETQ090gAfCODvLXRGlehoSWEkKY5gRYN8kjBbRQzPdbnWqApNtS
3DZ9ZMaqOd9w2UVsIJuMhlBKGJhCc1/dxv3zH3MqeQ3HQYj6ic5nhy3Y26q8zXzHuR1uNE+jdZbY
XpJTausWdNGJCyX0U/x/SjHzuCa+nuSDYcSBFuC20Xl2qjjJUY8vlKMGXBlX1Mm1UxErl2MRPvHB
w+9mzjZP5i/fQndKgtkJtfRYQEaKiiYv/8NPITYsNr/QWGtLRXSZ6Q4ocjTUJWAlu/uTmzPVE/yu
E374PO/sr6agTmNmo+DQAWOYNbr5xnz005HE4nk3MB2YC5OoNDBPmJ4hKcQmbWsjKCl9CZhxexKc
tSHP7yNPCuu/XNfGV3HsjKu9H3gYmv2DhRqX9uKlkldbea4DsWJ1JaELNfaOodAFPaVKj7BJT9XN
svI96mfXolt311tin1DMHZPwSg83N8EOLZa35VTg/TNxxRWSLUTKhkRKyXTFVYJ2QeTXwtgQuFgj
hyatBwactIEUhyFg2hIq9UnFU/0aLAuPlLC6/DHZK9K+eU5o+N6FJ61Ftnun6d1CKLmaHK9cWeDZ
9BVwAJgW6oWUR08lH1lwDS9k2phtcEFVf6dJQAcliyTnEMwXqcpJANEQwCdCzoLJdL8O1cpWG1Cm
GuT5UKV6gMtP/HtHKUuryszlyNbVdYeIjFJQZOu34kMRx8PC/EQE9tNhb6nY6LdYfE7Mf4BtUypT
UKlQC/urF5mO1j5sUKBTVzeTnCJLcDxjX6oaS/7kTdfdSBrli6fwmZHh0Iqo5Wc/L6ips1UTrBR+
KzjDbnTiqXeEfqKLd5CPvGf8NeJjvvKQsGXNwmmrI36/dz7Lky/1K3cbapdaohe0zwNzpvWXwhni
62t/jBI4wy0MKlaYuppKqDgkjkeomNuvhMx5f3BOLPXz8nI3cOxQauDMy6BKyVDonOjUnP1NQpqH
1xX5ZbziMHl07unNZKgoOqgnT74hh+CKyi1tLtcxY9OiVMDEyF2OwDQPsv+Of+3sWUXaOMo7VhPU
folS+zh8bFunhzakOpRyqyCfsEe1t59OV0bEqfE5XqbfQh1LKIDENqxpeTulp00w2/KpXCwj5qlQ
iMr4un8AgZxhXEGaZ7jtJYzndSOUOI4VjNabaCxQnvCUFaBpQSZ4gJ3b2LrelrS1ivWTAkWTYDpx
MLRI7WkndUvXLwyU3UbohfgFS9blgemOihA49OwV+92gU5P1UwdksfcYx95izmPcnr67d/XlSDCm
qv+1dT5wlw4yvgaQSkO6xyK8BSvCo2LKF9kl4dkkqj8ByLJ6J4rQ67K6IHKxhRJbOLseQC2fIaEh
jb5MbehHfw+HSCJUoVmmGVe1pLQRUu8F6OzlL5umpRsSBwVN0+eb7jhdGvuAWocQDd0hb/eXI9zU
MOTzGHBkSsEb8Ab34eZXHtPkA0pqQxEGMIU83tGlCjL4+qIzQBu8avR/5XAD4TgcRW38b9W1QVaY
4GkyKMDJiJ9/cfbzJaplyfMEksKacFbxJBDDSYsSGDRZnZWbqTvpotSDtutpI/hUTxZsuc3DyVGT
aneQqq1l3hpkulnJf25fg2lxhoWPinyyGrl91wAGCO2UD4fiwykZzgz7ustgLTJ5/vW29JrA03Fv
ZOKylKS3oWAdPQTjHIHvrCIfwz6lTfGUwNoJVDvuQr0QNoigJ4cu1Jelly7amzQkvj/PI/u67rFh
DNDMyaFh7rkusUphATSdzuv8/U7u1jIIx0T+RzFly9P/BPZTlsvJxprFPINR4l2/NMefUUC8dDpL
slo9agO+DFov0M2iA12vzTbMHdHcsB/CBJ3UkgQGkDPi2Zqc3Png6ujpclXXb19AaHgAXbxMe/Kz
i0w6H+DsVhJdXJfy81gI6KBwdKb/vhCNd8sfHHACdmxeL5qocgbieBz/G2PerPQjfslsF0Z1OvTx
n6LNRSGLfeBwSpoDF/QcvF/0+/SnvsH3R2EHrvWDwsaVA2Q5wNZodtLF8BuxBJ3tsNdNPYK2m28n
fccOvN/LBd7OBWqKQ+if3pSLNi7YEjUvFREQA/yAzGnFBr5uiaeBM+V5mTqun1ucwAWnhbdASpvU
T1nPuTeYafTuK8PQYAFclDPNzvwp1JTB97ExDnwY7i+F8iDshYAJoecvbsIrqkPVyfUlzKLRhO3g
y/KTlURL0gudSVJStGvshs0soBFZ6SmAUrNYCWDW9xdS20OmsPHYG2Zh4lTQ3tb737FSK6tRBg88
s392GCLSdSKDLn/YkERzR3OjAjWtgn4WRSpZ9ZC91yWOGdXkuxCxJ/SBsLmtcovJ8nuhpAniGTO8
NGHjI2AdqCXezk+KHneFF5D5w0lCFnD0AyiC1gOnyJgqNKnATen/w91BNJ1NrSOOhf5CLBhFxRIv
nkieP42XusTiDb+b/QlGni5htVtN3X7/nn0eyEUmJm30+XvzSEFfo1mOTilngGSXxhJKThBHIzwC
A8CuKHBaLUcdepAzo9EVKRxNyQdyg0MQc7ftux5F6XTKnxjFm2JJ4oi0w8sA3d2IHeElvg5745hU
Zzc1lcS7pGiSGx6CmwLWyDIyhbR8PknPF7T2s/nb9T0fQEnk2GcQ2LwHDWZEi6Ye3bGniGxVwu/F
6T1hQwdytjaO3rQHMXZxd319ggMUijSSDmJnLEvK7cgXh3bi8NRk5IO+QAadpH7kRfY/SoXSgbsn
EAJqTocZWOhmQKE82ttXMH3O7S44ZjVY5N2ZTvYdhsoMsIjAuiFEc6GiLKNzkP/B2h4QUOqq9dhA
CF3G/LNBiBBJOQhRczNNYyrnL5iiVzP3Cxy0knz7u2GuqvzghoivAkc4BrQqIbtONOfz8JRIM8Aj
LvbPy5alpq5HCoGB23tQxGMIPw9uSm0Iblu/mqRwsdoMjp/vQzm5OeFkIMUT2bm7Uap4DCgNYJ82
6+NyR1B+TiOP6Z7p6B+zcK7In6P+NhEEi6m14gzvf31NPAeX/9g4+SBbeGQQDCQQfWbqMGkSgNSQ
48U5or7DPWThBIi06I2zK7Fkg0r7SR1JXrHWKrQfOKZVcqiEzeCYvn4JaCeiyaWJplm6fd526NUB
7v2CzL2nM4tGox+h0xBipEpMGT50lZjGIeJOkuNikfO+wIGWpAqCkazxP54vJHmhUKC17gDtHfXW
phbGUrU1xv+VpR9RktI2l39nOE8ztQbsRh8Fmn64H0sBGksRYEHjz+RSuelkoqvx8obvcGfnUA0P
6FT0V/i7EGJg0Rbu4aNCmiFiWjWsvKtP8hCYr2hHXAX9mEHGVE5tuobrzF6dVMPFP9d1s+UTtwih
qZLzbwkXXhsDL4y3yjOXEjoBgWrkcQfJLPYwedn9LDM5wcWfk+5kgVcF/NycnMxzHOcPABTJMtsv
v0MQMRIwj88w4RJRYRDpzLlRdIlSlS6P9HbHXp9u/tBtDdiQNzRIjsKiqOUYwC/3S7R2Q/3jl8F3
oUNqBNQmjj8ZQvG0ZG288XNeD80WDylSZ0xB4zzpJ34vS5wVL5mRR0yvE33Al696Wa3qu9yZh/qC
vSiJioqx7TP3ayFn/Af60kYLs60nyvd5PSWsY5M+2y/1dmUlTlvjoFBGWgAAKNt4/c4pxx3tjKyb
BNW/4aVGC1DtxDvOIwbiZJ2qbAIuBZXdWRT4LHi+XTre48P+wdkw+FhtDwm4NJFRvnKPiSWP2XX2
gEJyAa0ErZqUKvilwxnZN0NDFCVeL6+JVKjIkLG0TUpnAOOow+pWwwUH6MNo5a9/Au9t0DuptzqY
F6AdJqhKwDvLsnkaM6Xh6wrI3YMba5jsDy7hIhHUULj8i93B2PbvEPIYQrzPIYh3s1yEgkXH6PTM
iw4MjZwQJh5nkBj4Frzv8bXtlcyGYpv7fD2+fMHsGSzi/t60WwHAH9jjl4nJ5UHU0E/rrFX8ujJj
eiM4szUfxQ5WIv1TGBwSMRUwddZOb8TaSnBwoCsJqQU0HNWFYwqzQkSohhKXYatln9eB6W0UOnva
L3SwSP0Q3iJ3/3xTXDEAAnJBNpXi/FKF8NDQbpGfvlnAiqlJSvc+xRTfif0fNTeQ3FgosfjeyZ47
2I2qI/SboaOz+lQGsdQWiVDk0a5wom8SB6r3mhiTNUfioG/z1E1Icj4OxoDBDKIdbrJJB3/gdvdc
Yj8u53G/fcxUFovkgaERHlb78eTpAsH0SqFpUOyVZQXtKv6/DKfIaZEbEOesp31tvC5L/agQcN5X
KbvGCy3Ej6bu+kGFu3zCK/PFbx+dqKGzfOe14ZfvkYoG2qBgeAzpIhg8UgD1KreOiTSvEPtwajqB
h08roLrP557UMwkOtvwTQJO6gU+Yz5AmVhtvV2f6vdM4CMzcyWn08rBadw1tNsaHr6prM+IEAWMr
Cw5Oq+jE/JP2SkjLRXwjH2bINkAMh+wDvTS1Ms4pRqhtP5x57UWIjMAbXXaEXiQUn1/tJT9fzWcZ
GkucEzBrEi678DcrJynSBhkoqaGvRTwibVJVtL8qfM/uDF7LJClF/QzhhWazFBDmtvPwUnfL8rXa
Mv9gN1sTEaRVGeX0xZjYP4UWAesjFmnp0rUnYG3nAS+6wNKojKQ3CeDA5aNBIGc3AyljFNIWc1+Y
U+XAawAwj6Fcf7rjwkIJPhwLgCRaK0rTW/q3IQ+S70kd1/IxLpr4O+XhFmsRalu6H0NWtv0BkBVC
9Wgm7l9cOQ0GiDqFtiKh1m98ViC4rAg0b2YdAd9Qif6Ws8jz3zJ3HGgnRSZ1JJ7KNxxVGtlUo66c
IoF3IM3NCA4mvGT3IRb985tw/jVb+LMBg7sFshaiiX+5eLmPvs38R1k1L7zcr1DbaH20nopKoITv
Cs084Pj9h8syjHNg2SutF/SLiWkDvHNI2ttTaTb7HdWk4FIxxjxLbZV3syoNWJCW/yQE4fu6KRcI
r1D/IH3W2yyoQSa9mo2YuVwVUZLElZ+EyV1JVsyjUzlUIt1P+7ZBuNsAitgMXoqf8m4Tq+hOP7Iu
CkMRzuz3M340w1k3b9CMiWbqaU8AKu4dtFY2mrvCnj5AMuxkbCG5Ld6yvKkyuUSR5U2IvWUc1lhT
/MsmiYaHCoqZV6jsg2Cu+u0FXK7ZUQX4AAHg9ugPssiPauTU9uWEdQbM274OTFUg6Vckx6nJAgWT
BGcmVNt0+KreT94RXvgtlEv67adiLdImJxHFVrMDjbZpcwom8bQwpUXyQ+4M1x8ORDCkSZBe28uA
LPsEQF+68d5lGORS2ZOycszAKlaLZqPwR17lY2hEJSAEyowL7RzHwtospBMnwLFXc9MWGBU2Xvsw
mRk3d7yIlNPI45Mid/jqmcrpi06QfhuYIfyZHJbKJkOFmkWVUwLyfHXi8ZVx73IwH4skqJyHDPND
1OWuOEXdoxjcMXG39akcYRjzVTStvlVqPhf74qXv5PFhb3Q9s9q6hoaIlfPAyppvGjMiz24hXx99
+jQM5ftz/ciJ3JbARGlmhgL9wA7/8GvP4DfluJI8BXMACgVTTb+nJM5Z4158Z2N3wgmqmfsYuWMK
h8F5ulreOf3/24E71+UE5CtYfNVIkIn8a59O6ihuROVuza5cD9PKGRJE/hKYaimJOLcxV/LkklKs
x+9uBRiSDvbWLI9uIvbic9jHkyi2MEElgldwaI0CMaM60HbqXwvoscZjv3XPo05e2MsZ5iNH0BKQ
A0+dFcsTKUgcRmDVjpSgOiKt2fY36ftdcpWlITlvQ2N/DAgkDRP0OY5w7Qvm3I04IywGAq2gTS4c
n/ozVMwmyO19pEhEczGWX3jgbIlPqh+0YZmEVNgyxYQOW7pJGzLQzUgu1PkT1dVYqsTkVHx09xNC
kTZwi/fcMIRBXI0bH3qGlsR00eamkNmkciEHNoeVhsQr6SnTAleWFZcwCMGETBn7xFMDIpkQsuDU
4BGKhQu0t+kfGDe8B2Q2iL1/xApoXOVOJ8pdQ44GVwXwKPf2inLFnmUzv5Og/Fv7N+YaIrxEy6jl
99keNbr73dbb9BqLne7Q5dZzIbpxTlijAClwtM7cQKV/No0/FkwZFhv15Lu/yzxKAAo/+sZefvRI
RN3QHUw8Ms0pQN8UF5gkoCV9GGMx2uXBhK80c8xwsB0xKp8J8mj3jlLX42GriF0QDi6HSsxxM0qN
9vbI7wnZAVkNiCwVXIb3dfkygGWLraQUqcG25MLfS5iplY9DDZLJqOePMSy6OQmasPC1w8ZAval7
2Fjj24dLO90Jmfx74kQdlsbiE4Is94OUN48Yu2f1Z9/2BAR5Ev9Xbuqr86iJFXirnW1M/LUG0gMk
nXo+buRjfYDKhYN/jFZUdwb38jrtgjzOypr95ta8cblr/dfdEi0k/wryUXaDrKs7tQDIaTRJ6Ykc
D2RqJ6t7hArzmvgRADU23Ibzw3PiB+vT/Q4gECG/r3GKVj7AUJJsEduhKlTq/xUX5G8DKcwRHxZn
XFxC8Da0zlrjIPm0EQ+XN6AKQbce6py4V9+i26KXU0gWD79XdbtcGxXORqLr3OeQpKXGqgfx0AIE
agTsteLGw6tC393Fo6J0lroM8/fsD9TRxTqZv+WcouAMrs0wBaP5EosH2yFG1as3qMon/odjLjZS
4YzIijB4fIWT72hyW4ihCNWvz7EElLBYJxVKo6osVszAtN9odQZLqNOeYI/LKa9aecx0AUOAxBJX
7DILhoj5aRpTtepmOWnx9HiuPzroOpdVmeAKejdqKz7JTUF2I03AoEHweCRA03mvODy5ZeqTbWnT
QS8GzcqfTH43LN5LtAdTgW7jPyYG0CyPBifyd+A5tyJ+mjqm49MHeA473nUWuW3QrtQ/v6O/lSo8
1nwrc+QPk61e6233cDQeAN44U/iqMQ+Uw7K2ITN9UQh89idcZdns48ob0kKP09LevadcE1GLs5Tt
J1mzpM0iocRYUlMT5eBqiIR3Br1Ow7GWFsrAvj/P5iPL7YS23UDFkFXHS9r6AR+t+odxOdYpLbbJ
d10X4NXsS3rJEc3H+VdbeFU/85ZwJwJaS7PzGekOJFRGe2h2Z0ncBsyHUZESvqaXMF+gKUKCEIIC
pvRy3pr+VIpgLQkiRbdfM3X3g7DdC2AxL8Mu7bdmTn+1i9kO9/bcMGKvOdcJQP76Ao4Q86os+H5j
rp0ZlVXX5gFye2tra6eUeO3MPUJK+j8FT4P6KGyvvIYekEK0MGrOX2+gWsykQ5LhLVJlu8Jpy+zw
2Syt4znpqIF1wtam+BxwN6oTjd8DsihGZOMYQC2fygQFxQ2JzSs3qTZMC5W15UthvRLcUCHfXkfQ
St01Kd6wGorJ7eW7WTLmyVuovh8vtOmhxy9b3Q3eH8Mx2vRLxNgGILcylmFBHJ9jHp2bNnrG/H7U
MnKY5MmVEV8tS1pYm6cxoVFOj5urUZ4SENqeol96f3el2Ug09HZR6LDREpyEwdj0/0UeLOjtOqy6
qVJ5V01Bqh99bnVPnEz9ZUi1R81O8bBExksFN7tDBg8bauJJqoeQAhoxQCrh7o+7OP+Eg9hr0lNh
7KGDTlxTCPadDUOxvxLtmke+CSdxXZHnRTqSFbFUK2/D5+Ch898cSCIb7mftux1n5j8hNvqQjhs2
vdYaVa7zXeKfIIQlRPL8ZtoONyHmqQQttCS6MNLt/iA0JqsmQFICezT2yc4WxDZa9bjNYO+7IYvt
x/5/PziKQ2Qt9Eb4Lo4REF+WgoyXDO0ceizp8OwvlOoumRptQGgXFegVcLcnzeKNDWB4gW75sUDb
f46dhEjXjtVsw3HLk2vkS6a4AUlNFlZbYaQr2vZFCZQ4v8Xl8l2qiuI7ssftG5MbcSRoUQVzk/92
po2JJ/EIjd1+57MUpEqw8IbtFJM9STMuaU/Hu6Z7IIIEZprwljEIJKUrMZnrB4VeUUo1KIB4dcjv
CzK/qheDMdkAlun9f2rhReYgNwkAGSFomu7vT78ebVxyHzo0FiEQ4AyvLmt8p3dlrARQaa1EnpeO
CadTZd/GsaoWzqX9MfuDI1jrDjBz/JkDSw1CJ17jOnduIZZ3oer+9aqMg6+AX2ePYEjCRf0eMwdn
8iX53typetwMYNq8VN0K0/mtbSQ8JsyId/KkKv6kQX1/20oMqW3thChqr40U3YOsnsu084uWerJb
qAeqKJ2GTP28spm0i8PjqPs1ju2MgxvtM6/y1iyJdnqLEeUAMpSIjSOK7AkQ2ebrDrSm/A7h5fSH
azUC896E92P1LX8n+SqXd7d15nfcFvX/LgIylmO/S9RNGOWRjCtzJ3cL7XC/fnViGTrZxXjMAFOO
eyNYPc7S07bYzcdNzMWnbClscSTQDAewHyYmYHXpsmbeXZ0KoDEX9HXk7XF8/drQW/idUlhHSAyP
dzWQtYy/tIg+62B7+ADkck7Inbfu7m0Rcz716UdS05bHc8WnKKxC1+PM6MRoqe3/F+uns15c401c
GpYQWJsBaKyqsqSzbgzZ5LCvPeOto52KWHi+nW8VQNjEdn6R3gcct0Gh81CjwAt/phqyxHZsZzLg
fFcwYcGtOAU1pLQMcTywYsD7U7VS1oohVb3WWnttu7gVdztBX4GTkK+ru1hBZpw081U8X5q/k1lG
UL9SftzqHeEVSGlExWdrTO3LDRtptUZKq3Wjbr06ghEfXRP0kLAtQpQ8cR7+AdZNrDCzfCle0Y81
ZFnd7+zlcYIWBXd324+MXlL+kPbgyELZ8ZFmbb8NYPCVNrxwHUoWFap1iDQtMovlBYW3ifHXHqex
qURuC8OUJorhJXkCvfxACDl+zL0g/X9tJKCNAbvsa5lpIUJbET65pn9q5Lm7W5td2MmYdCsnCDk2
FxrCJhR+QvFurlPk4UmGmGE1sVPXYfEYZuR8+sUP/I8Vyw0Mucp7kMCCp9ECp7H8e6/1cufcqv2d
vPMxpk5oMY58r2sMnL1F4BqJjpDyk3agepGZrmSEH66wIvgEdt7aJwu/wnpTffwl7QgaA0UHQncG
zUXOgzsZOhFD/kTj34VX//kkkOj3Vukp8709VV42gPSdUmCAy3jFwxka0LTZ3ndAdMfHEsjoX67J
HonXFmt62lclGNRywfAbCp4/2G0Ff849+UKTsniI72YFK0y/yiOGvQ+rHIHu7jUkmbtfgCY0r6sa
XFsFc1VMOVn3kKSGlzPeDPGjza9+PfawEEjajEr0cV1Eq5J9vOG4fxghXnloZ93wp01sVtIwj84T
r/kUFmddKL6pftPZgjDkLn7LeO4sH/6uwEs4/4dSGeqH0STyxwZzUroUr+URUmr+hmlPZaza8+1t
5MSdFfTReDUPl7AkkkVX1Vih3zJ8E6t6Wer9jDX/sSEhCkTNE5VxDUaL3QgWesugU8SfDgGKXzOT
L7IgHdllAdt5O+D5ZuurwoO4fPrJgDrWZb5rTx9T2U8ZVmtm/Qv8bvscFdLIEictGdINDXxj4443
7C1jgMZu94iu62Owfvp9uCMJX3fg9T/QybVhkpZssGP+aw9c+Ah7J6zN3+UhWj+PIYr3QBWzN88q
gARoZXlOtU8u8tDeYg61cHnome0iyO9en/qcEOiWZsldghgW4nqOKOCUgAlFK+V5b4M/9JJ3+iPk
zM03sgDFsC4GhkX8rT/P5pnd9XzFTJPTYwmnC4/se6ae0JriSaO+JI3vLxullQzN1aYttni/vBSw
FATpz9kSe/tiecU5xaTv+QIlUePpUIEigtXpWHWO9l4B0IWJ/a5H0AhKcgWW01xfrd0oPm0E7W4+
QOhGf0VbfyRziGLD8u9N5+S05hTm1tXJZpC1L8q2EtWmXQ9TKq/o5kgupiO1+lZJWCo9N/PDuvzG
s12U60C/U2ncZDF75MFYIvN57MfF418Xl9Ps7ZOPnQO4hFPeoNBx/Fx7eWk9kfPvYt5jWIaDRme1
F33f7TiuuryvnoieW+KZn3Fqxeq5ZL74DQpszupRPRjkrxkSI/KQijaekDKkNKcpJ/vXDjPkUPG7
DMwrsQ1NWVeMcCFzVrleGAV9aZdl65UBVhGowwNcQxJBTkQxcJrRVOXs1odM0oKUv1RgC9q+tG9E
vCFxcAvDY7kbCY/K81DKIDsoS0GLEyYJUmdSu3uKRh+/V+ssI5ohNSWe75pmOMRidMb2sPn/YeDT
lzFT02Lg3oVBhfNseY2atVsLwtOI9ZsakoiGYezFQdlVWAER4gzw149L5k2qI59Z3d1tMxc82Mzd
ehDYkg0mVtFNpI9h+UTmJK3QMcGcjhQxc3726ZAAlxNfQaSD6bcvfHhKsc/4aNcgxubYtH6dJ+Ys
Af+gcosc5eNFf3UkylypU7TFlXNgkXE53SRjssu7VrWu1eEE7R93EJ74Wgvd5TKCcQv/WI6Vv5O7
/PlRh/onwqXd78ZXmu9X8y1cliZLUnT+Vi2mHIO9vTTZkHZyCBr/58KnrKC4JI3CP+LlYx8tXCQx
25TuQhv6c4jnRwUzXTqg17U81A5I3mZxg4x+eQHXGXigCbSZcugjDZ8jsbCyxGiMMXYBa8D/564n
pq17v+88TU3n178/Nb4aq10yy406HZPUzcSmJYfTtw/mx0PtGpdffRaA+n7HjHrXOETRchBL5Xuw
/jYNggZ1cZMmkD6S0CjEY+hUn19y9EWiNUsVB9dbBG8W2yJ6Wkvk59TY+cfi9ZowI/4EG02XFNFE
PCWt6LnXOA8Kj7lnAVfxBXUsnisbN9jHkP4UkWL1gf3+BfKurcOVJYZIBcb+BczM7k2iQrJYzWi9
GB+xrnVgT1R1wT1/bo29n79gDIm0DYP9nhQdhEukNNTNb81iq0CPxxNvExwfDI3NMVS6K6zCOfJ2
5JS2VnbiV951W1L9EBiLgmEYJJ3JPS5U1AlME/oCRA9UDoCMBoY3a5J9aaxeitCbDRRJ9MTAhR1b
680+DTwwj2cCU1zCefilBB2GCM9KDeRSUltZDog4+llQCkIo9Ft7x8Eyli/vh5ZWURNNra8Z1UGO
Hh+GhPzyslD8hGu9/9zCy50aUKq19ma5ztiDlw2NoJv5XFm9ZG8OtiepBG/acHZZ+dAcp6CL338/
2D98VHqIcGWyyTstfZ3BkyOZEmKgoztjstevYu1RVtycaSKBC+EoUrEMeO8So7l7T9J4CN2YgtTc
O2ukeC2DeWVB28Zu/3u8T4pPxc8xllEiIuyxjIrxeMS4jEvSyRCWZwa0s+kBWG2kt+6rees87xrU
7Dds++Duighr3oA0q/DpScBUgCKPOMiI+le+/7WwBb+9C26+L9IG6k6IajhbECjK7R6idC4o8lkS
2II3Ozcgv/yNDNYsTpvq4oP7qY1e3AoqV5gOPcEq4mc7xZrsQpVjbUNMAiBKoa2DN6+IYfwclzj2
1J95j/HP0g76C+O8/v2nl7lM2yCXufbDGApULMY2P5Ofn7olrG+nSZrjKaymLzDQzIi1iQFhNJx7
hM1+F8icTsw3fhxpNSkI+9BzF7WtDL8r8qkbRkA5n221cbI3wh7m0cu93oUOh5MiF+yBTaFIzjXx
Gl0LIcVy8OqmFx/r6H3JicKtLhEs+3fmP6Lc7/aziVkib3FK1zlrn6bP9vzW/SE5DsoUfJI6cnxJ
7iuhnfxaS3+U0ecp6mkXGPJ1HHfWuCuNeh6pOKEduWvdO2JT/NIotxKDmvJEI+U4xpzm/0gHq0Ct
c3xx1VMumPSN+zoMSXDGx0lRg+bxSd+ABXW95kZIzr03ZXOzBY1R3ZqrIz5aCsGvqJ9Mk57WwM+I
KYiKBexvyRYMRag5ka/EDYT3rDjUy02Kzr5o+dCOVSI/ymx66QramtuJ/e4vpfS+nvzUY6PGxoCi
peNJeAaakxHHdv2XguYWWKayfsL0+HILgIyURm13lTTHSFrRPo1FT1uf6f5p5God17s9KXZ9kTyM
fKVR97u6jc4OIe1QWKZXxbOCjBlmgVNcro13Q8qRjcnSfvZj+Ikju3Az82q2UOcJLCe2rGM/6rLm
zFSyhQ782yzUUrkLtKDLpoE0W8E3aiz3OejooFLrM46WnspzHWKFeU4m0TaXAwY8vrM9QP/ZZp8C
cNBb9koXbhK6ZmDx6U07d5LzVm9OahLZUav+NYfAh3DBJbZz4vyhfyUZM+bhM+MltYuinydaEgyq
qBql3co42INQkeETxlq4/vFcAPRcxXcZRYOSGO5i/gLzP0YDExshM/Id5f8sqgJk1W31SWImkhJB
BaOEF+h4cSb9WWZY+xOrIzQFzstanXPcpfjSVvfUAXR4uS3O23d8LFTC48wwDm0HbdSqcogYkmur
x+6Zgk7PripHhefahSyEmsYvIzeHp+d4rWIUIpUKRRSDyxYsX6a4IJDA0OUrI4rMNV+OXcPO+UVr
3n+OW6+h/TGvzTRGfjUBu4JcMJd73Eng567q3HtCzmWb6Q7gCDLgRM2ev1Yrh4ltsIAmshoVhxEA
aj7uKUNLgWJnSzALAdsA9r0pgMlUZo95mP+cMZUPBZA6N1rQ7fwP95YUkMKTQJNX36V5oTYcNhxR
3UPgoecodkV/d7Zy2NHZRxOf5wtPN0XD33RpkUNUB9LVIaMUJ1243nskEzEl4L0wuwytVdy9e/3L
Wmu0/lcSA2xAOnEx2kMN0rzbtOQ3TEps6OOfgIzvIyvMUvXH214xnPsCBXba9rK+uitfIqnWiZuU
dmCn4nY81IygeMPIE8CZNfDNJ9WoQcUB+HYun3lt3Bm0/jlzLvwBJIvrald8+UCx710Zf56Nh1nO
gRiC2wb8Keti38oiI9Q0py3rKRH2GAaOW89dJdb6P4RIYciuZW8hGVuUm7fGvkvprM+Awk1NgcRg
WX0nlqiwffGYhzLmB8zaKYBc2DDpvT7dFSd0qGX59ntTcD7FB9gX8Akw34qRypMleSnJumTb6NHw
GswktUTngjzPt465Dfy7xgVbaLkrACVPMlaDfamZHzPXZK6kMYXtmJ5Ls4PsjsLlhQf9131Ub2+m
09CE+mUKih+c0u7PR2CE6gv0dP5cZBxpO2SWkD0NSptw9rMoXgBPoywDLmAOAieKVh0t5OQoXIWn
QtYsqLS44/J7llW4nbDOthHApSOKWkZXTsiPEMJ6ePFCNcrWQ2pHxH9fN2t6s3QPHWgaun3r13yB
aNzx/SP5kkFRIJW7DcSn+j5GOpyss48rOh3wWdgz7zOX/ljgaoNajWgSKbwl7wTHYeXV68pAVLWC
T8Tu+K0tu9ZqiNhpq5RUv+JypjwkXurbC18i2J0M1tK/xNqqGFQ5AToc6Z4bVj2SA8WghBvoJTCc
m2y2Jhwq7a+D48yUWnGU85sBy5MF5jdwuXZ1Kw6cRyXxt8PaRRoovP4w1kAJEfpPB+Ut1OkMHnRb
ehAsNkL1SvdUaK35A1ZjS9847lDfV9ceiyN88KkU0a6NntBq4nC8jBu5Mk+eaxjKdF2zTopB0IbU
iOOgd+lHa9PiA16IcBZ0G032zRkGg3/gps4tDoTTRiC4PGwPGMZLQcH1lap3/hIgpjBUsh2YWyyi
fy9wHLjK89ZlD7O8BAqLZEW31cCUovsLgni7wriFjcDxWXWlM5zx7NnGefl04lDYhOVUBexPy4N/
E2RTIyZcGmQGTZ/gVmG5CeGQ4PahOWFwrVbQbt4oglg61dR12ZWrEOKO6IYEwekNkhSFvSv0Pe2a
6edcX02pgfU/JTv0oy2DOhQ5edQaK4XxhqpYwD0/r9KCKDfD5MU3jgsf4XrX86dybmLoCYOJ9M0z
VKhFqenQ66HOVWyLyciybSEDVsMQi+BIibYGnRmZSXjLLpZGvsZ0jgUi+vsrm2q3/Si8uBMhhFc6
Fz+qsv/BYpk0mMRynVyD7LCIvqY8rqjJ1mpZqN8zpzHCcQoqljoyitUl+SGBnsl7B9/vhP7LebJ/
CnHMuQDOOB+Y+Ho0UdJPORDW3rN1ZWZ7ZGeGwd5OSzOrZuDwvLuDZ/5V3l9dZLhHG9uPSCJsh4lH
Gm8VfoedA6UfmnMV8AdWGM0/X9eLbRkxS5OTdfGJ8qz6da0RN2XJkWn9qGpJJnpBGXQ1cxOUK3Da
4I2JkaF1pT7apL6qYlehs5emWhjuf3cHq+s5BteIjH2bVkH5v/Qxb6UUB2yFiQ5uerOhrISy7asu
H3jsAxtRNUROfJaDawBw3GisMOjQ+10g6HAf+rrBG7OO/SnZlWHCJ2wuo4QjfReanq3v8kfwQlkU
jk2LhClirZ3RIRs2ni01kQG3KUaqFG0zMWZqVNvvxjygDRuiyEvSj55RvZsq+tMvfG5Y67F3wBBY
HcFrYXq5jZxqWgTiHlyfLPq53AfxR7XSaNm7/CHbAyCm9h6Wna0X+UjrZPWBFkJHvJPZ5T5YxfC+
4pwRKHg+Yel/v6/vJz8e9VY73tbVHL2VLOVN4/vtqX1FcpgBDus6hR8EW7hrkTq/IkeJl38p+JK5
XWrdOcomw3oCSxf63RN/qGsS4RrgLSfuSw4LbD7JbVB/3WhEAHoyNX8rpgQaGE1YvpRaypSnhmQF
Px2VYFDI/Fwnq98kgZNRUXmlWLWh6ezS3dkG2IISAzvOJllwqxe1VHD+ThoBUEx0bqWfB07el1Xo
RbSXB7oDoNGlZNKPcKxHW8V9+0Na/JZe2gqbTlFZ4Cj2dKpN52zazVFnJkY+6nmOoBMSBvBNJWba
mv9zwVdUTf4we+45lpEmqZN43TlO4a6AQR4jdKfTP5DRyskYBSIL5d48gMsphUYRSQC3hx0CUefp
+iIcpX0xwFGlEkYeMiQ5GPz8hR13GUrEEdEg3/xs2djjqwPQHa6+PzL+PwyNqq9CPFLVoq39sbPy
kXF6uFF9MvZUER1g4XWvxJ2ay/R1vNo9nwdDw6hfA16tJ0KdhQpH4JVWABmg9UiXeeRUCIf0rH+r
Rzfx0WP7vfhFH4UqGe2UAPyPBlBcSr8/cUGCKrsHjJfdlYG12r/khEZSOHMOa/ZJV5NZoYz+hgvn
cW0hXMjmPlbudqOeQR7texVB+MC7ERgNtkualvZ7VznvDVzFUF/3/cH28FwCyyTUNwjlbyfmhKiK
iECZipJH4MKAV6KM96Ut+eVeYHKW283pWX9Q1wQMgOKBpnfYo8jEe9ufsQE5Rf1ex0Q+Er18u9xc
3lx5f3QeTBcTGdWew/JsllCSdVFd8mGMyOfhOTJEG6Btck2m+F0d6gErOr126INroPt1PeDV3WJF
JuEKNKR0OticRkU0FTJMGtQ/6NewVhNcC4lWWVFWm5BQ0pngC0meJSHVaCUJnEu/aeVYxHynGzdw
n8nZpx7ex8GB+bvmOMIz6eidUHkd52NJvqJuO1/NwBZaTQfmIfLE/uNV5gE2s38iC11Tdf29XkxW
h7AWOQ2qzKXQexFK7SwOao8OvXwmjKgnMP6TnLwfSQMB+1GvuTZPt7e12Xrk6hSeGkoPYcegbFTo
EMMhnggsrNshzb3tXMpR+rKM3C7L6k6WOXd+nR2WAJqVMffGHTnUXF6uqgVmGCHyeJU6uVtnuHmx
DEnw+2BePc2uVatgZ26cDVVO6JaJf2LmZQteyWJ8U0PYWey8Zwi2dRlOWeV9fDTM2hd6Y1oRVTah
KXc5w9yn1hwSLKpeuMwzdI4i3xZ/t6lZshGrTp79AJHHugWVXs1H5Fdjc1PLylG9FOHhlJM284mc
zK9C+sUCiuG4aouzZBD2tLCmb2neTKjYSZEFeEOfxQcUKJsndJ7U+l+GLtJhtH2Q9gYw7paxupH2
KHC6J7iMmstDil1BNRkWgpeONpI3FpQt3LGw1aApe0CFpRMqwDZWneye3M+s7VefV36Q0dT+3GJq
2kbZ+OlR1bHUuHS0NGnJuiGE3j5lKJTWTY1uyw9uZeDeAt6kQNPdzKuTuSKFjO9PvPyoGTSL4LO4
PuJ944PxqllPATjf4ShWVpa+tNGHmfDQU0VxzQ5+X0wNKOkszcrqynu0LBKHVIeF/stdmzwB+v3X
F7qa00opZhj0Ms2VuRl6vsiRN/5MmXFmBhaR9wDCgb8jiiBDKlN3biYxmZIHHH7ez7Za6J2NQUoP
H1J/BgBZc2dk+qv+n/fpocCfeiQNxt5HdfMIEht77GOfMfs9hUhkDxRGQtaFhy0zMDgP4gAafADK
fPByRske6t/d/jhh/q3wQfgln80mtEyfQJGdkgRpdCcDkxctXpaO01VGFuLi1bTsZyhf7D7U/hG0
6da8VgSxK1kWsPfCQ5NvoOi/3Y9JM501I5IOtFNZ64LTkehqQims4iJQWmml/PtupT5EL/pXPMiV
ZTAmdQFAXSHzUBLPNGtKn3ij9iy0Y4lLlziO9UU0H7mNsVnPUxddnlz7E3oBOc2XJsy9JUJAO5Ti
sUPweuryse1I8zl1+QKxTzv5MRPc4CblRHhahs0hJT8EU7BzQUgphw07YHnKzrmouZ/7lAfhEqnu
96UqUMZCPb3Sy8v37+t/X76RXUCNH/kuU+KKzweWim8bLXDR/zCqZUzQtyPYdSO+/SW6Y0bp+OfU
C5r5b9sVmUsp6KfOM8U55dAsCKgIUCv8MoJjM6LXaEhbICArrzJ8WHgrbIsiuvydmtTGxSyB/QLn
np1V9pXjSVIvd2mqdMp/FiJUiMFLxcvl6sOsYnff33MvS4Vl/vKvGdGiA+lI2WI4MP32DiD3fFt6
z3rzUORPHnBdsdgg6zZDhmZeL/T2VXdyR85OkxIzoSkvu+LQnMn8SErjrpUnYirYeMpK3f5Ow8TZ
EUnS2mUGJ9DLEwbxpsSjpV+Y85Eh8R2DRRKUsYTAyoTKz0g6uPzX1c/LPEIIgWEGaI+rYqDfktMa
92j+tkvYZqcYL9P5JorLpwf3bchnR4AXwugm9i27m5vz3eu0FNjVKfWPx52o4l8rcZV6rXnqYepu
f0QCFYIIDQTJsVNTHHv65P1bMVrulF9rvvCazj1EjqrY1htN4invYfUORnaMfybs1zC7Z6om7oTp
I9Qegou7tjIt2gxQhilIl4k7dvQUbF2RLWCiRzGf+APzKj6HfWDrTqkiPearHkYGTtqA+7S8Rsf+
FCHmcFyH3e7z0BWvYOlReNyp1EGoLOc4d0X8LMpPioCb2uTq80jkrxob2oAT9NqZZvenuaY6aUxs
WAxFjbLuwnGlGBKTkPvr4HyMMfbdg/jXwsV3PrupRdEJN/aG1zzzikhPoHqymyKS8L4nhdugChVR
Qt5fz3FtRBmHUx2xT5FzDAsV7q0F5Byr/oyoHrOvWYEkvK5KkahgXzHVn6QQuHvKuhuUP4wTM+7W
sdLigFRC0LIsrRgZxW58B1DkRVnOA/9SYr/HSbb5BIVezXLbX140ad1deeQhZ8intUoLK4AnQ9Ue
XQs4yvILIeqcpWK22O7v1EGQFPaEzfJ+dPgsBibd6ybZSzn+KgILvm7t6xIcLSTCal0UIG86P6Mu
V2LmgiaAf6wXT5AAQCnAa91U+M1A1g6dBHqMA0XKJJIdlgNaGWUhllMEyAqxfFBbndtWTj10r2n4
o9QCJq0OcegZt0K958HRsQXvIKanIWUflglhV9ZA6yr08Xu6mFokZpspWeOsf4x3dIcL8MuuB5Je
KBLfbGXKBQUZO21GekyJwxr9O8CczBkVU5/lu/uo1ZVPfGRELT+jcsLQp9CEr3gfbRDvANZOadHp
ZsYWO5IZT6JR460+ymxP0nVjnKIVXhlr3FvYqtCIsd/CkoO3jJxm3z6ZKc/iwzfHBVHWXAjPZmJH
1L9fIPQZKKrUXduV2IlkmIPcEF6XxnTrg7LLZOjuLO9hMptfr4urocsUXlePpcfY/J+lFDoTG+z2
PL7JNgyFqFyKEPbsv9bnsUbHu/3O/enEQ6uVr0fcGX5wKMfQng5CoS2RgIsfFGG/DsdY5S0bd6j7
T4d07m8nU0+jAgm5CdURJkbHc1ah25r7FyYBGzAHyfOVl6yhux1kLFYWVoJpB38xVyC7xbEtRdCA
iNemuli6B2g5FukTsfKKLRjnoSMN1w5QyhKCygVh7DVtq6d8xb+n8Ei1JcamDlVNr4SwEGnkMOBm
ZjzyhR6GfyoRGS8KFAAC059LQWrQ9ensLWuE0Er/CAXY4nKjraUrxYFW5/xctQZfEMNctv8c0EN7
JcSiwo3AFaN/l8WDbZTRYHfKPJxiBkj5lUfzlrt34ehY3imUk0U/blqCO8LfHCXBfGfoN/x3IYXp
Yl/eNP9NAOTCn+7QEq7CoBSbweHkVuNttrkMGZSGTMW9rxAFDKAA6gOd1ap3tiDMHqlQ2hmDTyLm
9iOjRWG5JWyWpCVzGj057hr18X9wLBKDMpW105MdBxcQ82ySqsjXa8+r7/6AZLiM7AqRIDLwBQWy
LjloU5Fbw9U8oDv++0mKJX3pyqppsAaPX9Wl6tkAqvJSJ0bJX93oW0EpQozSiiYWBvmz5r2zQNTd
Il6/7vNpJTGpsOYm4sknTImXgnyi89j7VCh2vC0uG0Q852xhiLK0IjUFqZsh/NqLNhwcGdG225Kw
Da2sVcPq+ZXGEpn/rhGAd4buYTmOayKTCWo/vlJBlIyfRh64rsdatLVIx9FmWmQe2O6YHPprsUSF
MKFstP7cFgKY5J+V4n/WW0Hy4S2VnxCvqQVeRexuH3OrnV7FZnbSRzL/6+YjyFGDTIXuhfZQsY92
9cglOAh3eKnQpDuz45dr7Lg04CJ0CoRaaGYeSb60TFQzD9a5Ma7c7SrxmCtWaw1vy2j/YJtbNCbi
Y22wWPhGdbe4/O5FGNg7/Qtd//PDfTatD7o0jwOY+Aw8Ga4q9I1u2T++N2UXYRPBQ35g6kRhxJ9D
v1EsHtY4y7MJyi7yeLJi85DNiZWmEQlY8jNJevMnD12RpknNSjBVdwlh3mjeWIbn8nEM1wZgvXsw
VZzAG5EypgHmAcn1e5cLa+76ew5PJnih3VeKIizR596A7FN1xmaRHYtfkAv42eldXpP/gTbGoII1
8ozX8pDD28S/kJ4++b9/aFZjS2Ysp9/rdXj3Pn2wOb2+62oyjGJz1Wm1yLR6cGYTSHLus9995tmY
MNVUlOoU3vhjLE9gBNuKn021zUCBxIfmvT3Sk+GYNRJ/JuVcMVgc6/07wO+beaXD8+uiFoSdmkgp
F2K3CDc7OWbgcxYbnGMLvo97HBD56/4n8xrifvtuMJH24oTq6Ldsv7Hehak0CmZdhcaUnAhRy4gR
Eiecj6dGB6m2qiY1kbOYOBfDOdVktIommevatCcCQsVePO98QftLlUnpGoPWWo699Wqut6tuadK9
p19yG/Zn/xnrm6VaJq6Lmf81d01cYgp7GG7HTgWxeS+HTBJxpmU/A6BlW4g+W8ub6wBlR1H7FL6s
CHezAYs7jxkQWxhvj0MfHlVeSlJ3GnKWlkciV8GaKIyV59HoLIBMt3lrK3as5xBL3yaSp4Mezbpb
e9FypzTy2cmP002JiXGaGDtpeG21QJBc6ll1cJ4/RUE0RmQJdZ4TyvX9+hKHOuGU5flqtqVzxRvG
nMEBb76oOYDdp0hASpxRoEGLsFb2qSS4oaUgeuLyl0i8yVWL6sd7Q4zonnILrSfEVLbwGAXOZkZA
gXdpi9F60YcSw2I8B5M3NsKAYWefixv4Ux+ksISR23hboKeFdRupj/FCKegp21epNRTzYzd2CbOJ
++702pq3S7i95+HIq06YAV6aKBGcTZ/9hg5jcSGe941Xu/n8IuCSU4YyZpE7r8V1/k/1ngXGpD0k
wnSs+jHjNeNG1MMPbLFbInMBHCxe4fqvK6vGob4gcrTjOObu1Da8W+pSiGstr+U1x30PBxhUJNMy
RQEIgi/miISAEh0Ag/EGvPgs6k065eCWT2LFdma8yapS0S/kfOsZqu0U97Irs2UAYiQDzocO4CdD
XQrg0DXcO7cQVSOs/oeu65y1LyPue9SK3fLnDsay21gzjqEEn6uMWrB5Y+Iss5aNReClM8w0BrBU
V53xXuo1GIukv8hhCtSpYOVDjhNIBdyHDP8XOv4zPGz2tCoISGuTW3p5gBOVCPOZ/qE8BbYQeh/4
mGtFMzKi/M+QNdDI5zIw6BM4n8811h5uy/ZPQ1DumQtC6aMhA/ySBJVmHBLOnW6nc3LLk8Ed68lq
9/nbAtoKBHAgZYIIUmYhzt7JoEjbkg6/YE4xGzIHezD4PNA+3AS+Mm2PE6eAb6r5l4dmqncNUpxP
/H6lNeX3xfND4ZvRrkGZZQBAsw9fGB0MQ+n5bvIhYb+4WnzfLTnPczpSekTPwm+QQTq2j3LK0uK/
ejFw903iAO5s7ihCBds0OU1JSmFBEz9Lraz/RxNtZ8v1mhF4PhQHyErwOpNSM8THZ1N7x06C6pS7
T4dnPa+s7PIjILF+aD0AvFBNVXjXByZfInfpAkFh5NwWvF+67OYJRR4bavNXVQ/0U+2MnyNeJVwA
wQhznGgBtr4wY9fGX9fV8VSiyou1iNXTOBRoTrGTPQA5WTFM9ivQKjfexxyG1KHAHkCrkiGwJfeo
7fdhr2SMol7v5+ChEyY6W/JmM2txoqSjPRojqneZw7eu0NQMhhC+SMI18B5469ydBEfXJ5XEb5Tx
qY83iYOoa21k5SVLCz8q65k/prUnzHSKFQBaAxHvamkuJPd2DiHvh4nvsCFrQcBY9wVh4sSL1aCo
FgXr0UI46NXwvyJsklLrRguv42BBgp0c4VxZpNtMPs644Y8hvWCNW1u+kz3n1ILXTchT8wJ840he
eskwAQUHSx333w2g/b/zg707xRd9wrkMPJooJs5AgUDKyz6zu4Oy1gd4XVBWbmpqOMdh8rFTEg46
wmY/5wDi2zuw9mOwZsRzDhwDPhSPbqFj6cZqYS1F2rZ/TcR+cJniPqCYyvbRil33WArI+eND9Cft
fD3ioTD54Gmk6O9DMT2TkENS3DCmkDfCKNNljOJPCTvIAoMozO+Rpz8JMuP2z6tQm6UM9TDN/ZlX
tHNUit7udyMarXz8HLeSgeiIv+pRC2JEQQNJv423fe41fP5E2Q2wpnq+/nW6Fk6AbkmI+mHJJAN2
ggu1iCWHe+XW3KrE5saI0x7kkZ/0EpozOVvklaRkJi3KaryABl+RCwy+mv/hayFXeUvQeQ6Ihruo
ksh+Vcop2kZfk7fJizlr5R4s9Y10KuAL2xrpTUtWEka0yyWU3ue80FTuD8ooius1pGCkkWSLvRyy
UUU8CYc/hQFc5UGv5Z6uIxhvr0kHLI9ooFfEhBz6fU3iJwu9YTGa6e5fFvBUl0FAiMeNT6dGHwOD
0YtBzDo+gzI7Hw0717+OS/aQ+OokttDouapmpDQFVVttzIvGCW2EX49ihnCo7SU/2Dz7qf4CPjqz
Iu9HCc6ROqH9Y6EX40Zzxy9uTDpkquXBYocvDRwVmLoHCsj323QbwE73YcqTNFDrrJTW9ej9BEe1
jUJtVt8xEL0CxaCF/T/wHKmGrfHUvzC3K5HTXn/BThNGX0sOpXl/kIFbRTr0oIS4t9dS/3jPcJbx
xzDmwomO4tZ6M1uEwsZnoQBHnJiTQtQMs8nUyXu6MoLOrae721gqWdehUPOENDNpLc/5qI6I3GkX
LIu5eyF+gvR/AIOlr0nD8HaosujpuPF01nEzM4hTPFXy3lsr6V9g+35Q/GLsdWo+apA4khB+M6MF
9u7tmPaCz8ySaIszvAhykio943nikkwxIxerALKCNln9SND4zjPyOdNPE9DQ6VjqutqlvRrDGNy0
xf0u+2McwnCNWIU5gjXlOi62zskxG2LZOfdRL65N5b1OEAZVDSfAst6X5sFsF/t8SL7M+xagPRJ3
OcNhfHMURHn3Y7YAP3q8zlqNVoYRl3GJHHrx9/8J0p+9AYnF5TjAdMPDzvRJm5CeTtycJaz035UQ
WRldhsuFtqhYTvnDwNts/NNreRh3p0UxlmZ077+DQrQ3VezcVShN9lO/LupCsKDe8N21d6A0yxSB
Up7+OrLKQSIdH1j7fwaMcsOlHh+sUVnO1MGzhBIaFuZ0s0n17Mw/zvmzHqIUqzUhnSzAu0NTLeGj
9oyVcomJEStYiWjXRReRgWeAhk+qhFskAF/HkHio2G9ryCu/0RXFTNUH2yHxZCqCd/ubefw8RPDP
ROQpPouyb28i87ltm9mhjaex6y/BNHWIZJWff+cdeg+g6BhijAIMO+3OAt+/AEhaDTdshb7ldgTG
+QwVb+qIiTgy8J544BJCIFGdngPRNplaIc3IkFNKG//j+htxCGEw6CoyfGyVO7cD8l2wZddUgVu/
cavCQcMEAWoGn6d0AgbcNxWZC+JWgUyO1+lRDEMRzXdT3MssOe4hSIQvnZ89DXjmN1AiE0dzDewb
XT0wH7l4NoKLI8m+9PjYHliBIuIZgl5Jsdco/VhKNEoK9JUiPXBTIpnscSY3OaIAjW2xJjUaDzT5
B+0pRc41nDkiS57awPhdJ/wrtwbXtw1DkGWLbf2IaaGqVhmxAmtE/tbkq33N27IhiSnTutpqPS+2
wVqAnszq8nNeJTftiHNKPxmkep8ks9n5Alysww1RgFRLTQSyJH/mccGz39g8ahQKQxZsgWcliEkt
NzGGohMrSUazOaL4EEeAQFA2EzpxSE4ZAYEpFUedBe9N0GU4DptoQLny8OFismlBSn5KZhpwHYwG
nb6d2ZsW6iBf/eXojBrZu1wDoM/YanCELskNwpBBaapSuMBK/mO5wZxhnG5anGpfT7IutpjBuJ5M
8aCjogIb1YsGHZhRDxH/+TYnJAnlHFZo4NtipjfXreGf7JsSrRddDliDstDTJlpSvcKoMmMRB2j4
vW6O5TAExKsfq3b1BCL6V50Fixt1X6LUvQeAjgyI8/XDxkXexpJLW+fPLnAhRWqG3kXQzyXRBIXB
7297av8b/3CcJfG4uRalynn+03k+lfHLQ9S3R66HPGeSKFIxv7sugn0hIlQu4J82hhX1X4dm6rTP
jZIeqVjZmVvJdc61CE3fl52hpK4GR5KNvhTd8NJu2kQLusAhrmspYR6+KxQv8LKVAhIa3hLLbr6P
/K5yx/wLJOj9IiFpnqPa+t1j7TJ4jU/Fmc+MpM9wgh0Dmt0ocPsRkZt0uIpxkigyJR7sPS2oR/Ao
0YGSYGEe2DMhcb/kZduYBodjw3GzjekEhUfaf0gQVg8lBQzVlDEZXlpJUgxwltJKL0+qxXpZcpn/
TcC18mxHBEkfN5L+5aj0jGd8Be7q86mccplx6L9xzoRi3wilxYfM+bfheeQ5UPPoeoDT3doVZ8Bd
7C4LXMXyVmAeLbJKbkCWhLtz1k9GCsHj9EiC7Urnl4NI+TrTegxhKm7cRPP7Ons8DznK9zB35fDs
I1uJUNIfo/XPCp1ypi4mUEv9gdWWkAZRYmYo3FwpvR3YW+68dlwPJoxm0i3TX5wUDvqhAIxt02yQ
7kwHoOKbxDqZVhIV/VwqWiVXM+wuNBJJoi4VjcJNIDGwaJdrqxmkRi0Y3LbcWTvZDs+Ea1xVvxaP
IFSZ3yyza1LcYy2ikXZ/VFiJU2khlU0Gjk4Wg6/yLgJXV5y6Yaw4207LB8cSGZo1wNBiPWHKRoug
y8qfo24zOlUgXxkH3pJx9v30GSfYuxah5lWsI1E1kOJ6KaZhc3HbM2MiOsrqS7Vy8hkXlgX7Tb3A
bfiJdF8loXUc4JEgvNsXLUu8MaUzH4E/VMQ9OBZsvgVieVA71tIloRtk7LoYKzv7Cs60OwcmQJCe
ugSuOTnNHYsAeo6tsXU8L0S61sMyTg6kry+eeQ+UGN9/aNt0C958+MFfWjJAdjT0pWHAMPYvHRBE
RvA7wt44FfDW2U/D7w2SVXWjs39C3x7uaW6JkAM734uYdNx8L94o7RwTMjYqHehKghy9EIKbwemg
JC/UsOPO3PbmSwLjkIfYrDrqDZlv3own5JOgMkk3cgD1XtqtO9nvwIA5YkQPdZaYrNGqgszO5ZcV
0dl3OzzMY0zsL/0goZrfuKBWSe1NoH6nblyzcnYjVJ/SEjYfTz5dRSLU9rwoIrSxkYN/UCASjUEn
y/szaVLa0RrfPTzxc+pV5hgHUlT64ghQYcfTFm9mUVwZ2s/k3NGhdkbigzvQA+qQsir4QIxn/3tl
Z1OjWCI3FSEq7/1Qe1F5U+W+kA7I8SXN7kdMH6I/4bGO2OJxYxIe/dFxfusu2Z7E2kZ5YoqFr/gT
w+yjou9peonci9WwBPMMyrfNMg83kYcKAGbaPMydXfSDTMLJHC0TTcf9gQ2mkKiIgUAt40NPzBO9
oPmTGKWuVwUNpGlWJ0XOcQVzmdT3QHps79S8K2MRH8TxmIGAawXC4hkRsIF1IwVhiIPDiE0UnmDF
iaZ1/ZdiCKgR7XZW07W+IJzqwsUGCbPob3A09hb5zSx82+SMMzlaeAKTxC4nmgDwFxWaHBE5x/UJ
SgLnvS+VelQ4LyJtAixua38rBEljAn566KixPh80Vw+FYx7iliIUy9MeLWteOb3Wm4NgDsH/anXN
/j/i7e4KE+wV6BGnOL2Fjx1XnrNQdkQFw8PzAtRLdupt/qTfUFhCC2SZcb934XGx8nTezhVUIkfq
xJpxckd4ceQda/lEsPyGymb7EcqoqJcS3py6r/mCTTzvwN5XVSYu4kJQdmbS3VkPMigiP56DAr7L
6laNfJakZ8TWNXWRpoE0YYv1raps/yAgp+25RAeMgxMz0aj/NrMXVjkXzogPeoGVwCo+RtLcZBLj
BAWII4RKRzlFP+BvbvOZYds+TNYiz8T9hmMFW/WTXTRKBcrn03+it4uzAxkr8AyuV4ZHG0+lwmMa
Oy+JTqbxTtH7hbKqWaiedyNl3nRBPMEp7a0L+6uH7xjGdJd/mTaJ1nPEDkB1i0GBQACspMcgZgoz
Cis/HIkW9x0jHqUNkKai4XJFCk1Zp2/rlLVBs1zWoEIeVkfOTJQ/Tv03Azl27AEZO0oYCbxYfPx6
/E6X8+ChLB0rT3TWFks1DnNaILKPM50uRwIfF7ZYbKKebq8ulAW71XCLASIcunb56mvD5r77ME9G
My46Oh6IYpvc0k54zLjAFKRZwK/b82zLHMT8dJbFJKde9TRHtbTUAPqI6QltV8Zq9OAEP/ZD4UzK
8wjlsSTOwa560eYCOio8rpP/dBN/nbRxojGbglhNjP4MbUhlps0ZAtR4GfOHKFhT1zQh56jF/bjb
+dgiTAarY2orPV7bNVpMxPgBxtMk2kyQsx3c31ek0UGlra6u93TfveW2Ag2LH2mc9KY5lE2INYSv
1M2lRgIwg0ABbXe/OyF2oqAiWDcy4wwFFuJThnMfwDCAFAo5sqeKdwLANsgM+x2DDAjrlGU6S9yL
d0o7qESoA6sjHg5ocOmnLW0tCHJpFkI11cNLJhXcWyWbZYLNzc5N/tnppMO2KtWxtOkDLOSACyDA
EdVIU8lkPJ5YsNyTE8fzoURHAHmUa6IdWaChu+aEmJvyQlu9tusWfK1j5GD7dizSOZxrzwG8TBhy
ImrYnbrohOq8sovaWzspfiQmS4M7cszGVnoWVYBriuRbeneBGo0PZvlglHOP9rahA22oe08gc2Sc
SjQHpHMQ3HcZntOmpSimT2Y5ygFqf5QWHALXkYjzYKrpy4f2bxcHIAZSxcZoX3ZPxsCiBmTYbxuK
BW+u7TLCWphgiia+T0WpHioeHwKmFcYI+q/QbKQ2P1kvP0Mk3Jje4Vj36D1Lkx/7d5XdM8msQwtP
YV5TvHVt5pcCDJisJPRl2XMOQjAPxksM4+OIEe+ZmVbDLiSIKlTWnCsnjgCLcZGfev532VgsEusC
Xp2sEuMN/Oc8+cENoMqDwUU/ynDfxO5zwDvcVJWrhVAfFt94LdvPcwR1WvukzWtylTckcq5ARo2u
nHZtQIptIqzlbnWAq9cZ5zMs0zdPFCaLL3mcowqrqyi4nBwpPDlwK1X5hJ/fp+vchztV/jSVjIk7
IjC/Mil+Q0PLpjWHKln+XikNCWMeC9BRbRBilKTEso6zDaZ9JyA/LdTiIq2bNozUvNiK3UnvI/7B
JazGmixwZg6d9nIQEqpKKHWjvUm1xwekS0OdjrXtmbrzpkFLk0/v4F+GG012ktRGkQ0X475RMscM
7Z9ex0t8GsbzYLzDSMUDxKxecX6K/Rtwaew+B7NG0uyOS60fvhzN2WUHettUO5/sAbVcOqXu1CU+
OJs9X1cQ7RsgfwFN8qOH+PgQ/PJ7RpgxW9K7CmRrpOEEHZc8cFIoavvrM1S7ID+crA7O0lFNazn8
2gK8MuxEBXat41eIYrXgRnmJeQNd6svKWT7/DNjlA5rVd6hedlYvglKdYguy2v5eZUDWIHoaB+k+
YK3/aKnJYQ+Z3p27548zWY1MNBqqhw+VisOEugWnay8RfX3XCDC4h/8Rxxc33dpz/RZDbTpVojBo
OcByQySQR1LjfMMUOvwlozPpTKsIfzd8fnm1qLG3EDtIBtvWFJvRrMiCrWQN0h/TEoVkipZDu9za
PrfryACibjKO8WWDEnBMAN21H33ZVoPkynVGbLCFoqATrDp8CrWvPApyFzM8shQNW15H3C96aZmr
wk0orCSBVA4cDe6OaWZjMx3tg5xFvIBRUV9JquxvZri+fI3S3h7iZsQUbyys//4eGXCM8ReImv33
jhV8xTXoignVoRVePrQ5X510BjJvlvbrvdnsi13Ckvl8LlyVdb0Sfm84MMnNy9cYLsylM1Kx12i8
2FnU+V7jljN1O8PtrPKOC5xx3+o/1acOO6pfGAnljwY0mp3tG0HFsyhUtxSScT3ZiL9N9NoST/Pi
ZhUs0t1FgQpBbUx5PAlnz9yvU7r8LrjFLLcTscdToPS5cvQ6Wo08mn79ax6Z/zKuRKwzbgcVciDk
3UNY1B3v2nTXhX7ljKi6hX/NLqVZLqXzGDsI3VNji7sd3ZLfc3scHZ/tHurvypRhQ3co2Lwc2RJu
wbPuLYkSPpC8B42E3alv/COCDXrOyaPY76oyaAiZ50RhxNpbzXIfG1dN2BYrmZ+XWHDgzZnjvZCj
aXHIYPRBJBkUamwtHgBpKSdNB7WcmPilN4OtR7QnwYq9RmKOMuJdnjAeBZKHDYcRoVcNhnD15IJ4
pweo0igZcG+F3MU9eSqMTKlE5I6a6xw12Ixm6wBKGhvV73uQUvOD1wmh44/3uQmqjSGMmFy6D69J
tQyw/xwi7c20E1In0sF2/rt4oJYX5P4T1cweEM4PcYTrcVmxBcKhCQ+falYXrRLz6w0TL9L+34AB
+HspXtAK/1Qc6Qko74io7YL/+T/9KzErD3YGeGFaNhsSkaLKYEGhEn5PU1u4lAnMTv1oWSt37P2d
1gusf9LOfYz5XR5KsR2ZRpT/HrxuVKr6HQSKSf2SA33XD34VsNq33mqtPAuGgaYvxOS8GsDJUWCg
LmZjOXm25GtyC5q5lfuBLjoO6gb95D4v5YYx6BfDFLlWc6wXmD6xYgH8aV00wjAGDlJtVpQcOYqF
6dUz0K8Zl4/NHyhJse40NEn98K9Rmr4IbAkmjKWRoSZpYPc+sYg1pibbxgPfmW2bFK2JcEJGnM5i
9ZSDfMyO9LOGUqSc45AMPwqNBXF16fifaoD9m+i+YHfUHFu3bsyE4zMScjmcEkhsSTSKVbg+lyR2
xRsaAUq5jMoE6Ws+uDF1rPOECYeAgV1RmYfJOFRNagGwq2bl1dcrWQOwXw8yEg6W5qPqMTSKEkVY
glYoe44kYpihu4tUW22aV+3DswzIYB48DLfj5/JYUG05lz5lCpwtjHu4q91X7StQwI8zE3jiNoBx
I5fz2uJsGhlKC6aB4USgVwEMnLq00EKzThgvo8cLyrD2w0Vy3gtfOmD3cMJ7vTzmYt9t25qqsdBK
0kV3Zfp6J5wyNDdmES9yCEeUvSNUZJ/JI/wZ4940zMAZt+/bMpZJP1FsDF8Tjt4mpxJfnzXlFQIY
wzuokRueoGMLclxhNsGdysnCWTUB4yDikvIf8CsW0VU7PYDroPG99tQ95XWSDzUDeKu9yITTbJd3
ZMzBRGRk4xm6+y6JqgfiwxiyDWHGB4AKrZ/gKd73BINsgLpQWnIb7la6+WZevyJtYg+uyl9Drkyg
/BQtNSDXrBdcYGwkOIx8wPK55RHkXx2D36AF7L2k0w8pMMuvo9En3j2IfWQlLMq8VIAoi1SSvuPO
JquxLMmfMYHXMrMbCtW1DUtfQcUYyJq26CLTSh5FJ0mHogLZaTvDRyzpAvmCsF2LvU6kYLojC7XO
OcuBvL3wv1QxnTiH8xs8D/cV2AQfqr35mw+mNl1uoq2cUW79G3aw94GQpdORhc1KYccfxgAHnYKa
05p5ITILGE32x/0vA+T5Juhn6t9kutS8Du4WmelzTKdSWkM0v5c4qkDiaCvmigRFL/2TnwkM2e1L
xq3RDgq2KwA/eNHlhXcS9WPjrsZcFel099UwLh5IX+S4hxXLHzXAK7DS6Owm3wNFmQRbvgTpqmrT
HRdBeDvOx3F1pj11KYVA8/S8Oka9RGfFXUiW90oBT6DqK49V5Ppicw4bZmeP6k/OUqbXMHIgormc
4godzMrXdyTgih+uOhwo3fxMTIFcpTKNqKG+8//BdUTUthB+N998OQqVYUAQ5turw3kh7hQpcYdZ
6nKHboEtY/vEfhtLQRNOoduSOmqzaSjw7MvuvVe0cI4DPX4h1VNqploQu0EVlDCF2EnsWxTHSk4M
LL5NagyRiRMq3Lrg/uP4B00dhOsgIahLLFUPaHPFsp5mJsUDh7+2ii+jjLF4pxFoSdkHbPblss0D
hvpWZ5WHJle1/XPXdFod9KjZ1yuiM6iFz3uFlBfUFxUOSlibvjAjnQyWOaNWGMbbvas/+IOha4ea
XgSCMscUirkHSYZt8kMYZ+0zDqRzDQaBw+FZPvvaSPZMT1JjNu2D1HW75vNAp6bHDuYxEIW07Yol
kRkjrp7wZQOJ5Y29yExi5wcz8GCiIcftJmhcs5tv1nky0ppapYvP+U0r6dKzWe3Ph0EsREyWLRD/
QxjlmmssDsZP36ZRLmSwiI2M15qwpcX3TJ/bMYG+9pNK0JubRA3llV/aQRIkLRjVbu/eybSg438d
cvh/hAEgfRoE7bmgpVvSvXqgV/21xOa6m4GPQJ8lWB2VOrXjUNsJKrlTooo30B7WYTYteEXU0/yW
Zh3diQbUxALmALqnBzErukj1tRFoVFVt9UAKPLU9VTwjQwWMFka0T3FjKf/3JP/FEdJHKCv90GyK
ht+pkeJ0EZa2F4P1lLzFinMXp8HzSWXQAy/u8jnmSItvu8qJiQirbFL5PDObs+2EQ9QBpOUOQ1Rh
qDJV4xEBttpuV8RiZhuUZLWxwiERcvHE+xUmDLAUKaYDqU8oIvAd0WqUGKHUfmVCUzviuOGNHoVa
LyOb2UDzd8ZzQsC9hw+tAaFI4UqE5xjvSsrz7JxTxdxAl+K6PXi82m2qTIg0brGYeFF9Lu/pLyKB
dJA6Xix3S7S7RLCyWUp/+As7T+2fe36p7q1Rx4cHD4A4/gd3pKmnZJevPVjE5F/DSS1Nr7sj4mgj
JVqkKUfjUkQY3Hpvb1hbVQ+6OdUibxRB6rYF5wO0jLe0OZwoe5F3oiU3U8uredQ6Fggl414yUSEM
VXr98IGJgS05lHj26iikhHq59mgOhB6cTayhk4SpvT8iT4/DOtJCfOu95XYczOQM0PtfKzaDS3WZ
kw5GypHZ50of3KsjY6WCTu7DSDz4vhKc6wahpUVOsvNlO7Sq0khtx13qGHL4z3Y1FmXdyFRNMugO
c9BrAEUxMVgSM0zYawMb+aeqELAjC768t20qUf8GL29RjMCZuUh8YaCzAEn+vxKeeY+jT1IJ26BL
C4iZj6iV6NFP2l5ym1S4tZpOTckXCdBUIHzEweLC7RvlqHTrHua6uBt15R27yZnZkqo9e5/HfBY+
06Xa+i6BJrWad2/9qxalPdhaXx1S4kiFHqpJ+eLsE1io7143TXLRhLRKmDRvH2bqQJ/OO7Ouiiwn
TAJYBNJxMJki5djtNWY1NK6d9wDFxl6l8OEMERRsO30hxEABKuK9916+EM5trBzvrEyY2JG9+T1A
EM2WGB4Z2nf1+2MVZkkb/4Q/qOdvzKS2KRHCVpQm0sugotOscMRhjoXxAElYPQFL8uwT2wiR4+LZ
w+TejGah9vPPPWGbCx9fALIF66+LkSa+0LaFsH8nUf/TnMrB/dxAX6fpWZJPyDyOjN0lGQUFqgVJ
rCnzDfBAtemDuZPiYR1mEM+almBk42xpVSMeBGQCxF2MZPyejMRjiDvSRZQfswqMhrt5aSSuBMj0
3pkVN/nEcJbs5661vWcGv0tShrVw8l4uwiG5nETNlOffLf19uq+C8vCSXjaqJL58UlebehtCyXMy
jZRyfQxLcaOtFMCQ4rKmDgXux6LUH5C2u2a8THxx5Pdt1h8G4g/Sv0H6gl77yuFzjjoHCFmIsZoX
sXb5j1oge1X8yejgkP7/mbniqmn1cVCfgUFNsTU3rQhq1XSwCvzjvuGv8z6P01TrvAukTD+Fa0E+
eYbbr4c+9p6G2yzQU4RnSV5bPezIiTVXBGnE//He3c9MTLWqXYbN2fnsevsBNMKOkg470iyleWGC
jttWpfkPA+pNcj2DHu/BZwmdPIP4++iOQjrvyj/g/vJlKsA3ThrvYNNze/mUmW7QScb9BkLB0vw9
MesDba9/W6IRdGxqHP1yEYScZ7QHFI3gxHgU46jIn+vyqWRsnrskyOjzOkHuNyQtiqa5kOhuuqt6
RJahTICs3UxSIZQ1f+vaNDZ6iDP/sj5ctYzYak54RjQRpiF14MOxlnGsp5nPTnomQ+jP0Vhx5cI8
ZLljfb3pNrVw/sFWuPnW5HtH0Iu+fOTJqBDoRL1sM7gRN0QaXHhxrM+DxwJV0fqEMLaqNLBJ22VY
6McpawcvTIfaBF/p5ZM9YbDrKl8M9FhEQwpgyE4sIDU2WnrlGm6NowFZG2G+TyS0nz+9XGuCZaOT
glz60MmPJnCCcRpVpV9IMyMaCQoHQl+7qd3zfvHFLc2kU50Iv79ezV+xwi6u9h5DjkP5yyJJCs9+
o0EOVDP+DuxOMqRF0O2y2CjwheRrp23JWF+cR/zH1XAOKpmeVRrirOESaVhd4fP4d2w7KOvCt8Xc
4eqKwqU7yyxPizIcw7XGPX7M4h5o7ZfCrx1kNsZKv7GIpCJNv2KOgLYjiwxBYhKEsR2ChtJovy+r
3Q2cwcTdga/UkbCX5T/KLHmnjE9VoNqfhazjA4jYtQ+H9C8t528coZocJ6p8WfHmdeRUrittj7Ak
a07v2Q4a/P26LfnnVHLArfnSpv3h1UnNAspX+zr4pRV+ZHtsdrCRPCqJmxX70G+78Meuegy7USOQ
iMzQ+v1Qt31uY/qXKVS4P8iYMYYHWLDWcnaPKKCmw7iSQ1iWeZP7hT62e2nBQeE8PWquRXvEHJ9f
PJFFqsL2eN7Zp6UdLaMeMWIqob1dvoVjvtHrj/ZRf3f36994guRylyC3bNS2t7AOR9XvZtgYYJNa
542b3y9dhbs23dg0Q21Jw6sl9Zza2U/FanNHPVgx5JvHTJGhHDuC6V97XCg6v0UJF7MKvBST5dUg
v+scAd4SPkovB1U43qzQeAKMHShUqUS/WP/t6jDrSDU2B2VmDdDi0IwCL3kc422cFpRVHndwZrAl
d8hs8zGszGMAdN1fO7kbzOjfM3nOYFM+8bmTxTyxd5rmzCLSyGK1BYgkmhlrTK9P2iDW9H5CYDPc
kTyh1OAUmmjDOdOyIgM2qjCD6nWByfd516A/cyXGThX+GF0tIefkUT2o+x5RVQN5sF3z9LJF4B5d
Kf6Fwdlxbr/4YIocgJPYZEXc/ATYpikRljK1lFDAO3oqN6JVPjrPx8RkwltHadqn9k8UR0dww7b6
8b+gjhLc8XXo/rJmB1MJtRk3w5A3WFGfM+quLYqEuq4fkR3YG+JZPuu25v6b4f3nYfenggDeb211
Nm2n4sG7a3Lj/R0ZjWQmDMu2O96YAYQX04+RwQkEcXqJKweD5grM/y3HdRXguRWby0IICcoPscIb
C8qsssHmqvX+YGQDz5Ih5D+p3uNYQHX2JdrT8DON+HHGpLpSKwFFXNw4oshglHgGH9V3g4wVeNnU
hR+kY/mh8UFBvfIQFVR20gBDOrAVMfwE06xDI5r3NTTwnsICvBjKEHRqsPfMS4AzL3SuF8ZxPylf
TwUA4dGwelv3yZ53BcInCAQD7EULtVyiLar6VFr9ekWMURnr06PAujTyoJ5B0tJoVi7HQEM3A2Co
zG00ygYH/7roAg9r7Yvp2cNS+DF0vQuFcHEBH/42oKayyCQOXo9R+KhB7qPCHsSwOVyUFc5xOsnE
Gkq4CcRpYuPIuXZKY4u15DUtAKAYZt0Ln3LigdYIRDfj23b3GI1aLE1byfjBz27Mhd4FIJoIie8F
fo0krauOHcW+B6IstG/CNqN7g/UKNVc+yJlEUj6xYHkivnsvMGlBwghqQ7QrVofBAMjD8Jm1S/VP
zlpZh0N+Uy6LVswopTKg5+rSlPXkWbY6G4ebLH2JPzkj9VqhsTFuyfG8U6xF3bUSk+KQPYDbrF/1
LyU0oHzZEIeyvOt7IqdOgb2j/LBoyE5jDSzDteoloBzdV4mvYcFMouxpxIxoPBfVv1H53p+qH83I
7E7QPTch81LLeO7zlHpwwA/wa8NGQhf4QCVcRV4qJkImmgYlz689mX3a38kJ9PLV/h8MlvwD/JFM
60QFOdVAB3xwH/EbKuiiA7xPEgtKE8/4AiBo4U/9HAEqBn65sqSsjp0lRWa1BG10qnZH9a158MiP
czGeNvOFD/HL955tw+M1Lym54f5PmAXA2bNh2fQxRKht/GcB/nNxbBf74NqrfIn9RzCFj2QJemOQ
wYRQAd0QBeZtAeDTje1N6fvNhLIbH4xsrNUvr2t2vlVArIp0PjN9u9B3B477NiK3XWLFXmtC2lou
Cu+TS7h3yXd6WwsZoF0qC+O2e88sY9vRqDByw3uWHCFPw4P/Ltr+jXV6J7PCqIH+rZ4c69303RP9
WIodAQDT0ey3FSC1bPnBBUmAibRe6R1KG9t3oWlsrJZTwCdorKuO16EITItH1lZC20ayyTF3pcst
6mz9RcSqX/VOT0zech2tbhkHeTAGgZrFl3oJDt+wnHU8af0LWB0y8Lhb52I5zbiT9vg0UaUap77a
JYSef2fy+A5bSo6po7CW6XgRFhnHU/+zLeONMUEU9rF9xtWbnbS7HshOwuZrFiVOKr9UPbE4afDD
LLMhA8SOlweHK4uJdK2DWtuE/6bXlLrM/KkD7IYT/bcm+DeX/6xka8xcMcXwEUmCn2N0CbGosQSl
RRDEUCIgC5wHmY6cbaoOMYjL3CrX8hKAHIHFuaxfTY517tolyIhYwuYrRwtMKKGzN2lOwbvUfPpN
24IuX6SZrvD61Nuz0emkK4y7ie+9tztR9J6U34AGcvhY9EDnTtsjm2dnJ+ywOGh8zBGLI+urwwa5
C4+BfUU8v1BSR0EPnyGeSgV1sZTQ0y+IuvmqBM3oMNFqHJwmbkgJBozxwhEMe3+Mp+OQy0Je+/1p
8tFAMGYd/GNnRvQ4DQOBwXhuNPlmkrygwL6vJly97sIYlkDMr61iLfuabu0W6Xma+AQph8j+6zKI
eA/z9qzawTMBvEgzI4GVeYy6WJgNXbgTvM1knsHQtda/9jyy05/0+UxfhaMV6mjwblNurnRTzY+s
/jdq9YoMv/oj9emYc27ERIJxPTU6neTAQRMsJ80nPWE76SZY+wGcbmqHLMnWrXY7kgNGbaEZ6oIf
bis5WatPNrGoMPd748pzfrhNeTRc6AeKliSr8k5GDi1QjFX7TNETle9G+svSPvFb1eAaWPG2ndew
pZDlE3M+4aoLOz1pWr9YoY5fMiX3JA+gk5of1ecpLbWbiVjUPZI/05A0cT/Fc3AVp5rNBkXGjegg
Ls9yardGw/Mu5mjlysiNO5kvhCXFi8tD6FKgZK8bR0aWZQyyR+IQ56Etwo3pAXBwx1zjIixjMkrK
e13quInZHirG6j+mn0EMF9ifG+bnNvokLnnlpu3WPhJV28B0otuDjxNXBpYjDg1rNDyo0yykZhiX
TXtROlio4OhQBkX2M+1MhQlEi9hMt1EUfRnPtKdBTk0ZvsgwJMMfY2mPS56CmuAHS9UrMExjIcwt
t8trCSCKNxHQqVgFtcPOGI0VtcLBu3q8t2772gurR5y6tgwbVC5/MvJ2Wm0AtIT+xLxWOyBlRmiv
0TeXNDAJksGigPhiHX8dg4eBD4KPYE/3IZrw4r5go4WGnPWAoP0AH67noTogc85Qi0IbG+zOLfnQ
KvjsGM7HRzXEMq0VT52EwAxP+/o4pboHl4IE78lgwTF9PJcxNeCCWeVNjysamxTL/C1L+BBccyFI
TqoAbmhO5TURtZNVH7ZkEQEYrhdW2k18g24yZlIXpkBAa+4l+pDiDWhl+h5+YiqHbdsF+zRi4oXx
VVLL3i0uB46lAUBje2kwlGo0PTCXQrPT6RNXzoIBvHcoD4mogELoywsMjFXq6EE25AOcwxpPdA1o
WViy8Szv2xfW7tZOd2O165RiygjhUQvNGiEk3g6XSy5N16kO0KchICUq1d6l2HDZmo81MEzKtiHi
1roF+3QOO45HzeFjP0W7v7xuS74kUkFP0s598Ri8it6R7JMiTeF1Glj9skWMS/tUlR3UwKux6gLw
WqoQMdMsa4unXR4elP/NgU52pLyyzA7jkjZLSoViJl+C0qHYoydg7E4MK+DRHpGtTY8GOeShfQfI
rXurKTBQXaJcf82EBYWq8NFd76Js2c2f+/vIo26tEfA74dRcr3kV+XJFhi4Zoj4ZQyonUda2HtQF
1fR3s8Dc4VgO0nJcm9sa064pV3GPTYp0etf7tCW9CQg6h7sQAcdwE2X9PD7EE1R1o/4j6KdN56Q5
sndScQWoBFOcHTlLpVt4gaot4eB6TfBZ1jTqJ9PwBgTnt5ucj7WDpCslcDlPzxzb6W59R3FQrMGd
lSx3R3aZqGs4MnIWCrWq8A85An6lpVkl5+50E+2zAfakMHHuNzL5Nn+rEpu08/5yCy/dd5OBxPnW
WaiZqpbdmHgfnrcU+ZX3UfgLpPpIZvwwBcc+xjGz1NXyjZo9xSSgDOw+slvwQ/xgeTleg/StmjEc
LKvlSRjGEO12xXoeI7AGYHE9wy/rT12k6zOTxEnFvnM2SvT87CBKz6eiiGMLZgDWkL0LNSeZwt0J
SSi1ye0/FpbqxLxBOSnbOn8pXtg5ZPpIzPnATQM5enawtTdiWXnEI1DMOkXjXbmblJnVQB9fe7vX
U2R+8bPwqpCMDbOsvsC6xDnva2P1wYW6EnxGhzOCHluNw69g6znTzQ8Wb/cvPGjUMPxDYvlye9wE
2MNPUcgv9otL8EP9bNU4ONOXF00ewTu9N1KgjXPiQE3RPZzVSiBhVcqUcV/HzEkJ7/zacOfrkqLB
dV4/zeE+hyvgwSeRtz1lG+gzkqBi+eZPCYz56QnEvZTcWk6j5K07TSWb2eBrgWOVjyf3zbJMRdy9
aQoO3D2QOffP+qB17526dy8SK13YDvtQq2xC7nhm1jMQ+j/+baaP4EvQUoV++vDbFxEl8Ry1u99W
Ra/MPd4go6eRMDs8yt0Bbw2CAF1U+YM0XwFneJpVBeZc1p1+5pLUI2dRoJq6p8BYKJZslH0v6dfQ
d2OxY4wwzWRcTCjNCOjlSAueJeCQva/ZE2qiirvRD1nCC1nKtX9VkIxPbD4V588qpyHZ1ClGasH5
1mZfl0y54PI+9ZCtT5VA5SrZ89nCFU/f5qnvKR6q7JkghiNuuptkY+AK0BaZ3mTqPk5JcSMoPwIL
wpusyzSfbeeFRWM//qQmAMuWbGRLB6vSJCcJ0eByUCqPPUD4hl8355FT9eNudyoCbQWl05kWHXGp
eJO51BLGZnEcTcLwyRd3T+OCrxsyjNZ24n48xRAze2Q/j7/Dmj04f1OgLOoJRo0OtJg/jrHpPdt9
c/W+V/QHfWNiueLIwKK+6Rfw82jPmBiiNtgh1mdFK3yD5ua7V4i3QfwTmAlT36+KBD3MVDI+K4dl
ZyRubais+JPtdFIRwOmWBQ6jVpjT3t8k+/IAAtitTpAjQcU+h9cpbVeYQny5OaaZfHyotVQi8Iwu
N/8PPbU/Swc+/AIgdzK5/ZdTBLTH+A4k1axU2u8QoqjYXUJD7my0CkxUGnHHbrw0h+pI3bMEOwqy
/fSZ6MS/4GDgky62/f2SkQOc2Ylvxw3E58h13P2Ak7cpTNdRzDgOfkymu1G8N8kAaFqS0+0zqZ1n
SjRVoSN+rmQyMH08/eb9BH6jaqsrbH2FgX4gFMKksNPcsUDYZi4xXAzds6QiVw6Bewk3rgsi99xF
tOsLnIhnY+6Q9H7yaItmpP+Oau6Ts7KZvaBJn1PX/hHm1sgdmFrAxWpTuWOnYyF39VXNu/m0yHrT
nMMym3WQhcfjU9pEUtVtaSRZYawvonfq3KuyReEJxxyAGtUDyWLkNJDwYu1MCG/zI/piH1phTDCa
rN8KK3FJZmeNUAda9fN/z3IeHfFg89qiRquINQlXWGC0j9oQNHe96xMPNwbQjar2oJEAYrhnsJt6
saFuU+r0FhPS3N9bu1QH3zg8rBY6B+zvehgDrOxUwmZoF//oKX6ExXUWKWC2Q5ETd6t3Fy9gADzL
I309+tAhuEl5OOgsA99HDaUcJCrONR5kUTTrJAlYN7YMpvaXhOf20IgMRhgFWsHKy7Rv978txRgx
+HQF3S0Lc8NftvBut4R+HUE0kWLOQSD6SOQLHTqAWZT9WaPjZXO3+K+jqzAIMqwAz8L5gS1VPmWA
tX94KNA4vjO6N0No8KbqZRmj1L4w6U10lpZQDubhA4s77Jg5jx0gw37Lbo7BND2HuxLO94PlUswX
kWG2z8maxNeG9OVIo2f1cBOPjrdF3hVFli7M+KhbcZrlZ1UrWCKauvzfojPGRD0I2z+Y20kmrm5f
1B5/IPnWxsGlkLXYgQZ/bHzdhtBCGAd0528J1YN7BdLJLR2QUZlup+ZkKbPUUUhIXWs71g3gcJvw
HeoLxuneLSNWE4BENQ001QM8fTI7TmU/iUaECVPun3tyEJykaHPnVIs2rfM4HHGgeR2U2iLC8nw1
1W35dWYZe0R8MFE7eX2wEu1/u3rdBu3N5x+jtQkUAKMrx6OqGOrSqLGAYw4S30FhYJhvT2eqYMZx
ZeFH59R5OHhJ7+fqtZJSF+BpMCOkkkqVMfVls2uG64jvOCahEw//Y+pCJnZavbsUeyDCpv2vTnrU
PD1aIEX+wvVrFB6kftkwesjl87PubWTX0xN6YsLP64oRMEyNhb8FARtHqbNzthI7ZsYdu0gn9pQm
6ZXVa5D85TMifhlL2ckZsbq2GNEFmHhQoYRhTfOYMR48NG9MnuIlNtyfUhWpMb3eZZTwi6tbgSt0
9Gt/qJKWkzSYER2OWI+ljn8Gxvi5kj+wUcUm5h3bJU2EHsPStFq/TGiF3u1/THUoFEt4gtwyS/yj
XVvAYACA7FoRxqfvfTJEAX2ukKK22CXKgeVBt37I234F6muDzws8V4rGCaCH7yjejxqLPx6tLXjV
ZMXl7Y7dMapcKEsoas3ytqRQQMJ1AXb1YeYGnBYOB4vdqdwnENmFk8AXtxWpkOfbBb1JV0QthNTC
VeibVl1k55LKXBAFBLhzuQ6ueCZCfN2U1p4p36JuxjsBDl8+MFpbazP1MDbl8hNMrOXoR4tODFAk
Br7Qlu4yoNHNXhQiTVuwda+M1JEwzenGjucKXvx2PziLKHhghT1+snKUqveN5BaarJU1m6c9IF+/
oTg7BrLAhafmlaOXqJwQI711voNH27e38uslbY4tR6iC/rtegnSmCODuA+I2hOgI3hlRxy0aW7JD
Fb219W8wCfPU+s2WjwCca504zNZdIEdyTCaBBAoYGSwajm6sjJQusHUw/rWsxODMCf7harwyIo6g
WiVvXerOJMtMIKXlZ6Gjsg2KGDgsJi4Tklz1JhHD6FGic+OvaxKCAZlvZKIw5FHt0IlBTXzxNgQx
Ld+OYPUTAa0srEuOHUiwEHgbOyWd0WsELJPP8DxiyoqQd7avr1AU178sF0FgMhglZ3zrIppIGMMP
zoiUyTHYV+nvGrMJoAZ80B8rHFirF+JN8nRR9g0bDLMghhnSCW26H3qntngp09VRsprAZW5uGMGp
/xLANki9XqBM3xbBXnWRgpoSIFHNOi6Y7LDYkrHVy86/SikyFcxlwobcB3FN7dVzn0es0mDZNZ6E
T3qAKirPc/s8CxTpmyytBMHkxZ/dRGoCfxai3fdeXTvzeABpfwyIPaUlLrIbU3W35AVbrtbDcIZB
769QsNGUq2PUetQGue62Ohtdd95NnQeyconyFW+++OnGHwaRV0z4uZYwGDbso57pBDPH2wPUU9zR
zbDQXKNf4B1+ophHLhXGV7rkGBkW2kl3TFWR3dY+Z0ipQNLYF5BFF4Ofz6bqDvRtOIcfr1pDqIql
o1LfxVMFHXyUgWiYrYe0au976A3+rYDfwITpDQvC0BaYQDzYpGRgl06IamGbXzXHMCwC+LVRnhEF
hNDlrKeeG+LvkZccWnxqpHr8YmVsAV0UioTPLYUfI9S0kIXiJdEjGH/5Xqjfj4f2hPoEVcIWHbTB
TMAu8mhE1zJbJz2IfsirntCMJiDo+n+KZr7+t2vAFmfWGdnPhovMIo6rK9QCiZP6sSgfrRV7txGM
okLsaZZdjSmy8g44enRTQ8gnfyncaNacXY4SzDhYAGqNklty7m8/z+vCxtYwMJ0T+jahAipwI6kN
otoIHF7+4VE1JMvBiRznJN98zo/gKSUZ7TbvamyxEmfr45FH0rtBsyJ9KgQY/4msjD00s2/hIr3b
YMMAjo+bOKIbzZXUD4GPSsctPWazT9JQAniNTfEoOnKFRDXKyHbyrKlEasjSQyzuhbGyFsE1ZjNl
nCY6Nl+UwX1a4JNohOapgEgu7X86xxGStBNTTW0xSGJX7KhVxdKYXcax8Ygu3tTMSvgVKTpu873B
ozmzHYQ2qAWtr3jg7n+aZXgq/+vj7Z41tAqJrcoEY1UGj9xDJFOOFo+3DXjKthk3C/r4qY9tDfbA
kBmi6wtLXdZiyeIJRMPjXXJLBsaGjDXcT1QpjDVWzy2Iyg3+i5vTk+bO3x81BJPQlr0CWI12bd7N
bHDUUxbwFV9oTh5XsLVrW5TpNbMHa1xXmbb85I6PIlU0HewBeXyXgwBhaHlcVEPF2EdibXpum/Bd
SQF6ZADwu7Oisw5DSwr6thWhFTE47xwjbLMScUBUnkzqrRh8bKvd11pruH2foGBLDa/UHKgSVVbC
EzKBdVt7PinI6YioA0wPETJ8ydXnv5mGeG1gu0X9FQbh+Wlb1omyyCoLOU5acBU7NR9c4gH0Irxs
Bp8SxKYgnnTKSw4nkfRmEdscDWixMd0qA1metk9OVoeZVzyJZDR9Sgs1WQt11yEzAiDIBKol3wc4
gt0MPApYK4qK50KCo6fMT0jiLd72E0nNlt5KJxeOFdLX6ETb237w1s/fg44uxuO60dkjXVAEEQcT
MOvViDz7dkA1y7gSOMztEKMCSUy9YDxLjWs+W+Zhfp+kyaT7cmnAtN2OA0/xQ3Z+I0N3pPsttumt
5Pvihojc8bXopuZFCC1ftzu9SXaOC8MT//Z/MmmbFaNb5YK054nbegtN8dNwtl7BZt4lX/EjFzf/
jOFcRHEvDBm8xOnG09UQME/cwO9F38RCa1go12uCOoFgnnoSisBwHKobvbSLhuUF5UYMs7m8d6ST
Nl3uHjhWxwkxs8gZVhUKj1Qv2+RKblqDGxSrlJIgYTFUvnkDdrcFXgvEBGzTiJUY2sWlcJ2Co7si
YuJaQQjcg3GZRtHJ7S20yFxdSJwvxmd+BwupzgpAV9GW9sdnxc3Kxk/OYtLQ9ktEo9vj3aPXUz+7
WS7VDmOO6p5CCIPnjEzbJP3HbXcu0niTbVoKpBa9Xg5GZaWYboCyUvhd6cMPY27/hLAXUIN6b1uV
3n6tPgzWsfC51QBIK1dCdf4VTTlrcNOtouv6mipYSRBKUqM5kJCf2O4h93ZEbJYKy2CyLHtMm4F0
5kG60P0eqAnGYLaX5zSjgoZGEF/uqITCQbHKkXsvwkjx1SvJxM2c+INsxpiRV4jBy/jChnnf0DNv
G/syXBru3kwyUkYEn0YaU6gIu/EFZxMsgb1Iw6tW5aD5U5f9NnvQLPVsJxDjRmmYKTYZGme3WyTZ
psEcT8CYJEkPnroYcyFNcs5rwnVjjrm7Xv+6tyxQpyFUU5RA+TddGxBnNzgHg9BEyYqne5OvAkYF
Aqd/8ftTydSv82lb/NR9sfbWZhqspzf8wEhPYcV3B8N1aYkpOCJYkHcQWsiJpi5mcZ9Wzs4ji6X/
9hvnPsn2w4vg2stZouVdqzd4+H6jTiX3CVkZfAY5DovYgDfIXPD3m8Y0D8hSNi1/ziEObmiP1nqp
NCy9uUUnrIqy3ASuEg473j0dyyHr3c5ypulnSOxpjmjE/x8pvXmPnPJC8bG7GZrWp35z4dWx9rhv
f9+z5eQN5mKPjRPi/vxPY4xv7LqdVTRdHmVZyHxLwbwLIGlvgheAU7Ccyc1YM2OTLt/fNgPiAPWs
GRLJe3tUuKvRMomw4pr0F/yXRYQ42FMRoXbPRMuN9RDnwiUFVAZr2jvU/xmIAQdfvg2eDrc6o/5b
0v/vgMa7GnZ5G6Esx3szgY+a+doadUVmke1OWmpOfECE96JpSonv7/UhCT5NaCEds0nfgU1nR/Ie
Swxip1zEOivTvkicfzQbcypSiP1/q04Oe91vTbKOnuBIpHAll2j65M9uqi8PD9VJ3ieXsc3myuJj
B6Bx11xGoXa0k0VmbUvZDJEKeMO7vlO53476QVxZ+I3Sl6Uajbq3ThQr3gOywrqTRODTCXDR4oia
KY73bidtAczYQq7KWwwzU6eQbW9Iu0quoi/YMlzWV5+VcfmKZ6nIXvkrFW1Ty2xpb/iCLqDaYqBk
bzZm/otfjxF7Zm5vo3S7rdIQbabfZ2VwfAs9tMnck6U5Ixw4e3NtX2um6ksHiAeeRKnvZY2gvxOd
rEqi84XhkO4Vj2GSEBotScN/utOS8WnccMAXZ7YXe9j7usO18aJu0K3p3E8dS3M7Wba7I9EEZZns
qsCDPmV0YIumZZ2uJ9K0jkt3vB77IlaVpeFjfvgiVdjB0GChxA+pSdilcAmQZXj482vUFooBElLc
/XHYFff2a7NdTpJI3sNkLO1e9pO6TDR8qk3YfEkQ9HU7g3IEMibM67JzefMPeaZC1/rEc0bkEaKV
+y4ZPOfPdbRS1HUlJ+E8J79ju10YHqP1s1WDz/k1O1Jdpbaupl1V6KZTvzpm1SaDudUcby6s7rY9
aQkr66gX46bLiNfIZt/R6dtb1ihoH6uAUXtRSsJywJrYz1nZrrVmkjhqDQQnNaOU76GDBr1t6hwX
xDu64h0cH+OyWnwG3Dfs0NOXd6hmAzoQifB3cF1RIfWwCFTXoPkll4YbleYD+ZKcFeqhJcpnkWkN
9lxlMb0Ipkgcrmo7rmtr6O5SG2k/BQsOrPSmFIZN5Zpe7+6vyE+58jyrGUlCZ+uUkWJo9nX169g1
65lUIQdThNLtg0MzUM4ftmPo/UGmlIUaqDT7kThSlduEZTGeSON4cr8vH2v8F7oZ6Ezwzc3p2BgI
rtNmDMC0+7lVp3EBcfMDzmIQV05UxNT5eL1SfeeJkqxNSJVUthy7DmBEAnxda4BG6Zy/bAS8Pn3x
cE4MehI7ynmfgc0LjrbxDN3miDCNKpqNbA7KwfOXar+rPctGwFgcTQe0I3qOhRjtE0JKKkIEmy3a
3jN8Xt2rkuXCN29CrhkZMYB9ew3/IeCE8M+vuFQ5Gr1tNSk1YYysj/F0sz7mKnOiB2W+oChwGdDD
tIhefbk/fumN2nTQuwE07/aVze4QjOcd0gi1llQ9vddkzHpiqWBsJqVEsLPpHz8qO9YiwhZnIvPn
oXMHc08G1mT0xtaLrsaoySWH3FKsuLla+l7eBHUxJAVscpjeUeFZN1uhDcFaYabKSlQsmhYVA0gS
viYUQz+qivIJk9WoT6KjoPtKvolt6qedETrp34fHISGun4ex4+VjUDmY9Sj2X3vx8QyY6x2FUvON
8iJCiVTu4T0qkwPbWzZxjwdGYvGMqa4CqKvCyI39PvCu7Q2UHMcD8oIE55iqBHNc8Zl3ZSn72fya
E5BHfPzmCHHftxiZ1eFWHXdHJHvBbvu3sC5EWzrjTBpwC1rlONj0BSmKNBPMKsX0m37h3r5UpAyp
vSYZq0cWEcOV0b4/rdq8PAqOOfzNvTKOdCWgyrL74ZwEt6gCpXMWjtKYXTXpVASRNd4XTQH+c8me
kTW0WhdLHjY5q0FfAdta8XxSeVvhbuC+O9KiVGVCH5VKlunb9RZnJKpodu7P1EkxjvLXbXLdozqX
U7l/s8vlbTJk9oG8UawyY80xTtHkrg3SQocG6i0gTy5GHlXhhvDfqCwoFk1pjN+PU+3DhtUglTWU
CN74EEnKHpthHHiLQkSAg0oJ29R0MqOwsTXh49ikVixN6bEUaYTU1ENafCYF77R10MtcXW3C1P9N
mDsimfv/rH7pIpsFYDCQpKJQWiJR763Ki/Vo8/3yhqTQ1hydaCXnVaK04LtXHXu7KXo4A7LfuqAr
f2yXkmxLA7wpVGxwuCgzIGYq/iR079h86mG3zqKQQGf4XnwrS1VT96S1NT6jMsy+oexY5+OueBQT
NSERcgoX4ltM/sHak+U0JYW0mFAg2kkVoqo4jPRuLGKK3Y0eexIohpiZolkBtCZ2cufYYuQlJCzE
ZnHZehYBRSiFfCbzoU1rNNljocSzLcg+CgzwF4Z0pLWfU2lWkswlp1TTB445Dp7gEG6Z5Psml/yt
juUksIaj8AlJaKhBcl8TQ0TBWkJb4PfGhUe5ljkooVLq8wx+f4t4deEPN2AgZoVxDTAlgMw+B7JU
bF/l46paso4J5RnUXuyvkYR84GkUmsjXDU4OX7wD1iMTnU5usvhOP8/T6bGI68CfR8kDn608PU2S
iEw54xJ5FLspUTn2itWFb5FnJv/+NvUv9gS/XDz7K8Irok5s2yRdQYfATubU5bk/naIDswqVk2VP
BDVjREZq8rJsVQ03IDi/VvoQvZmdpzdY09/uD1Oen6jbQyWIkJpOgE4LUl7PxvqVDdW1qqMdty2A
Z0xT5i8uxTlGEQZI7FtXtNS/t8OgDR8AZ7S1IkwkbWRJTNym/jLUlOfxiGA02YQznjSjvr0LZ+x2
hVmUCilJgqhVzmnuFlUNdmTi8D/h189935/cRC1c90xKk96wAX60B+LblRsNjI8brgGOGEFyUcP0
IG+i3TnJr2U45B515h0gld1rUQMbAtrVEvSyl4t8fsOLa5LHRsBUWnSneFskPQHS7Yrbdq1mDwav
jppBQG755K3jLQPVKVmVbg0eV43OS0JixuAaUKd7zJAb65XDp0KYZLHLHS09W9uqryeMhlDEoMmP
RFsJvz9Fq20Iyw2qRRlNWIW4jBpzqZnxORPA1N8ereFLTjs0GssOSuI57brnUnWw6VT4gGE9e67t
zFIX9UogG/nDI/fphTeS0Rr/aH3yOi1UjTMGXONDbQ9dpSB43D3NyJacWK8W2HxeAXr2+kJELfYh
tDBA2HtFYn5bUTTuQtIvPDo+mz2A7WLMsJWvI5YBEevJO1MLhnM3gMCn2mGM00xOAx2wo7HUEdFB
FP0psqlC0A4cT+kJiyA0x8fZOxSWKUY8AW6OniJzpKgXzqPjTNHImM5JxMaHPXZzoM2x+E7maq4E
ThZA5KZS4ulw1PE1R8+p7zqU+KUbulIvuX9tuyKrsH/5I/ZaeeMZjXbbLr6liLHxTHjVP9wQ0gvX
VzyVbjQI7K6pJowaAsZS25o/+xxMufvy9KLafA8tqvtLAQHlZJy4PJ7CySBkEr1VphXx3jdq6UMx
Uvuu0no4Yq+bulzBqn4vncQaQhTJD1lpdmvlzlquSRNccA67ATUULxxbgdbb+niQXuk+j7NrJ1Tq
Eaagz5ZPYqbFqtaMQROIAU6wOl6j69qqb1cA6AunnrmSBVSEKRzRFcVz+OhcfepmX3zgsbL1ySWT
W5EoPlAvauJXyj5gRXbXTxZxYBRwDq23oPFCfAmxNCfxzlZc+KPuYaKSFPqz+mBC34kZxBTr5Ru1
UugWOYkO1GqGdYaBqs4PaV+PWXjd+e3Om8UxGExVl97ViNYUHgyhaQKzu8POkoU7KsVUS+w+WaHh
eIui/bp9nkUQpCN6TDMYyzzUtuIfaIel1O6QXqjXxOduA7ZEBUUgj35wt8EcpYAUMuRmojbcSimk
eYasmUncbt37sJ5yfoVcVLUeYjV5ufozFLJv8VsRm2fh2ezyfHTFFTQyYx7CvIkt9WeUjXzzloAU
pKLJtaapq4LhrBfIwcDeVtNtKbIjNED303QfFaz6k6O2D33Lz/fJI/AACyx4sWLuMBbWzlOa+pu2
IaqXvEsCIrq2kKogSt+pJcceulRpxDktwKz7G/JjGxyNwzTW6Eiz20k0h9zoZj8pbA+0M1k2LOe3
llwon2ITIPyqHx6m4GQG7RqxlGn8I/gerH0I9ocGV7n4soDrb+LL+RxoGIqrT19pGl+LVHQbYE3n
WQ0Q5WOKpJ66VB3aw1Vj832YuTRgM4nEIeke+FfAJqBrZHGFLHsHl06Cu2LGQhKVJzzqh3zIKJy8
I/5Wws1L7kSXD+KTTdOY+X9papkSUfFTO6Q42Aks/Tcv9LbtO13Gs3apyVWNKEOiPjAs2U1cyaJp
hH2fkc9PbtqsF7LxHr61BUMjg/9Sm6OOZg/3Ip6FTyofw9n7+Ii1uU3YsYLTAPHGl64W+SjZRhd2
bMJ+NsQSjARTlNn1lKj/1yDY6o7R//jijkkMAezSbU+wkBmSQCIU70oYzTKBeZeiZAdD9zV3EPkW
65/d6gQlLbkRYlPdGgUFYHeYFoEj9udtOS/bWuIRgNAzfLDW4tUvvAGoq4RctYb8uFYQTN7NzpbH
n+dR6D2j0mNYvNvYbbpl8VjwD4WPyTMWe1/gbRNmipYPAyR4I5XQNGJB48Fmkd8XR0pU6F8OfgUq
voQck98bsHGU2oapz5HtFq8pXETx02Rf/IJzd1E2kZbPCUsqEFSHKkSQbYQL+GZxh+6eamwQBniB
L2+DDU2930Ny6ONTR1+0QLTtX6l4B5e1rLI0LaK/ApOKYEfC+w7/bOW4vneSHGce/hnU2LHUrZKN
LYCfG7n/BL1Ma4NK721NHFm9n3EV+T9xygsUVdJVZ0uxw9wJFLnkBvEFMTJWFCAzcX/hFuPpMRR1
onlCFYUmlgnKS9ciIILesfvMkG/EqbECbmjJUqE2z0BfDoZUHzE9uqVgz3x/c4OxoKwwWoTYKMgs
xoWwHt+5T0WeGHLbjQ+FEY9iu4Mwg/AvBVexUThcF+lO0aorwuLvoATeUuCTlYlSexx7DrtIjkdP
9agwhefsh4N3fP6ljWUOjF0iFMLYMXpb96h0DPc6AunoxxYm3fKtnzs1Kja5t5akCX22AQ9GBu2n
dnZpCMeac8FXyFQab/80+zVNApdeWHHT8dncN7gGnC7N3NjyihtffBVj1JMnIIOz+K81AcnVzM2q
/0rqPpQPBtXsFib4ydUXDfmsdxvFceegy58lkLoo70G0GExNDb+2SLoE3w/3DyYJGG/bU7cVZ33I
CwA9myT98AHzkSrMxgwdUxln513kRroac+oyAymXasdMKQGHMsfybwL0fpWNXF4vIG7Vs9o/p3vv
GHrM19NStc3tQ7m6Zu966FhOG2Z+SxpdMyE2A4pccGEdc8jCpETHFdybsyhj5LgEJ5s/yME+TuSs
yRgdLQBRtnfdxatpdtfpzOZ9bXzNYyIWa/ka9pC6dVplNPlPKcYrlKVhuZ/B1+t6oaeaQw4GJcJ4
Jt3K9yUdxHWU9bzm4nqc0T8Dc7QBVcXJ8jhy/w6l4gdstI8nVi4PprmHjNbbho+VZXo5Z3GvAJUT
hrQcdYjH4yLJkl9LPRrIlVqoRVfIIWdMtKQ2yHyL8Ss1dG8XIEIUO1gxQ6cRfHkp4zCotL270NgT
C+lh/jNu/YL0Nicf1kBmSAWz8+Pw5mrXfENr4RSb7eeqq35IV4YmjauUkOQmbRln6YDauv7K6kkv
UQaWFhmaCFrM3rMkodRLLA9I5JaXAeUbNCUkFD24/PvYaYxZ74cwAmVrYhgphX+SVcYcEalo/JtN
i3bGU2KhoiiXCaQY9xgXrH6Kvys3X/XckdyeLmoaRqyxfeoqbuALSxDqhf3dLJEncSqMj1PEZuvP
zsHBM8Mm/dDq+p7Vc0GG2IykeVtT6ZZ4Z2iIsFsQBXYI6uehPfE/w8T+jFVgQk18xbVdTGAF3jlK
6pNM2g7YHWELCseRJP6TbIqPJTms8n/AFl41RfZ0asQb17zy9yYP1Ob7lEJMAznSIoyjAHLXx/E3
lC1jvxicMtiiblSvotw98jyZHfkUYAVeAi/pNasveYzfW83x4LVgamCYihflcke4KLwA5vKunSzs
sEHLYWlN4MZvu7/8zvmoFILHFJTP0COzOJFV7twvLwxN0a5PHYfag0G5AdPRdM5dPTYesQ130fFW
Q7/+mMZIM4/B40SU6O4/0Ww1OZpYyZ0CP+ipFmxf6c3uCGRwznyRd20urfvK9XVY9uNztKfBmylD
phZHSDpUp0sMxMEEnE0Tx3jbms98G4G+rCdbBKVXV+Px/Ufgz7pqfkVOgRJf0uj+pUOquFoBVVzE
JKH/6xNTm1+T7TkoJ/1mTIkGQJIWe5XKUVqgYewJyGCEkg1bynx/R+yYYf4AKyvSLuGkM/izvYaj
ODfX2ZIBdh3D0hF03uy74mxSbW9OFyP9KxPGjAKqaQazFOQnEQnCs72gPYgZvTbqp1vVNbCi7h4C
LIIzDA8Xjl6gOa2CznjdPKo3w+wZ6/4nRe2eD9mLnPb+gHgQjftHoMD8r3UZ0+Q8xqcAM/VS+4IR
fhrb3ekyGmOWcOG4rTUEJLXTIgFvA5BQutQao2ezTfXB9f9GfNIoa31rzlzq0aAaRp4KtuLc2hik
7fP+guYioByVt5jDrq4TE3BoFam47z0D+HE1xt/TXLxoIrCpmYZj/0WUcEzNL5XFAYT10gw/Fgs7
n7T0L29oKtu9jziV0XaB0cnwBaVoCldyMbdJpBuAdZLJE/ds2dY1cIKR8At1DurNJT1bAdvI+XeB
RQpdtrjrzPjzzQ3nfzLm0DEIdDaBTo4YaD1FGVP/2kL8t7KtrEgQxAyI7Ny9VpQdGX2krSkz38uV
L4mU2Dw7DS1E8vkvcWsCeRPvhM4WNOuQyRR93hoJPEfSEowIdcXa76ybCDlgkAwejlG/4qZ8B6V2
fLayObFL24fqXdalFetuNs5dYihHkZxBP/hBmgMv8On0tMWW8JHbpRyJELz3GM4AiktHzY+9a8hQ
KN/52oK3fD7/K8AZdyoIftmvYRiulNVo266JMqSy4GoPaMldnT3oOkYoQ33oMf/hDZWHiAGNZkAR
3zoJVsuieyhdgvCcEl4njJMzbml5fuOyJ1kUGSAWCWUpVXUxEHOLiGOb7C6JR6NlQ5yx/ptQD6ts
avi+hZOTAV0yGxaBRJs55z8JMJWyNdJiyDjgSgBr10D8dLr26kGs5gdUgVoPZUIACb3kXQjnYJLF
iTAeivG1Bvm4L1r8CWDlZDhYECvg4nZZnXQ2LtFCzobU3xbQbhL0028PpMXY9CCrloevwr2Un5nq
UJXANZNH9de71Pil5lzKx1Xeuu2vYsP0fB5RvtZbKs91F2bi1SH1ot/PPIVn4bewnnHOP4Hn48q9
r9SJg9qS0jLC9jLeVHGtUqwxup/f96n8IrFc84SbPZ67u8aP9qOS9lsTeFmz6rLbGFqqgLw3Imbh
JqGQdR99cjflbdztKOA5SECl+/nvgm5dcgSmOHIlGSsBJG+ZntyY/AqprCL8jtWTnMhyV+hx5EMt
FtO5tiSsxsv82NXv1iPzwuU/5Gs9YBvBOKdn8dTw0BKhDXAuhUddZrpuRhM5znx2hdsDOlBLXaMy
HGn3zRk+gNu2OnCMoyg5nSSMbTksziSn0jDoR+mClA1q4UmX436v/wPscDcwHllgfV6yZLtBu29X
YOvJNMBnkABJ15BtWq7y4BZvdxgR3qfsi471diBBWRE/Vhw7gRf/5D9DpTBQjt4e/PALN+VGqeey
yfnMs8wfbh9AjPCzMS+wOUMitrKpRquE8S8QRBB5Nb0uwyHpGCoHlPuBZZ/+EFaxfSUY0BV+wmV+
sPSVsqCKw6BKrZW1ZGvVohQzCUQrkP27jv5PXRphNfGQYRSsrSPpWgdRh3VPdBVxT9NlwEw5pCmJ
Ykd7Y0DDklBMaMWKf6QGKDYiqPkT9iHWkmOckbTT6L7Wko69/+OmwRic22+lGre+4aqMJpTZDnf6
aIs6h6uBQAYHAW0acywR7kFbabLAoZvzzIUB5ocrt+8DPdM8j+YJvWw4Nal8Ho7JtV2z549QgUC0
yjG8X6XTVBDGIC/o56X+zehA0RfiFoig6XG5IspHJ8NZsDmSeARzh3qEodrYylrnqTkVvqYMnW6W
SJWJTvzwlKijQ5Y/+9uducm/RdZJ/kkQ1tJjxopWlGnhHrsE5Hf2tw3w4TR1Iuh8IgTrEy0mZQXk
KFIxwgG0ACJz2EqeIxdLxeDrEEJGQroZ7oGOuvXH8fLjI8pSpTLOlpiCnH8ddOADHffYiUZvD3Td
4xQsd2jZxnp6cXxx/2YtomNHpp8MNgBkhRy/xc6G9Vz+lEgYvXlZ/wdyJl9GzebPI/Jd1wsz/twe
piQkqDTK64cXzgNy+39NtAQVb3zak/3QvgbFIc/ZsQARgDPCmeBUcoI2dRrfKtBIHxc412dCy/jN
uF90VK0EQKdZsIe3Lr6V2BW1AQTi9R1NQOo2StJ9nAwoRQ540Zl4VLJwvrVwmQrpscEMCZLO0N+F
MS1hrJmnGc/AaLmvaA+A0AmsLNR2SsJmK6tJe8FH1G0bNVPFesbZsiFuyAovuOV+VcWA1Glkl3Op
f9/AifTWQY9kFku0xTCqznzyo8jrQoEAcpcTzUS4bCxnAvl0fcu0HgidvZbQ/jFNcaWdc87TI2DU
YnlIPCU2RX66RWxqr+r6Pl4PD7bmH42Rl1wBq180Ei+lfMch+iSZcE0S/BQUlsZf9zmqLxMzaK69
uoywmEF9ZzMagVrB9lLIhNufGgYgTBUnILAMElnPZaLu7EU7TR/+rSa9HRUljBfREN2qRADArtQV
6IIDQ891zDcI8bdUFTxSQeRyBQJ25ExeLChymmnG+bgCsNPK/AVSYGGvoBNt2e49R6RTF11v3aQz
Cc2wYJSZtnAPg55whZuiogQJ85QpsSmI/al6cVKctioTikC0latPYWKYZdfilTl0m+zO6bkjQ6QJ
U9WD7410VnBAXTYgoVGZtg9xtL+Kwic0pWz0nye7JxTtd00X+WOQe8LRaELqmxU8g9IiX2zImj4S
yw85/Lw/HNdMmIwV1mvY/lKYN1ZSp1CM9eeI4ZDZ8tl2X0pvmD0HB+X53PH4Y9FIJI+hhuJ6Tzv2
D+Lr6gZG0Yv5rwhnh5oQkZpuCkV5oobD9FmmzZ14pZEwr95yqCG/UAV8BWqo4o1Xn6/GvqtzTGd8
bEgAHsCs6AL8wHxLVqhGLuQ2xKaz6DttKwqd9VD5aoyn763P8G8aHVAt4brHQkOPVo6ia9jIWex8
r7oJPj41ZPkhFH6BmT6OVKEDlj8IFK0LiTGQ4FAm/mAqRC1Oskc/QZuFjtP0YgI2w7QylpVnNhno
VMknmYeL3EDBxBlETRo9dX6FDnes7xtHAWVEIS7THABkUtMrIwGmp9pYDxoPSpMgLvtgK2C14wfT
PGUyrI5ABIM2v0mT5YBIokBZKZnwve43ye68AIe+pFQKNV8j6gZv5lTI3XI1YmvfLOEDqVWnQGgp
jlZjPYSNuWYOm5JcElXDcmaZLFiPtfLiZS3BFmJj1xJQHmPGhutNwmUf8CUfqCP1mhChFuDf3ftz
vQockMDFcJno9S3vh+QWpyFcdul/vkC/TPGBy9U0o++PwX3V5zbuBKJS+HYgryvpgZY8acEcrRSk
OaaPuWY2Q1wdGKMGUkjqVD5sN0t4bQ6cpQO/IfxHPDmq40v1GXckK6KqlRJytKf8KjkbuQKJpX2B
Hy3awt1jCjtBAXqfadgxtKtvP0r0njVLJuPa+SW0fS0aFQ/KkuHKRdlBVJBrZm5yBYIXgtVAk82S
t4vZAmYodgKRESZnw2XDLu5WiPOgk6LY7hMHoGGE+Cu44DFtOOF+UQeZ5scgDrUKuc8+TW01uNp6
yjSlqH2TFuEx2H8v0LsRMhb5ppWrLiTPB+QwNluBl0C3Z+xrA6YdIc8YYZ/dzOp1Tz4+O7SISWMg
sWnqTvEajxujPNgUXrjFY3Exu4L3r7KOGRMMm8eFuJUxapI1bqGJQ99XYv27ozeFyJLEyv6lSA+F
W++6fa2HzdptcN+QbG/OxvBOJFbpseB9P/L8wet0W21/LOEmkBEtPnejNyKid8sANCUdI/OexptW
CTVitjzv4fYctCPQDA65KcXEOANouD937Fw3wSgbRKBS71jVWGp5MOgNt2L4FY6tnXxZVDxYwMh3
KQMd86CGWseGzdrrCxG4ISOqwVMLs6Lxuz7/JrcEhFqcQW1XVPgzHsYAaXeiwzSrn8AxKUYKEWSr
GCkKeszMd8qvj/9xVjff//QhCVvekGc3C7uWp2RflkcvI/nmah2BrMKVRrSy1gRLTjuw94V2Sjsh
sWbvRuZ8KwYRv0YyN581ZojCTdYRf7Mfr5OBXgM38I74n/jZmS3dGMY2cB5oFUuUJEqhxn2ChoRX
uvWI46aH8zSF3ZC1XLItPCi+2tqhVNFxyajTGQABqsWVxW4cVDy/qGtMzgc+bV1OSH8+wCS5Jpgg
VwRaP/gIliAYpzpK/yecwmWxPSzTVFzKzE3Yol8BkB8qsoqf0uXeUnkPcyQgQCC67xYBpC7gpTwn
FX0/SYGsjRIW+7FV99zykAAFsuds76ViVvdiERybLmh7N+1tDC4TI7yi7mDPTQM+dM74nvRr78hy
zDSadQNHSFI8saMMKjf3jS0s41nZLDurdPhoraAJkh87nacUk4cJRbQ8HulgNw/Ct20OQKrHPcxl
Yv0kzicegpllXr2EaX6XWYBMAszlVx0Z6yqj+Yb2aJqfwCdqYqs3PVGIwaeo10mySFLfYMjAJhM3
nlf8+e+sL8YSbhshNx0JiZTySYtfc1Ey7f6av7cHmYHf59PTh1Ax1p5TLJNybexp2eyyGnrbpPp0
hks66UvhKb+Xh0co1QDxq4ESfQAftGymfvVnh20wEWgqaQqWQQsP0FT/yBedxAs6uCLTGHHci24h
eeSsMrYX/zP+syUxUBxSSnzw6xyk3VPp2Z4Jw4tMbPpxubiMQ2KVhYhI1sgIn2NEzU/oiWmCxIEm
z487MQ/BZGbo35sZoacaWGdKAjrdFBSefTQiABCVtY/XJuKqxTCqNWPhVhqjCHk0a2XIlsplqUlK
Es2PDb9BoIWIQGP8+CZ5N7pr0PJNRZ94yZ2CO79skS0XFIELbSEfYf336PzToqt/0grZVYhDcMco
Y5DoX33MFwYAtUePqs8U6Y4vUFRNZ/ZEQQIMzLpNKN97lB3LgGjU/JBaXSu+u0Foeoko1UKhgFjT
J3XNNKFgsVSaTa0FSpV0+aHI2tML4cNtFp1OEhvZ3C6DaHm8874G7FZhwV6LAXJD6JSqwFrbQZDr
2VFPreI24o2dOTNGFdkEymcLuoiB033zblMewA6rRhcZGBXY3xD0Bj6VeFdsTYwbw12gMV2Xzn/7
IdI+k1oVKqh82PmsIQWtTLiP39aH/c0LLDjecLp6KHt7XrodddOdsnRDWQviTp2n2nJKeOgKWCHL
MmmzVm8Z7puQLUWnc2sMbdVxoCXlr3VnU3nazf/mZeVT27mj6PAAH74SNs5TBlELeT9JehbQknn4
9vOMyAr76n88rg7sMs6kIN9UAO15Q79poXfQxv8l421fJsZYBtAg1iEjxemU4jpGLwpb9JU6pQns
wOIf/ZYSmwISA1pjdN3eLOBxvg7R0YFxqF+se5HkJdig0yGBadVtDHIWBCS7LocQ6S4w2A7nxas2
Suv3c99l0HzEUJnvd8EQuBBe3vutv7xa+39YruH3REm6a29LJLohMwqQS2Ays+dV1cv/7i9yzN+X
rSRSXYJ5kMG7PY5y/rMPEIpa9C/plZMgY/Gt2KrCVYViQk+Xlitcaju+53S+EaIiRfZVD7lgEPQX
X5SaBEaUca+RE8J5vfs0GFibNUmmlplL02uQQ0dxBKldOAhaAgbNRb+lgLoAx9FFT2Ze9FUz8tBa
ByisrBF4+Zeqf52jptkYi3o7P4aEyARu0z0bF3Nsc+IsCdy430XQ70c/WMgVv4bf/PHcZVmBRfpL
XxKCLtoXtDt/xRY8im5M+JbPc5TT9a4zArnUSbA0egf0Q+0K8ZWfuTtrSL4qYOqYSvUY6NydwbLj
129nCGE0MS52dIXGcG9nYIF2HdRLDbJzPVhJMKqvvmJyQ5i76gOS5yJKMukI3BViXCEWG2uOohs9
A9bf9wNMwWiBRqHzOzg4sz1ngVnYDLUjRnITjglSZ779kTXWGSGeBLwKWmppUu9G4hIUVCGturc7
h0iA6ZQnw2abflNBg7rjIVbyC50tARdyjSPVKuWr5egHwYHM9DcVAXlZD7H+/Ney2ZPALhypr+WQ
7t2Vwytso/C3NV5JlPOOYCuFNTF2GRNe2DWDVd4Ty6HpPjSrCYbvlgH08TuPfDlvubacYjsV6/sD
z9CgGMw9mBCQ85CrWcMjHyxGo0RF3QacDaoC4BCXmOKxb3Qpu6kblNDN4V3NqAeSUvp3a1Lz5GMw
bC9MF9Tuu76MtAvViPrf7DudPJSd3/hWcxn0g/+WblKC8+5gZmpabv2R1agv2pYHWED301TEkKhn
vkQsu/hqOp8AVuy7vpOvTg9jVdcBGMCIiPjGvYywm2hA8dt+w1hKGRC+qXU9mQWnJKeiJqnnMqCq
RaFybCVtWLVSVlRfeRmS1kHg5v3IPYrzSNEVL0/jlI9PT/snhSn2ZxKqauvPBde/U3pnGADJMv2R
3j9p8w51vaOPv2xJ8efF6KwJ2Fb7byeV2otao8ywG3jtD00Eat9b5aJ+fQSJe9M6O3dZLf3jb0aE
K2QCG46BORvqXpKuMjZBxqfA50qnPDWQsZaVXwl9RmLppSrHagRQNXCK60D3lWTQoGF3XtWC44J4
ovTHF46AAMExLpb7DXveHHQdXf7iXB1TCuQ8MW4lQhDfGjxd1W55giBejJa44AEAt0ZZahm35iY4
IgT/5hOuMxRBjPMvLucr6fYyakSGcW7FP3ZPVknu009ypZt2CyPJUc0Bt0A0TYgnVV8gL4aIsuGi
61Nx0HzkBRafRU0pw/GxHcFjOfBx1k7j58QeKPWbjozWFaxzQQwr0gV5nc7hw6+MbXPJrzR5QOtD
4n16R8K3l1bP+liHfSFJjmCISDwJm9xJ7Jtwz19TWVfunz8ofllWvLdtr1N8XLX21FbWKRRuayJA
wXyEl6W4/XjzVsUxYu/YBZyAucsG6sBTEmLEQL7m1PifsWLa1DZQDo/1v82NnGRGjJ+vLYui+HoH
KdwQEaAYQbkEPH8fVASBH/Ym0n1ywr8hhlkIjptUEDxKsieSRaqHDNnrK/iS36bjDcmmPevGlkMW
062TY+psn+rxtErKXwsUEK+3xBExnLdVPoGfroqKmutRtTZq2egyJ/cojsLz2q0TEPusXZAsoPRm
C6VrYaiZ3A9LfoN+NjHs21GC4cxbjyKrp8luBT9YVmQtr7WRJT9qG1vn+st+zB1LfEkxg9ytSlpj
fIRv0RxYaTYh8ohM7J7BwuEcRnyJT3Tg0FCw+QhLwv1Qau7WdPpKek/drmIF/O34RcLiqZeyYLNP
NepNEqHZsNi2zWPLVW9FL9+JhZDFrVK/TzMJsDsPOORxMJA8VD9bTPiHOlySPEjGgo+PZqfHyM9P
FACoQciDBCL+n24TTP5ijuNSeYGtV4/pOFI3XNYVto4cS1S8g1gu4sdigotC5myYygLvJ6JADSdp
FiSsAa1xDB4p2R8LSe6wwjJVcK3+D0bVNUWni95GprPcmCdvHubQxpUhONdt8HMFRerPBIqHd0ob
dBscAt7e+GKtcSZ6DsEuVxMSI2RuzAXhXCZCLqFbj/iBBwRrgPVG1d31wD7uA5ImiURS4Xlis7FK
N8gBynMkpNv3BKF5IgBnkNTZ5oS/GzGn7BqCTzBm6MOnZzCzjv2B9kDgBHzC3gdCgVVKFQSONT/+
OdadPs8GiDMUjMCIL4FJ3DO5QAgriQHCWHdKjSUyYYWSivTWOwUWA1xblUGHiPHDCmY+nNg1ia+C
+KKRRfMGChlOsKVmk6TgKMSYZ8tOuZAURrJNNSA8nf+RqZ0CL5NeiKw7Fy1BSu7sn51+VdORKHdz
XLW+hbqVk8nycWA3UxWWMivo9liESjSapmOTerzUqjweOwkoTz1xoAuTBz5XUNQm7PPaOvaWin6g
feojhqMtG1EU1Z/7xwrvfZvcd+B2QxA7ow9pEzs8LVsfOlWcY3q4LCTwb0TtXbiAaYv3gGXpWbWl
6q6fR4PbCEnDcRRjGbvPvyKKyv6r0QA6xUkmKZCyUbvB6D81tsMSub8AoM3DxClY+FFzkilgBx37
9IiMMmkQ3j+S2Sg7z8mfQERHrT59rUGG52PGlTC2EliBFyqVEFx3M7+iKQu0Zm2ynm3qdhJiH4GI
wOiCEeYomaO85e98wp0wK3e2Nj/WnFDobP44omGRrh8NE2vWnI7P02dMaAGioFsdbHrZYyZfuzyA
eD3WNjJzHCg7K0QLN7fcZjqSWjFOffeDFIEsidMgNI5tiHGTkpt78OQkpicMf0iz39rcoB9cob4A
UPwGycGnSq1Eqq+ifVzX/tzPp3/Qlaxa4OdiScfk1VNLK3KuzH1fH7PzgFq3mTHYwSUTZbiycxiP
pbNkjHZNA9kgPWnKp3IiMB7kX/rHNRI+aoEjBS3d0HYCTxgooyzy+HoW/TPf1Scp8yscK5qI0Wsv
r0zYw/Rhi3K/M2bjDupC/ASbHCbYuyyaZEnhabILGh8rIqaC0JfqLHj+vl/VOfevKHMoobh8ToDc
t8hbc8ta+cUbtI5SorZRPYaMGj3AkINJIQSXq6NmMeMglrymoVJLnbZKgBX4HN+AzfJeuLk4TlcN
DtwNjSbG5fhxJZo2gwjs/kkTRDZ2v9eZ7urX8ZsPI6TRMKxAFOXUvn2Yg4JBdwsSx35TjbRtbhQx
BZhhwnXgeQYj9zoQXmH+uVtjGI6PX1nHGaJLac1dPhWDl4fKSGxFTUhxzXahShxVHORh3OueItyw
UiNoImcO7Ckn4CmLPvGFIrjBCioNJLH91teGGEDeuzqAMPN+bHqz/ABiINma/o7bG67ZSak6+iZ3
1tj9rVNjH4e7lxgMj8aecQKlyf7XAyOhp/ZWTKoCgPwSfQZgl+0PHNac9lckWjGTV3e4V/bIwDXZ
3ny8+muh4qnwa0dvrjsk92XxdKsg3/79RMp8DdjJPL4FY4H/3VEnOBZCHu/hHOIttxh5SqbiOwn0
ydgRCPQOrv3NHlZQSSVI8HhHupH8tPSCrHTQHkAEnqk0rTcrwZv/gJemKxuJOyIR3rQwNL1xBZfb
UtqNSikIzsZR36xyypsQ3Tt3bYjG7lJsAvPyYVjS3y/rDB6RRSpf2Vu054c5LbvrM6L5VyssnoJd
3qELkSHBBsAxX8vjVRrEjN+g3OsvCQWgUIpWstptRbOrL8lr3T4SAjCGnS0v5Hq17OxY7eu3Caip
+pQmuXiJP9iKAhJD0JDNp20JbJ9rwyHE7ZWLGvzrQGbS45zfY7eT/uLvbp9uI/DaL5X9pcOQ0sDi
7WIKowqpzgz8C3lmsKTBomolc4gnNsI3SbxA4GUoGerxiQqX2fCulEtrV999SqzySiXgyukX8R/O
K0q81N+qdak0t1HJtiM4R3CYZC0wMPDvQurrwhmq2iWybisn75zAfpMxKmKv6Q2cO1C6uaAywd3z
3Va47D0ofVuDJRRdj5fAdOSXhnB/mlYtZIAP1QTbhqPYsPxZogDsjUOKYNVFODaUksRRuJ1SviIF
Vv4JvbJGr2mtqpgQqn2XnZR8hcaow/ABrn//jxWKP7CuS4v4+VGptd24kuQNX4x41yDFhPRVjoPJ
dhAecNzOKIN72rEBs/27Dbn45i8XBBPKPLN43xwFRmHsplcY0uNeqidxouX2Ne8e0Zv97MC/ARrA
kfUfqL8cjopS2V/9hbOAYsmF9wJ629UKei5nu7AOGpJ0GOxoF81oL4rnBjnNGNM3xgEFRMJaRpE8
INuXodi6HiFaT7dUg/PXk7L20CCe8xygBuIextnkXcIOx8NpbbiIl450cxrRBSoPTe7biOCUC0H1
X7V95e4oBddmVHXdyR8aIJdOGd8Xq2GHTlnErYnseDuTo9Db6pCXcWPORK2iqv7bq3Z/bxQskV/P
iUvOsy/Ke5gWFILa1A231FqgocH2n/5cBHEZLC5evDsW4HnmcDZjmtr/2sbCd/ehGoi+bRF/Edlo
6p35lf55wOURmrtmmP4moO6TcP4XLHXkiyChnacDsFiaACACrVStrSwkGRiUxDUs4imRX3GmF84s
NjmviLG0C+dt0L51eoCSkBCi7cAbgFkVnbJvhOnzjVN98TpeQUnBug+E04CU2Nj7eLp8uOmFtx/e
e4hXYcGrdV1GuznCuAILWZHNP33lA1QmuWytFz2Puyz8tsDtxGiPL/Hl7NnxSRqLS/6sHC77pCZk
0c8WG4vLvxJUh717v7XOfW+CKLC8Emd2COfoJwb/1QdQPfwZuf8dw7ra3Lc2KcIIki94LM06aohq
vONqu5jyHAwCoOzhdHNxqwm3AaDBe1diovyeAv3ug8P+Ir+LoXMsUh1hvTnbOMo46h2Mgzd5pEkl
O/Lrj2LWMMtCEKo/I69KkAbfoUzlAEsZdJXmC1umYdCy64ZufoaEgWH0CcVs8RRmz1Tgd1KZ7710
rV2izJi0xu8e34HvHNr56SOuFETv+Jfbi3G/s/q9QGnMreD9kiPl/iAv42tjcM1ID2Lu9f2+O2I6
80Wvq+ZkJl+CPyOGbS8WmlSMnPY4+ru7LJM92PLkkL1CiCC0lDoZky6oSAYYGZ+BcOlZOYI5Dx9X
mVBfEqFUjJ4E4j+nX+wnf8/bGbeJmAmIbvgQGSvzrl4fWwiBdjvonUN7Ak+fSrEP5nj49ITBbGAV
f5wz50rWXm+1fG+azQUXUx/KMndjEyS36BFNaEywi7P9WtKJkKknEhNbUk7JOVCqK2acA8LCbIz/
xRuKGcsTPbdArqTIJAqKYyTA8+oAboQ+aEkFuJkixEpVGuDncTXLpTgWMjnibJ4D9A8gbXER0nxv
svmOXhRy/y6Q/wHOrrFiWsxyMyRr9+UKLjK05wf5Qt9RSbfq3wR/7B/NgeC1olgivlM1qIKzvg3K
Ucywe/K0lA4r7x0O1ZvSV0XGqGFrG72mrv6QOmAAr1hv7PuI+dkHDzZhJsEFJjLBu5FBAp7U+lIz
sHqdhXbyGHMrnuaUxtviFfYWscUUOt742y+RjMaJGncVFHadsrsMBDliehK96F501rjOnhNf6we8
GP9A4IeOk8rO8HLzHItnEOB9T5NBK1za0QpQ6+1YPyEHd7QI/sW1/O/6f7idhaLZZHeqd7oQAWxD
xFgiAr6QIiisjjFnF9r+JxVYwRWnvHbhlR46rVeblkcH+WFQDX7lu9zE4s3MXabkTT5x+KC8LAn2
59xL6P6fd3jC5WO0sZUyCXbry7CjfeLd/r/UNaS8NR+lk0kKwz6Lb5IT58H8bmnrlFZGi4jBuata
mywM5p5xhMAsaxRGtl85/jpg5dPmo1Q9dXGVflsJoWUWKExFDqjf1JA9JY2bzdBtrCTnENqwez49
hAqtmnuYkj083P0N0dHTW3rEAUcp8yjt7IfFSXQjZEihAmHY6BVwYJgs/XdtiJdE+p3jKae8H7tT
Jny9d9Vy2rUjEMgaaE58Y5hK6aY0uy53Iv1e8Ap5UAFoMmUmtPA4+q6Gs885/BWRdNLHO5SAqlE7
N/Xbm3nQ/Ci+C0dwl6S6OvA2UzZfGFLvtoOVJY92bL32w/gM1rPk7uNbqmbTYfTKo2AktzEp6Hs4
Ebv+/MGUDGHPArdXdiFdfagQu0D93DzfPXlJq2tmGO4EjDup+mnltbpEemeZ8+svQg4XqGL0z7Eu
JSKXU6yBjhYU+MmjJ9WB5hPHz2n9kdHOzK2UzE9DFjh5vvFw2k7dxgN2Wq8m2P6zOK1lCCY/VCDZ
BrWZBtYLcABpK8JdNJHr5pF/gWfInT6gkqGWNb9+CqxQKRcBYrn/P38eUJOBfWbdsVF5tKI+rA0h
dmuf0rLUBcTXTlOmOqQY4OVaapLCBBIGg8COw8dyina3bJ4mXPHmxtMa03MkgcXgaB38FC3qlm7v
soDqMEi3DNJP81Bc8oQYX3ulwdNF6Gvi9jen/Vbk1PUQYTpkE9B0cUOYGfqTATugYCb09+k1ed6l
lpDTTaNos6+XrCLaVERPPoGS+4b3B3RfTiXFR1R6HVsQi0NcvFevH4Qmr6j8eyb7zMi5FQ5vGRST
sg0QhiJVPxxq+ORrxtq7WD12IQY7z32hTlASdrvioZkS/sGxurzn+/knEbLRu834WvTQ68cP5S+j
g+ZvNhoziAyvCrYQdZ9w8ds4vEibwrXlxRnhhyN9e69gfynFRSua6DBZrbgzlAMpmiJEV2myAxWv
Hxs03ZH0IQUkNJ1zr85sv3Jxc0xYtdwLHLmBVIaaKDSqr8x6XeSB3WOOdbuYFjIhFLLDvspO1rqF
lTtscK7iFxgB4FcuXa7SThZMlKnZRHdb4jhrSYZ8Wgd4WZ5Y2N4hdH3+dcJXcARjDL7qLc8bLPF1
wYiiVakAkG+07N8fpe54+Zbob4sWcQvF3OCkJfk4vY8Fy7hNG5yLPAkCTtYfHhXubMHeKe5rs5zY
CaUYsSfe+WjGrOsEQihHYVrygVEP2G+X9xbopDcuirys4dTMqxDcX4SN/T/nzyc9ZF5f+eATPR/y
y1Xc2w61l3O7KB3SDbBCsA7fxgXLT4HmXt6chCfW0331nPytLpvivkB406zx7it5Kb6mmgvcWry+
W/JOtQqbcBq7FhAlE3oOqCl4v97wOAWCij4COIXZzNTH4RC9MSULDuI4G5oFdcyb8JTEMScr427w
o48gBV6s7ykeKpN8rG7oMulSOyo8/t2NQpC6s+IC9wRtz54pOYPlN1XklKGK9bi/c9tXBFXikhs0
rJCqVj4MocpO9tnU6HaelSgeVxlb1ka3JhnQ8saiu+p2fTMV3fspiPkk4pDeV4oMPH12aD785Ovk
qA9znX04NSH15k9gEStz9phpZHSdCaNy1pOWHdPbpd215xqfrxVKjw4Gtky5YQTY4P0LEs0DKEZX
I1UoYYDCiiMBXGICg2oeJJJGeDpOE6VA0H1yJJo05rnf3hL/2bdDd0O2iO7McEjrxvT4/mqZXNKv
1gM7BQkyum6hmCbnGPPVIqH5XfrTPkKCjJ9IYf6Pp6FqnW2hVv7imUWkM7+oQTNlDk9NJTliZacL
YwH5p/L0Rax6M+zjgaxLoHoBgIKqMFOHiGbfUnWhToAM3N6FdqmhEgoEnvS6lhin+Kkt1pGNsQCQ
+CZ0b+XfZtyKAKvojHNSijv+wRUi0UgQeH8exbUdY5eOqINBgZu3dTreKqnfiT24X9iLLmWftjqR
6r65MNQlcUuiEcwmjvFDFzgPK5z2br7EK9BuXf8607BSw5Zzg1RNcc62WpmD6l7UFuOicLnAmOqI
eM6s32PHPqaYzYyX+LpyB5hP9JtoapLl0Z96BRhXVZcesKwASbEYEhRd+zkyAwuY9AVP29yn/xNg
Zje3vZCwfp57BV74/64MfxjuOXDrOMn+wjgjesKgRt3jseshPUWOpNP2RTWAaR4QFvlbi1OUPitN
bpdyjhr4sRqUhAGRhomMDCJALEuhlsE4NypEO0d3g1zMwf+GttZRr48ZDxlwmaCnbdq9Dzcg9ggX
OfCu9rl6CED95d140DApor7yuaVd6bT1d91xYikXDtNNQwbxjGDCh8Q5tfF/lfdmJJwfPm+Di0kA
zXehaVxKNyGqoSnZeJ8l/0bZcD7njhGtSweQNKrE/5eAWrWRBLF9lmwAlsfMnvqLkHOzca6SN0jq
S01DVFLa2KJLLQFsVp3LrFyB7Limx4q6BASEJkPbgnexwehN7mDJxsRu0ytRpWoZwtAyQ5bC6dKq
957hIHEhChuTW1QK2dEy5NpYG7EeKkrngYoSkzg0BgFiGZfpmjdbcypExB9rAOzduY3Y7ZerxKrX
6P4gU894VZyr73lCzww7JZN44lX2Net2PMGYoZT/wrN68gdIBx1BlOvyJnwWoO/S1xdnSx2OzVmg
tObwZKbUXoK1yh/q+8VbgmXbEW2yzq0GnWklQR3bPr0bXFqfvCavWJDVGQi1uf/oiq+oh+JkhyZC
FirWQ65UPhIzuDxFAYT8OND72WoOldi5fES9hxhm19+TdGD5IUPIcgJmvzXchjSZM204mosCtXcA
l56w/e1QJ5z7AM0i3w4Dxy02BC2QRJRtk4eSgFSVU/iMf2LWJPz1t/G7xRcmCJRoYlebxE67fVel
+JcJ44w2CKFk5AJH7u0abRMHc3fSCcq5WdgdsRJYRNZ2aA2D/gkmoc5bBXwA5yWxftKUF2aW5iEX
EU8wjv/DQrR5iCQUrqKW/XpvFj/54YlCwgB4t60Il/RoULryGO9zs/+oxeic4Ipg9A5INA5A75RE
VPBLILy5CiWOe3kQX9UCH8c2ASgDIXg8t69B+oEVqPIvD2XOs/u6jJs6srqzt/Ptls6cZCynK2J7
9kHmdBEbAYa+HWwc1O+zmNZWzrryuQvicwjpG2tgkDCRtL7Q5nCcBxm1vDzFo7yueP+T/1fJbFzA
iuPuv8Djerdf7NTecrV92BXSICMBRutiXSbZhH3/8ZOg04MgSegK/MsBHjPOugNizbsitYA79StC
P/mwolThvQ+qHT3o9hYVhdd/kOVgFei5oI/4THY8qdI2YqueAksIY6TXCBiuBYmtuScw/BpuCtOC
krAvC4dMX3y/pdsCeiGiNjVttIPQd2wwfH6NLOXy8p7yTQ585U1vt0SvTxgfquFZ2eF5cAfCeY3f
/Di7IfmdNTWBn0JDFwApIHEoggVvZTGyJ0TZaMFPtRYIbuQX1ueTS82+NsZt7GuBy8iLYEsTsVvC
PBS1dEGusxfTFTdYClbYGoACM6w57KOse9EOWTWcBxzyGhdgvIsnN4sYONs2aLnrnyIfAWMoBWHu
wjqQ/6/qWCYuGE5jQ7jaXQ4pzENklHl8yO7ScJkmAvOCfB+z+WvcMevufD7gYf8e/MwPisRgBIKB
oKuEC4jiRmIVymzYNfYbEMCMN8nkq75/KIoj45y3ZjjaiK1SIjjNlv8vJg6Ev+aLFlMDhUIdT895
lZqbVmFnelVdkJolPYwjNDy+hVna/nMg9xtZUjddOjmgeEY3WeU9BYqBO4+H+omDovKp1clewUrs
TXArGNXEPIdXr2eSKSx8Q33xagZoO0/uOhKDA3mk+7F6p2ZRkNo4gvoCp/a5psU1AgbEPU/naiGr
gDpF6IzTkc+Knte7BBiB2bn0EqfKLWqc2p4vCFmhS41hgbtYw8g27RRkN+KvAHUlOU9ffi7NTrUC
6edceYf6zp3NHlO4Ee75t0+yb/MZSD8d13VX54fmyOEKSwAZSs+dc6wmnOnt+QO+mnaZ7HHbda26
coDXowEjqpYuCtdQEdZ+etjHU49E+7aX/GCPgdHApHHV7qTE06k4PmsIOj/F7QY1DpFhRDTjAfja
PjltzFjZs40g/am64hdBHvm5ayi9fjFmPKplORlAKgbYyRZkisVVpZn/Q2HdLtuusawQVXTXfsUO
yUorIA3ji9ylB9dFMHjW5Nghn+lXmti078bPCKtO2+B2z9+grB7pE7sOL79zLcP0CsRHws6RSEOy
3NAiVOKgOEIygTfxx/RfOMwluSjUlkEigzJlKumRsToYwoyMuGECJdUkWcVEJHVwZawW8/aHCQqP
riiMgi6SW7dfRkzpuVY+5HAxPu2Ic6Kx0hdmY6VrApSFUNszzKcr/iF0g95V/lrPGO38d0wangXD
B43exmQ2f+7+CnkqrcoK7uR3gjutINLySzbV0L7cf4ToAEf5O44BR64T+ORTmjClyK4MRSlkfFPE
02E8hSlrTD3OjbJWl3gfsHawQZHyu86T8GBv7uulSz/UNFY6UxsOB0gEyMeyh1PTSz0osGOO6lCy
2tTUYyyfuaLVn1WlRXlqxPiEYB+gprHWJxXwK3AeC9W0dOXzeBJBcPq+wjnQoUS1Hv94NzZa74mU
mfLs2quWwE234PAesKdqLs9IIyponJIpKfto2KDXZuvhusEIG7XwHljT+rwD3qC0442JODgIIpEv
cXUDDbyQQc8m6BFU08LHIKVqBxjYeZczLlWToFmGRac3FirFxulhou8GWHamhqb/bGHYEb6QDo6B
qVYBLwk9XZNyoLnJIsmwctUbgpZxyau8917uEogvDTEnl5DmoWRIPuE/e7FpH+OmD6AaTf2/BXk+
Ko0hRzY6d89EzBPMsox/jkqNstm50O81bZGwOn4B8e5ZX0yJ3fFf1lyVNGIFf+mlMuwycQnPAgI2
Vz+lVDe35DSjc05EKN5AsPatHt6AJd8+hjY/KNu8WXsNPCTT64B55bO6yVL8yxIiHJj6rkgAlOOf
wEreG+JrPbO9JZdJvCo3E3kENK3JaBhCeSOvn7xolPPLGfFjk8185FIWrdMJl0oSZ6yPCHYCiYav
Z7GBJCu1o3RNTUeRQiotNxj6zkxeyL7LoEc07+tShWUFSTHwfJHjQikuxKYU7WfAmkgE91T6MBak
Vn8oyzx0zMj3JzncpYhk3LlFKTFv7PSfdcS4E7bT5VFmgzzO0y1qovjW9A+gmoCDpxSNz7o/xxLL
HbuN/2KugiBkMfHlGwfpRW9n728pYSPPkIQ10DfmGQ2lvMtXoKLfjv2qMIYuXw5PzXd+YChkBRCU
8eeqscVKAsdXIc9noymgdkBg0/kKgB8q4QpYh5xQIpQSUbEK1AWdsqcwzHVhGrPbJOBxySzIEnyt
pjUA7TUcI8dEwWtKLC7aL9h+NpfU9l2bTTW5yRqvOlxhXACak/ceusn9F3CSnTK3K9Nzq+3gAPOk
08blvMGnck0YgKXYyU4TWyf/+IDauQoZ+GNGfjIPMlt8IXlI3Qu1s1TVro1illl+AjCEbuxLoZdX
g9E/O/8HK+ahEJL7id1jkTC4ishOukOidDm6tjJhgCy7xUUH1FTbybTPf7TZHZV7Gn4rRsDGqtvo
b+JyI+dhGyYmJvv2atTSaY24xdDnaVaDANfJgTfsKEBHlKO8Azv9Ts0EL0Z148A1Aj7ey+AP+YXw
Yeo7jngnoNdSOWTm4+N98H6xXDMx+QjX3k59QkUGReGVdXRtySe1CpGQ96wm3AKn1LcFmt33Byys
4MSdnmqFAKBltIDMiUK2sMijwUT2Oj47tul76SK3twBCq8SqJWJFtU1jg5amJW0QAjo/beh4M8ge
CTEfi1mET7VfVmanKXEsSV94r9cE0KQQQJP+u/nLp6io47Lvnz6+4Xqbwa1UDGX9hbBA3UEcIVw3
MzKHgidzloDwk6RGQfpAOtUfuq0r9NOTseEZAyqMDGStDKrTUMh62nXbGpOyWfMxDRC3VjqSbMAV
3go8UBXeVigrPk8InDiSOSFBoFjz/yHFCdwRaXySxrBlBZ8SxTyT/KbEuxwQ8svKIM7eMhAoJj2b
QMpxSwWwi+gz4ypZtgpqPLcDXMVs/PQiK2zWbEmBnnYVF+4BJHsfIV0H5NS1vKeGZx7T+Qzicugk
7siXw0k94o8Pwbc20+lslIIvjzWxe66nRFtfxoVyYnrtEW7htlbWTzyBH2wzo/6FhIAjm369BUav
e9g0lCSUp0cHgepgUcnupQPkyQznS0smFlVEIxszzqM/mK+fu3JY4ay86HWPSLOtBzTzYUO8Q7At
8XiMEr16oAjfOq++PFJrKA10O2YuDB3HmUXRL/5yFfGRaaOredTpUnbX0E2S048YpPSbjG0oe4kn
y/8xfjbOqznn1TEnGscZdGG3W7kHJY0aXlZthQvgpnGNMN9sRIkasm06RKHn2/oG+KuXi9ky9DPE
twtYMscdAvfTs96pvp47KTXvT/AzZojpYQlF/iaDlFLyU0ABp0aqbbVNZuT+c/yGAeh+lidbZ8UM
Rg0ToXs5bHnMPzWAJ3dm+tdEYTDT0B7ZPf8hsdSwRwxziJEGkRzNWc5oaKGS4XHwFtiQUtp2poKK
RUIKNHuh7VbLJ2C/mi8oHb9b0bJO/5XUZue5en27LbxwXDfot/AbrHiKx5ZA9ubs4P+G9S3sXWY5
pGJFYf527rlbBOnIjbaPav6YkvDZWEIZfjeluUK8+Ve5bxBHfISxzfhEba9IFpjpdE5mNh3YEl8V
DKjP8pi3Rjyxg5T0BeqonvTL9yFVfvdYhSXjcVZUOZjfjFeqFfov//ZWfosNvOGbbZPJROxXbjbr
jxFJGYQdviMVie6em0v2FmSHXtvlZ/IngiS/0unodolk4vqzi96cET2akO+pwS+A9dVbzud8f/Vs
13m51+kcHBea1TbQ5jYNCny5w1n+A/e/dLotCaVhTQaBy1QNfWVR3H7mGz06nRPRfVz4Umhv6FtB
VKjCcs7xSTQWxtSVDcycHX9u4Cf7QJHAP1FsIZmF1esEM9K6pij2tcYbCKN6drOKS/8TmnC3Nk1o
ebIx6/pfOwD5v2PGxTNu2dKPg46MbAQqjE8jFMpIpoBsNiqTYfjNLJltY8PYdRX0xPUMjbLAS9h5
huI0bEAVJUoUvYUeYT0lRL4rINkGmFdMd3hpAeeg7KjJscWl7VXYqleHb9UJQreDWV7Riab2mTTG
1r43jFLZDxVxfc5rPqZBndpJSfQ6z9Rl7NoMjhSLa3acVnBEUGZYJbjJI49hjh8iIZwTHmMmBFFm
3k5odTKK3QNttN8d2cSrLfTYhgX5MqUdw/WcUQ5gwUTzSgO3y3c9K89MxbO6LXDKmPE8IvblhNK9
YJU/T8vkkHo67JZl9nnrCIZf2BTjEzQcbXidg9OqGIudfidNT7mSQswcdbL8fSL90r5nhK7us1pv
tGZ9xgygBroA4BEX+p5l2Kr+AHPAA0STxN5ghqb+A5LMSPDmgednDwXy/hNX1Dy75XyIiD1kKAll
6FwV/s5tESNZ3LhcEiAqSJth5R3qE5o2Y7bso21dLrW/bNxOTI9zGEBdYENqx5Eh59s9jJjd/tvA
CjMufoDqq1gpmiuWoQp7ZzwGkj2ccXoWYnKv1/LHNWAWAk50d8iNBfvFllYT8lmu6V4zBMjuG5Lh
G/pAbiLTF3FeB+EsR9qHczrQCZGHVOxl2TDfrUoaE00c6UEiXAOCFSY8H7iDy8HDyICXqCo5P1Mz
61c7Oglgnp5IArivmJHJV/iWRCthKNoPXYqOUjqO1Pu/j4GdVTCPvZgbtiTJhGb1sWcvaGc873if
CijaZti2gt2ZtWVl2KwvzcXUAyGJ/g69AYdTgcks7XWewu6h+1lV+pCARa+Z3YDNtjfB49KJiKbc
BQVa3Mj1uJ9lcLd7Mzx9z1b5jNFo1uI7kXgVIMgAE2XcrPT3Ng+eTDa5hBYiWAIFPxoq8GqlXeu+
s5Jsr0fvQnSrM/yzfMp32Qs8c0xt08r+WOWnJrX8SHKTey6tkg6K7SHtLm6X5V7GtejPRRV5t2Dn
2FjxTW8NOf8Z/Cs19VWeGEBEo+MneH3WMwXR4eamcpffjAmsH7KURnwsRPwqqbRIAPn/UABRz73U
KN0MVQfegw46gkJPo4wDBtoZUH8i1OCemeKUD4d2ZuyDl6zVojmmq2KfwOzjM+VLBQ6r0a9PRyxu
8nD12Ro7RrRcD4G0Oq1x4Hf4TogI01YyQkYYXu5aLalxZR+ym7HYieelp9Mp8GxG6tER2hrdf0NG
Fo1CWesZoBVPaY4wIsKxFrIY70jgWDgqbGCLSwDUSxFTyFo/I1zDx3RqvK/u1nKTifRmaTbR0jnW
jULCLQKMVDyNfgnAYfIun64TqnQeXIC8YFRN4Wj06VAf3IQcym5nWlEAU9WzqQeHX/DXIe/PRD/P
N9zDDBJzmGGVG4LcI9LNqPzxsReBFgmBX7kJ7M0aqXZCr2bnVneX6M3h01JNLobJC2GwVwb6SKub
jwreGmS/nWtnYnSB2t+pnRp28igk9xPoo3Ww8W3HfOEctu2D4UkReni89SvGiw6nPFPiCb4VyY+a
CvPNUSyg5zFQsTM3tJ81G9OK+lkxvc9ClfPXW1FuUHQ36RF+oYyOJxnHuHub4nCj/69pfP24R/r1
62vdB/0K1VyZVTad1EJsY09ha7NRl2g5Aq7Lz4zSM6bO3E1iYVd+2WXqJ0HjNCh0zbcC+RL7XqoJ
PkARF4D/m4e72BxprCdCZoA4A++bYM7luoUT7OWnmWtWt6Tn1PEqkRJ2G7cH5uHaDf7/KERQNolg
E7XlPBVo1F/ko/oIUYzq7qz4eHeKtLGyxR+cEqaFfRULI+NEaU2EWF+oP5I3avXuAO4ZWCta3KX9
EE8Bm0HuSVsmMpANGwRQKUPGp8CdTQysMCPUVytjnJmsFV3i1psc31xdqinfD5FoSSK3Jv8TKXsa
+MSvJWl4FthVce4qOueC8nvpXqVWBZAiZerjPKaCadTodj7HVdzdnoxs1BngsC7AaDcocJqOMHhj
ONfUwVqS6NBxB/bU5AacoYGjHpR3tCXGgpMJCnE2VG3nvWV8DCt5t/aOQZwlwXBaPXCFCRiEv/iz
ubnNcqBqIWTPUZBSrWjjtjRjuZtIeh8G6tkbcF6Is0Kt/Qvl4nyLABSWbyrIkrxRAP5Tp0l3ThYN
+oNAN2fozn1gwD5opUME2AoVsvfQfQJVoMJCofr784nnmZNtsCe1OG8Yg9vyRaCgCbi+pn/Mir0C
QzcGmCwKfZcwlcjN/cWvGidoTVqXmemZQQiKZk14SYQm2NA5ksZNwWojscp0cwepW7T5QSCrJa8E
I/OHhFqwUt3vX66trzp2ivr4wQDD3PM+eHP8b5YXYXlrIiDlP/ZEHxYgSF/CTdZN+1wHha0A5zmz
WeuXFGQAzJLTGFYf6tD1yu+5xH9B76s4DV//V++AbvrW1jjwSeGzEP2pTGbap6O3Sijb4GkkUfPk
6pDBp41simVxB22AksVW+Ppwqh6UWqXvM7ZtcAB+q0Jj4DaeA3Z0kXGFjugwN25olF9YDGafdU82
s+mzhYyFhzeko+ywBaJ8fV/1tN+f1ek3LbZCn7qruABmqIBnr4Kj3JtkoJflSmI9EkKzo7x8CZd2
OO1pMP4SP+hZLqJmOCaZwSjBeS2USYXGVzWHePD6aWYuHPlFU6Bb5+exkiO4tCNyxRbhWzD32DP7
I7pb14lO0/ZDscnpvo/m1ESxGMRgsKpJDIwP/dSEoFCLdeRrhkYVWuNxsQcBpOzkWKMrZwdoiAtm
+EmT0z8P7++KSOtHC7aTJdPNBD5jq3rUhSXX22746Tykecsw7s68kEDAkOAlqYaqEW9u9isnRoGl
XOsOGnVR3KpwE9V8y5lbk01n2oEP78+Xq4V/H0EFBYdyTJc+hyejL6x11Y1UCg1nqz6MZ+W2qBpD
US92R+jjolRMYchVUmgM1TxYIuG9DnSKDjX8kFMobbxjVLpHWVBkUbeKRNhxw+TBuMGdISKkV1SL
em4LxuyUtQZEYW4PFlDrXfPYvnunLRPCywchSI2wlimp/RnrWptyradurHEFWzUSAT0eXytPGFBP
mnDZow/T84W88+ZqiTvciadked0b7+lNgUzERJNdJwG3TZHsWaa6fZHVQzg2Py5kkhR4QbXkkZE4
TqNxK6kXK4cKQ5klDdW++ZA0e9nhk6fm1ENX7T7GIVgfYYBq7mgs1mRKqMVZ8UNfiKhTBZmwItP4
/+YBVbJtBtYsCnnpVBAndi120hon/ZumNbrsp57/uzIYdMbYZqGPLHP4Se5r5BUlh0v3/0O2DLsG
Uyo10F7jUBtuq2plP3XJ88zuhUPzzlwyreF49xletSP0myX0PANP5eDR5uncAmUGpPJxruP4ar75
CXqo5p1Dxv1k53cr+eEsDFb8fDCltq0BNC4FMtip9SYIF49WcfzyQHijRQazNfI9U0BmH9EyxKn1
mZjzJGrjLM7ILVcwUSN6r8F8k55KM/oJQNyr2H45Hw5DnTwh4MWYiHOgnyzPydU5VuT+xK+ECsAf
64b3q/JKERzz1MEn3U/MlG9QPR8gxbuehx/J1P6YNOye8ynMyCrtcJpB/E0zsq3gnXCBIY+Dcerq
fsEt9veaH6GgyM0lyCHB86r1sr50oEyMLy0IQ7wj/flWyOZkg5ePuEAfOsLukIxlFddbHAW7NzF6
2rVvNchL1hNJQEermanU7HEdgczLig8NOhDHgIFscGLN+BStP2Dq1kDe6K/FbLswJ3ciCZa+Fz9a
E5JCVx5xxuumuUYqfJIj1psKWLIKJK+qlkIatNLJLtFh0nECvPkQKtiEjfnSRA7ror4w05rVepT6
EMJ4plzExp5lxDHPgjjmCWZTQJfUBxCntAIvyn26LPAHuI482ogrGX1CRdset6c2xJU5VuOG3ihL
9F4wyjGo/o6UY20lCRA7Av9pVZX7qTEVMuNIMTagndbAGLrbc1QOmsSCysSvEFpvAfFIWqvxr7Eg
vje9bDDh1WN9ORApR6hUyNamAW4PPQFLLAePD4hLRAkbgkYeHOrKxc/K9sLTD0BncE179MLbB7Ym
8KiI81JXM7x72E6n/k18bC0MJtOLeM+IDhBodNWm6MQJBWYlcRoUR7H8/Z7O5FqZhrHyP8jsJS77
QG9TZSbDUVlKude903TwsrRi6rajKlWwyzwrlMXJXWr+7tJ0CVrl9u45PNDab20uXQfYCVOCSZ/t
EMiiY8sp2xbOSrK1MGYSHN+ekEUtSu8n+tq7hIpiv+JO4YgunneahbEW4vaSF7kmgu6W5Pn5YXij
3zwNtAFWIC3GGuZtZiNw4Vzb3U59fZT6rLq3G0zYBrS53uRTT5kmBTp0yAtH+1JG9EzMjEbMunDI
2x4mr6Hxhh2SejKY0obHMBFrB5vf0krQr5K0itsWVZYIiZ4aRf2mqg35Jd2gGmYuc+osdReMHHvA
t3BcSLH66tWjwRDJ/ESqhKMJGp7WmEuor4x6kcYrbsdhxMozHMqAjxJzmIBYge1J0MFdR6a3JGmi
Xj4+KnqOG3E1kTf4ybQV8X1j3JdZdt5/weIJaNyNu5XBaz6NkIo3KC2Drob1iHV3KZbojJZJV2dq
0t66j4uZrD76RvjHHt5Lb+3GOaMqhpT/91yQsW1GwvLVqsEUnxQdQ3RXHDk4ewFX9YfkANtGVIkH
m6xEYMUiVxnGdpxHDYm70vsVA0t0jza6hgICvBH9PuIN/8+lLjXgutcqInPFOOuK5FGhpDFUH2mA
gxq6GX7luNRKLwicBkHNFZZi87EsBni53EPOxPZC86UuQfaEKZIug5P3qwVASVyvxzbpXAkIKmJt
ulD/+vXMVieUkNDX0lN15OEMN9kiksAWSeOc8HY3kffO7HkVKDc25dlm7mJCCyFFaCqD2VhxirmL
j2jeFz+LM/Rfc6jI0XE9r1Jezjgm9T46UVUk03nW0M16Y1SW6WEYV4ys0F+bnMpPOZtoMvGM5YxF
ftqHLVNZHgR/cEPpwZfWGNhLRme/QvlLGna+YT6zBsSCsGY60yZ2RYth52Cz+rtN36kTOdVnN6Zo
73l4GgLMmSEwm6zhx67jQSiQZAF8Ki3NTXizmNfpFlrV6G//VBDeyhO2ESftGqJicf8+prIN9odr
JALziLWKEXZ2kyUfRFnEuWnmciMQQwsnXkzprFKEqMz1L4oMCryg/qK5GCrzkI4GTwsWTVG4nsqa
Ak3/9WOxmH80UHu3f0d2vrXy57+sut5IeT3jlgDxkSrggFAEXe0FFMXj7Lqd85QEydcChBNE9f1J
sIv1r/755HK2pluwvNBjv5pUtUCEugRpNfe92arxUTWFJR/IrHKKlcTp5sZa8aO5obIdSxC34xkf
O+vFFhpdBghMfuOjcwfIo/i/Nv7RSx6yPY85/7/uGlEiLZ6vjmECxq5NX6SmkmUO5obPYI5vpAbL
YwK5MrPgQQP2QxtA3/LXnfr0+vuLnqZT18LTv3VQc1GOpQnL9rv0nPRkEri/4La95ZAnObIucc7I
Ze4oprIGb/+DnwR5TII8TAzrKrulz/Y5cmnx5qnc4QwamibF0+4GtnzVyroFBeBivoxL27lrqZEC
CMQiL9PlyV47rzk90YIvkDvifs23vrV0sFClXLVUXS5ynYFzojTBuWO/LsSDCL8CSE2a9iDO1g4M
BQQAwx8qc4BAtJofafE6t/MtOJQOzT/OArCqGeZ0130Wlnfw8bqFzP01kw8LqyxgDJe7MWZWpwXU
nOCOQBn/b0HOWMfcSBw++aRcgg/jtOFS/kfJvtvwjQBaiBYCNzjTN70bEGPhZlHkhqam9sxhc6Zp
glfnC6Q32ihYxG0UUDBBVkjFoVhBoqIrjgwbNaKlQffvDxFkWrMmmc8o9H4UVSOzrjNXcveSlVCh
JiRKswlSBf5mqhYhnqUCftLyKeIXoD+sAzgv5++0fz6nzpchIJL9zPNq0DXLpobyBkDCvEsVOitv
kYjSeL1OH1RPYW0bsoTWPEMBKIfXnmsjNoYDdxjXa61go3iz6eqnMg+OE0dvCliQksrOzc4z7Kp6
rQEYP79SZ8nG/Hav3KIJ9vKCzYM0Gq51OIdZg+EZOo6aV20B1mEUqJVypq5gHlje7UtZfJNgLCqX
8NtnLyA9UEM69sqMN4sZxBP6MCdw4WmI+jnGP1TXGFfxHbg+gH14fwnu6MYw4bmfY6FIODMyuWIX
qsqAla9eo30jxcs0XRkxMUdXkokKE/wBHsOgcNCNMSo+El+sjrKzp+jd+3786DdYfa3t2lM+KcdK
/PPA3HZahlct/KvRxDkhCj+0yIV4TER+6MPIZXIhQUy4oNc3+L74y24x3Wf60aX4LicQ+EzpgbbZ
Y3sW96opDw9Y9jZclLndkj/ejCCFaUUKP240JFj8cZu6DMuP3HzpmVoCB6/nVLpN0U9hq+E18TIp
Qrsku3qI3Kk1AOl90KT8ybILvq2Zk7ZGJUXMz0gqhYEVn+4FW0kcitoagXOgGv+oZB1hhmG7K+re
N5JottYIubOq4JKyIeQzSeJYDIyASCSB4OMixzcWpoRp7VZPP5MYfN5PTo3xoC6h1vue88fA9KbU
Bwdicx5C51OwLATZfBxQPcYjOgEVXC+eMgJAW1WhhCa6Y1JVImFNWvTR6dSST5YAd1m7PJNHlyt+
XEf3PGmHT/pBdKYszhuFM0gs91i+F95rHJUxxXo+9SkyUR188j2nWa92qSodDf7jB1vCQYT6/G88
9RiKajLTUZj3+Jv+Fi6jWICvgVdC873kjlnGRhiX/rOkeNHFEi0hZi5ln6ivfYmj1wwuF9SdVW9k
PSZ//2SO6v3bfpHbF7nM2X/ISmiddVCec+QyLQxKmBsd1wU+OgGesNZTdC3eI9oBZpTod48UWZVS
skLJj/zHky4j+s2tEkfyH2Q75udDeZNxdp9bVRKjf+0OYhmSDCttnpx659PTW8SEhqxs6noLHSfR
OmulvHqupxxEXk8CqSUyLgZoVBrV/dGlfpOlFqtLn3McFbLiJsFFBky9bNlGc4hTxYrZ/g9nmxw3
kzTp/MGgLK7XmjAqWUM5i0eGP85jtRpMII+7Q9MWipVbWa9V5KfBjP/UszGsHI3NHfgcKo8UXDZp
fzDbrhAWW1BezjfX6n+GDOfxlCnM85JmO5EnkYHqoOclG+CttTSKCWD+GqRCegniLTlLpzFcLwTa
N7CH/BNKVlWGDvpgnwiqhF44SzK2MuONc4PEc+ioGzi7vJc1cVqhZqPdtT4JRvFssZUG83fPHrpR
4RRSOC9D+vsDVnG6b+StH2bReyUjQDqmsqj1IethqI9IlbqHrVtZYHwNnWkcKmaXcEiuM11YixE2
7f/XVUMSoKPzFfdQ66M64+CNJFkfvmLO6mLC8bHklkh37OpDf8F/nULb2A4hsOgsXIjSEaWuoAJt
Duly2jmV2t2Aw5/A7izJf3KcOSZh5txo29Bo4GwhudLdBbdAv/tI9ZzW3/AelQkakda+ILZk4Rl8
y/g1kcWgh/a6gslVhm4PMTscwKf7Mvq9aiGpjZZ6oA8V80hFr+WDtEdvPYVD6MCopfQoZbS4YvE3
XrSUkTWYZleOFDkOTOTltENRe/t3qEYc1+IG0k+mNYBSdkvJkQOb9TuP3k1YRsVR9XEYcCoT0QJZ
i4acASVgEGDXZXx3eOJzgS2JFPX9yWRThts3X4aeB+rrEVT6BcLkN6Y8mN2/tkwiYily2s0MdXPJ
91ziWuQsAAhz+0WuNRGoMpySOJ0IFnrlpvgCcF3VZlxMhKtt9B5miJsn6fZcfQZzN5cpM+HJdruu
ezgxkfeXXmHgRCPUqbuRwJMeH9FeopjES++CFrH/Oeqj4h94uUcF+3kMgSJJlLi6g3+aEaC8NoLn
M7jFRkjhET4jvGAbgkRTe8KStYkf0vGoInjusG0FRVtVR56lA+KquGITLCvtd9GIfQd/k7tAIVGC
2pm7eloqBhK0eCv/tOHltc8rwqvMBIPqT4ho4ycz0X6c9xxCC8Jy8hLQeK7xg6SQUEGmlTAyhomN
KZybAltou4sIJPGQkY/JU+jvWSI+uHnnNQfsHDCfNkvCKaU0d2v96bdPSnHmnCXWBYCaVf9P+qe8
q/KMpcm3r5IzZs8P8D5XGLwHFeYPquMM+Qhov8BpWo66n6+bW047m/JiV7NTuvIebgdgvgYCdadn
OrD7Zgi0Ybq4DDzOF53i5sp2F/XNfbbQIM1J2ATPCaBBARpiZHlLu6oQ9UIgncRV4OavVhQnZOqr
IsmdvU8ekHRV7okrVPHJ+EjGahQsfMRTEb6l4jsfxkDV6Spi3BsE1UFljt0Za38xCUqwiMh5QDPB
huBLluWcpKZg9uEeyIGqd7s7NHTIPBhDNWsAMvJdnfPLnqMHvmttFUep1fUk4h70eCoy6f14VvCc
RygZKgpsNRgNi6funyRQRjUHOQeeOq8Zmve5/VnrzQqjbh3mDjBMvZ/1d2hfGlEYxrxSCGM1w10i
DKRNfvuZ+ZQ1V6If5XMYAAhfrWRnzGBHRnqAjGxlc8qlSpqA16790zQwwXQfUftgXED67T5CVhsJ
l1yAPZ6Ak11P/ZJ3oHm4Z07S78VZpeG7poIcnqyexsyuh62UwJ9vs1fVjzJNdNFD+qa0Ju1E6M4g
UQlJ2Ah9edbXqsbhO/H7Tok5qXlv2i/vj6t68d0hRzTkBLsYOG8ylPehxDp5o95TGyj3zQef55D2
vHrnV8LaOj0Afp3OZaKanEuiWVnkDNtJX9YVnTBBRtDLv2kMO9Lraj5+Og5J89IhWWwxNOTlo7gD
vQcu4qEqgAPr3FJiM2yq4AK9CvGqWZ4kQv/b8EvmMZbrdaezMR/TbWPQ4ZVulAxmCQSMfgtnOSid
ykcQ7pDCtyJ+FFyQnDT5mL+AdZ1B95hteMH5FFhY7qJJhmI3jzElG29+HfzVWiTCJCWtqrqafPve
eIhM2X5J+aX2vAn5zIRPXQHk6EDNQXeV2J8h2UxCsYfuIPOdR4Q4OcsnyRL9wUCZs+DF2l6fEk6Z
J+dW3dVlNnG/CNmUhzpZtTqTQ3Y/5w+ek7KkkiZ2SbZDF0IdrtISjioVx/Ej6Q+tFDVsYk0mrwTl
V9/6mYgUGMV8F6IQsjDkJrhGNX8wFBfqR0Td9xp97+X9HpF2xoYhQk11vAmfvtCEKMZru6Bi9f15
I7SZNvy4k8iNf3RhymL7Nc+TaB5u4CwofOblGDSPIQ3qSaXE5Dz7KAbwfXY4nBn/eK9Oxx0V113U
uPoRbxWPlLmFwkkb4Ynh9Hyb1gCiK0k3L0W33Nymtv++pD77cN6fHf6QkNVc7efaE/BKKZFcBpWX
3Owk7Ax6FoobrNBSH/FLeVFcveNTeQmaniO8FnLfc6xKKgboj7yonZ9zA6H85ZNKK+sPsjIDqWe5
6a4uI/+BW5CnyuECpfh1OQMmGc/JG/KHcJzOLGXjvE+pOHnwpB34chvcEDXMFaQhGD7KmQurQZnw
7lEomIgCwwd3g9NjH03VNPwxy8hsJM26MmnzvIdTxOAtDksPM89YhxAvMhgrL1TxM52r7/ucchA4
fXoJ+tnrZtQaAKi5NqLsttkz7SwA2qJb9c8zw75OjuO0wZFH1SwqJcc0yabtGriVD4Cfi+4WOW0Q
WWMHtUscZypi0x26SbSJKYoXb5XPhq9VbJ/QV1XqriKnMeUz2TUPz6vNTMYKYfroHVYhMNX3cFJl
aKfonRa+qDacNacVc7ypL6Jwn34q4cNck5foLKalem6Bhs4sfkJgu68IMJ+OlApNIPhpSH0geyfy
VHAf/lzkLuFaGD+RNirGsVX57l4S69s0Z4yuCKY69szYjSV8gw1gkXFwGenz0MmQu3fWF1Ev5Zfq
7IZLXhPYox9ZehEo09VwgHY01xB3rNDQLzjcMl3Fqd8Efvojm0oSEfBH1e2Iv0ET9eZMe6NYCwl6
/C9cUZpJYBhbGk18xgVp1y08Cq2TDtdEK8t4tmU5XT7/TMgaTdNwaws80KZWzltcDgSHOZiCclFi
W/xYsrJESBu/e61SgyIUaEkVTwcnI7LAMdeBScF+m2jX+0Bm6qa0WtmV5gL0qKyslI4tuAQaoNn2
TxUoB9UEYO2cLZanRG+upLFcwMRdwS6IsfhS4cPrPdpObKRhol31sDq5eDRS4einmBiKkzY5duG4
y8nsl/2aGNpx7j/qYFdvgnU20W0R1PIu0kuh0KXtfs6oaLtZnYbMZjeFxMmy1nJJ/J3xn/6Pu2P1
Jow1G4B38FUfO6gn2a0+bCzpSPtPSG8r4JvQNBnDLmUe9jnCXYdWzzchjJi0MgPX5tylvEZGXoUU
8X5c+iC5Ajz2sZWgOZDPbnVNzSQnZjis2PlwqR//rRdUZBQT/5ejeINuNjhbAfCgH41xD+AUl86U
tk0JFpDOXV0eKcLyyQXq6EUHymL8Z+gHr+e0CEcqMPNeXPCUMkcspSmxvEyK0uE5rgdyB9PnZfuD
Y9CE6TJkJBOfPx5vTwhvSl/zRJ6yoq+PxLMPjSNDGjQriMzwXNqeIRriTnjGIuHNz9hfPE0VODYq
rOArsOdsuNJLr38jEF1CpOdZkSeXJT4hvuIQFZvHdntc9zzBHvvALPQkn/q+kc26ZumlqxoUNIZQ
JqGT+nbyo9tMTyOe4VRec+0/qLJG2cM2gQpMvCcrZlxF0ygvbfaf4m0A4WcljgmQ4MUMy6TEj8xd
DLmzT3ql88zH4MdigO0bX1jqK/0gEKEQGdor1mbLQ7RanxnNeM+UCegHdtPXpiqa0/uz7BC03qHj
cG+pxzJKzvVEVBWw+H6KZB3Xqcrd0rJ4lfUfXGBSYQpdk2152RETBLkvkJ4VUc0ZCX5+XEaPePNX
JNyL1M3TD3GgllwJEEoOnO75Y/VFifMLU78HVtYh02bls86nvdAA98+aT1OAw342RxEU5egi/LXN
6Tq+sPOP0quchaW/4jGc1oWIlQD0obNljyTLZsrr9APqsTNWyxFuULekD6XpbqZKTrYGnBJpigBr
MtvnzQMANpn5u05/ZRK7pK852/5OXLn7gdm/rq57M4XLG4Z2DDYy4PeOUHuDrdG3IPPCH6zK70qD
bkaJYbwh1gKG3mCxh6tJ+KGqDIkJiaIHkav8ANTpsHu62TaA0UWn4jDsrRpDT0ebMl1I1R2nA6SX
YxoJqaTMMhbEUgQHAEOVYlpil5r/ZRrpaR7EcM13OKslYHPhk2RRxi0IC8iRiLFVBYXn8b1e8/97
bOknx8YdacgHlVrLq0+XeID52YXVFusEUmk6zUtbWpSaybpTlzPcz+Jk+PZs7+XM17qJunqN8svp
WfeGPQI/AjRdxtBazj0KigsYbbsTBRFLPpnO+G8Ms+6NIqZ2unpSzn3C3r1M/bFpOIZiRd8PfEOL
0HBreRYFsNsrWFy0uiDziZ/JFukgi3KOCDwjmd9FvnzBfvFFUrDUoi2bm7Xdj5MZmo8Zv02UyJ9R
TvD1Hdi2c3kpJx0yjr0AsTG8zXm0XzIcjJYzxDHO2FCrvJX8XNvyiIrAJ6W0d2n6s2yulPYPZE9z
h8VMYfmCO/5bYyjRB2ugoIor4oqw9I1lPBSmAFVIO5lbD/O9d3ZuAKhro9iAunnt5SZXx3KdwB/I
vXOU52DSLdfGooqKw+703kPNnNfc8g7/4/WdlnhY5jTELjFyV6v//qfwPVnRtqHJ3AeU2g+rRMpf
z6GknX7J4E2dMyWcAFN+8uG+/0TiX4UlSnGAVRZly7461EyIDSm27m+/A3ryZHSYrY/5W2IRmERY
5YB/ASQ2ZP+WfxjPNNC2OpWcrwPZlfM5IRMjF2AGgWMsmvte5FMYf7U+3SgEh6YEX7ygMc9tGfk2
YLqAA/H4BOACNaqH275QgyMpwL1zm+ZEcVNf8efBbo+e4k1pUES45As4fP+FO96DRZEQU2cKBHxu
jPGiB2up0GYYUTT4h1taGVDitCoXMgKBJmE6p4p9acj2AKDucAuwdAHu8n6xfzi2VOCNOWAzHVh7
NOCsPsSoRegdg4zpKfZU81PLZc2wQURCmICzLR4s0aGp2Z72YA/M9OGs8LZzly99Xt1Oe1w9tEvJ
rtx4m+uMChm9WzWfSwJ6bkrfhoWRUPkI6Wu3pyypR54C40m/NMyC+6YRDYbL9QAMQhzhdOToqp9i
3UFCkcHYNC9P+3Sqrn2xr9656PdvBE/xhLVWiPjoYFVxHgOhKl9pIZzPoDyglQL92AoatmKxobib
DlQaQoz5aQrFtBP4eCynoTIsQZoWaWLe4c9J4mCi8jTUUYm883PfKhA/0ZUWnrHRgPGnboxezvVS
ezxIcfrcMhbsvl0eUHPYTT+tUxJW4HVrx7o/QjI7T3g7BHGF/tBJfcV2D68Y3z5gU99NqB+AblP4
fNWea3/Bv+WLsFuMwq0wvjS4AobF916kVKpi5Kjh1ztCcHFn4ML4dIerPqX8/oztOCPY7En8hU3R
GHA9lZ+i64Nm3eSfr9vALF/FahGYiEiWwGJQv2hvaBw7Q2+sqHl8h5BHcL9Mgz14BhMDJ9yWYPqB
hI6oMo6YcaavXxFFr1vbRmCXkV1jhFOCjzgokvBPK5TN4YTv9QwxSVfeV6Kr+Ti7qQWc24u2VkCb
AeeaES2TJtkyoEJuEXkJpks/zvIRPAGTankz6uGcY3mQAqfm711Tc0fX+9qgqG75OXDn7DwDQj2m
De4NlD5dOZQXpqmfp+OgBUSinMAySp2BTZaYgZPgC4wYV4KOu3f0jo+6dD5qiH462cYIHAxzL/em
+uXVugaKRIpeYZ+Rdmfefm0BggeZ31qOK2BFRFlZrBXjii1F/7T7t/QIIKTUHctSDN7cF+/VzNwZ
IaYWl2NZIkVPg/30PMr/v3EzA5PaLRHA3oGxBxXK+mD6IcKs1a0S5j1byomxAKyzToMmWYb1W99r
BZ/nWSd6IEMOzkl/45DY+Y+Po+moUHOBAy8WftkTrsIRHLswjv3XrlIwPGF/qamQ0MRqX6dVB3i9
KtkM83iRcDuE/vU+esmdQBRQIcC07rOb8KSER/4rHoGLidTvjrEHW+Gb2C40SL5npeQjrh1OKFNs
iKwugsefgQlKqoiIAt9IlMrLqvsYmMD3kmp3SG4lCvHEDBhgCvCaX46xt8EdXLch2fcEpKC1zN/v
ebksUu4Humq07ozgR1ldoFGungPNK60uCjg8+4nNOFzZrPAAgLNR5QlFl5TDWyv05Z9VjeHBul+D
as+ogs1n54pFgWWpBVb5FTloqLXJo7FducPTeyWeWcajZlAyJyQ0t3MAopo0kkhoKeDDEXV937uf
kMvrHrTuJR23SAI/hWJUnZbXN6B5kfEsv1OfB2Abewt8P2GdG9Hz/Cfrq8GXq6YO/MsAj1xCbbU/
5PbSWHhEc14TWhurq3Q8g9S8D/uWDzw6daopLxT9wn8kjKYbYtGOCcl4TnB5x1apOFER+r4rNyal
wOzG+5rBD4DpRt6fKTlGNkr2PPumzlUTXfblM1E/C3bIka7ax0KON82XaB+C3+UuObLXjMBWztFX
b7B88a+54kLB8InUuRBC+PJ1iD7Qp4Q/H44TP4K7wKMisnHbGm07H51KwV3JrguZVk0vXQcprhjD
RtFbZ+SsyU+BUNRpWV7B1AIx+1RN/xZDE+7G3AJnvO5wFKcup0YeJVUEaqzOseqYANbGKe0UKYwZ
CPqVTcxCA8X8YPj/IXuR2k7RYKUUjIX0wVuZMLnYX8UjjKmjJO9OQmqSGsn2MJDvAISfIAdISy5I
cU6a16hUqwf9dr/exp1CA7HMiJpAsTMDW5F8o7XwlqON5b/PI278bIPUgwriG3gf+oY65OdS/sdA
OdS1tEbo4aYnxfovQ654viAPn130+5Rg95guPruRixTBegy9dZb+utXxN1nRNzcbPyKoykVMGXrg
8cxIB1mz1esI+8JVJbo13ENWyU2fGK7PMrukTazFVIjqq3HA6ASh4k6QryWxJ5XFguSv/t3zJf0U
4yl7Bd2wzut1/xRyxFqUFkasoXsc+pgf4aI9XgAYSy1VHGZ//Zh8dTusEgE8dVLHJ01BWtKlM9cn
6q+HGhchphbXZSUOBihoPOo/wzzwfml6n2pm6ub70mB8JhkZ3Tq9VVGqYMX0InRA1my48REw9uY2
UKSkLFlQJlfLSrlEVCP8EI9LRSoOfFqipD/2+ECv3OEyYMC3elaf+UbJMH5zXoUSobFHeOo3LocY
mcy+WelxUg1eA3+SVFu1MiP0qvAk9h2ISApA6TfcGeUyrnipFeZv/tcvtDMF61OE9D0MzfsCd9y3
lsT6bm2HpBXT20sIadqPXuhs6smn/WWMdcYQWnQnikBGN35aisQ0o8PDbYcpmX27BP4kUYfjAnpB
7dCofalMGikvP3fCQQl7gMM1Zq54OTy4cCgMxxHPTQ0iTDmsPS7TBCpV1AcRgv0IrFiN1vCDctJP
2zT0r/Cfff3xA2gwjeBFWNmet81ZriZMI3d3AECwUAt2Mv1umBmEASKooXK4nvTIw4Pv4gfpUsgG
5KGo/W3AAurUj4zp58zDdIjr0o0pECkpdc0bajG7/gpHZ3g0CPPDFLkQnvJ5f/Sd4X5K/f0NKq2b
7LUYUlIK+r5Pp48a/e7VJK0E/RztNTIHz3zf6zlGj1Ln9HBzGtcukr4NXJioLAlxnVrIJmXnM1yS
JSlHAjBA9M8/YolqLm2fOOmMHYFJCHFSfGBigDHpdFfc9AjoENGEbpMP6oobpwnuoJlBy+MpqMjn
4kyZbUEfT6ZlUcEEi/Wk9VAwNsVAwgJUVubQ/cag7HWgLUX6PRJ6HviWr7p02WqDSans1qeE8O3z
CtaQXwM9jAOTE0+rur5cCcAJkmDQCpIFzPKD5zsh+BHwaL0iviQcn2UCwrbfTtCfed8HvREfAjLF
JkKcUhnmltp8QzUtjukaN4ZR1ksGqHlp6M1nK0IIWH3SYcEx910Oc2KFiqF6lCUNyaKiqN8btQG/
VQnXM/Ja3aXHvobBTjGNsCsg3fRjYJIM36cnu0bh3ryOoHqYqOfdg6SvVdEmmA34eZF6FwxatMej
bRtr3ttRABxEtrt5b90nulcmeGVy+txXQUUEj9GgYtC8D0eXybbzGH2I/78aifC63JNxoH7NqHoR
Cr/dlnfPngIyUkcV/ZygSO0V30dlrR/sdAKqml1Egf8MoBbp9kCC6ETZQqRWIMrClitGo4X0E0zk
tacGP2GWJsS6cdYUMXZ+G+eZC0aUm/Zl9Wy+cIN7kAaNmzTKn0K/cvNGTT0eCoeTIUrZu1DZyAXw
s4IXWJXMuiuv3dmcTmvAO+u072kZh3pNgg5Ra81HkdzvT2bEONz0uSJjmF5aLVG7cfW9HBhM69Iq
olNDS9wmMaDC6dTW24ZezMx+1qEyQVJHNye+nuxw5tQdkLQ5b3O5SBQ6lQ9pVyPql8xBbcIAzT6K
GLVQ9gcUhkozVIr7PFJZS9Ffel1UUStEKvSl8/01I5nscyQLb1U6bVFjPhGEP/afY7Ha8gd3kDUM
9PUtpsZDNPhXiucmQq5+1iXEG77Bed5dhhWWCRVmesvvuFSoC8ffsJxuXyPZPWKMC+Gnx0BZm1mA
mPUsYgVeIPKaGE4Rm3bCDmrvfDjheVt0jnszbaQElfAdORtac3MzcZrFWtP1EnsvaSNqcbm4J8uz
ieUj2ONCbYMuUDOD1NRAgXFjrdieRW9RirErsdQPs+vMf/fP+fjPF3mSd76bNi38iFt+pcNAhFcr
H0FMuN7WKsgBgK0fp9SiA1x7+lpx9r1u5330SMMwzmjrj8cA+/kueyrQX/7wdNVyHPmOe2no4VLV
3p//xk8vMTPkvU2WikUxWgldIn7YXQ3X9ZiduJGtjc5lvNwrqkX977om0eSdWTzEFo3i9hydm96E
WiKN+kIw5sBxFTFuad/Nbwledcb+tpaFiG8RBLB0vs5Ad1wvwVtqRBEm1t7wPQl5lwZ3Sl67Gv+y
W+mHBOyzRJlqk+EEN+qKWcNLXPbbRKfJBD/IS7r/1nT9HqNo/7oGbRNt86ucLRI2brN0CnRIUKcQ
1NSVvRW5l0UkaZnmrPH7df0wlEbGAY2towsaLBsm39j+P7eaknMHcrRsIS8jKefjpa7xxQ+MnB1c
Nrnecd9XUpBKBuW3EbAVP7rFixDghdnVPQcR/CNJTzQH4fhmUmmqfJo6fZkPB7LXojGnrVdBht84
TOKKIZzfVn2Sn6KNdFdWDEDMSWMSVPLjykJt2BEz3eNbZalAJc1Rng277G4AEUfi+mzzgWbujX+T
tWqG3XzMMFOqTWpc6iwk/PaxMPsg764FdXMsSXHsZsN/2yZhwL5KZN6r1NnsMUpAbQbSWJFeIvKZ
Zk9xzS/3LMOyneSV5Nt08ZfGIXwFn/n2Ug9GEgvotxPp/qK3CzxuUjjJswgr44oHpAzvZWVK6699
31I43oTYDjBYXLEoJ2E7xiy4SS3wxgRohptxfcpp3avfbLh/k6wBZb8fpc6h4hB1qaaZMI5RXGDz
zUyIdy5Q3CK6FDaiuyl0sTxvFfiMV8fCGZUYQ0TSVKSlXZ+vTKVj0fOSNL2ZGX5TSZGp+9Np6dhg
zgA0oYjRLtSkpcJXenNUsMjZYgbeqUu5TgD/dC5rgYK4RsLbF9b/Lvdi5mrlaxSLNlWb5cxebhZp
kolOesOcjy1ZydxxVgGp8r885QF0AbH5K9MKL+GhpOMJSI/6ozWFdjdHMZjWMxFjGjaEw35m8+BK
8a0d6AjS9txVgZLXDaJTmQ4DYYh8oMlsiX855FxizphH9bpEI0Ddi2xGakdLBuWFXHDlSf6nsQHo
Si0uQ9U6wn+and0JiD2NrqLdh4Y9QQ7jHFTRNzLh4tN6VgRRySAjtYATgT2EZtVPahuXqkJWMKS8
jwr8qf+DeJ+Dfdz1MTVvQLTUJ8RlnF8SmUdTWi7zXUi17qSHAGWv2U8LpLsWDiD3SciweSwDB2Dl
fM1B5xzyhn5fdqB/kvhPwIbbqbw+ZyqoHI+Q+kU3G6MOiFAKmDUMzTvrDNxpABjgmlpo963hE/WN
icn3gYhb5EXpabhUx+mNsSucCnfwzUbHYANWZ60yxl1aH+X4u6w51FRJbcSFDVGAZVYu/oIhRjNL
q3XbLo1evqXuPT77cQxX1v7yLoUoLjLM7x8n+xUb6miEbRQLWGbP4zrKZga2RyJz4hvhDUI26led
wHaGohhmPlHW3LechitvtjCvH38NBNciy83/yQeCCICYZ/mpEpwHmSxergXhyol78WagM5wCdZik
IY84bCUJguNSWn+5aIE4ooG/GkORu3o8WtNbrpM/nt4HzZZbDXTwajEPxgfRqMc9MSOoT9nDLPuF
H3B6LLvTGdbx8lS7yoT5pLayp6gCc4WKvEKvGLAn7OtbxFBFD7T7KjDGJ2Nwl61SujGcw8sRg0j/
O+AZOp7b2dZytrKmBjgtxNbt9T4Y6Vry9icTGZDGQ6LkJ4aJMnZ84hFUQGUFzFE9wEwdnWF2elwy
JvPFAy+RpwLSM64cZTkmSkbOjRD/31kczrPCGbPY7WJndbbRaEzFClalEIP8k4T9GZdUt8qZJmkq
IFfUMLncD6YRQrbfBpMtKgIxKzAKW44MO2KWJdOZMhXmDmNKt2AyblSqNJmts0a0BeWAtZ4mYdzg
iXRMVNOjfiidOPMo4j8jB3uVAc/3TkxX9ezslz+Ptn9BDHgt2J1i3TktnZFsdHw0a1yMVO26JWiT
F+cyK6W5k/bABekmI0lhTsIQqvpljA/FytmtzhMuvGG8hxQFUq3351S7V5bJEPsB2dYm4dvzMtdw
mWsGy9CuLxMz0KV1d/swIGYgoT+u5qROncfPgj+rYhbc1GqRd+lpyR0hjWclMCZ9ZWcE6fqPF2TF
jfV8YxOTp/Auvy84aTqBSdHIFaiguRP5Z6V4tXoZVkiEoAqSJXEur3ue6pj4Nn4nZfQvQgBLDdpr
cXiIdSmCLnNe2exNTJZpcIqkvX2g2atCLTSvZ5BB9rWfarzYnBgfMA/X8EGGggcTwOuzLxs5yUqe
r2rNCwhV2CdZbBIKNVgZieVmgDG0NrmgY6p0/8v045XlnVD9ilam9zo6wH3Es40LGmhoqa9QlnLS
uUO1BdEeJOJ7HgohVd0uS9kakQYb9BOO4hN182/TnUkQHKiIGdvFHChcjA1Ny3LiHf0zLU4uxvGX
OYJD3zN76Wv1Eg0LTZZXerJodhpYsYFXjZ6OYn2Wxr/+ba9zJKahDVMmXrutqkqtVGeR6OuM3X95
FeAzLdKOQ3HuBUQ56jUvjQAp+U+R4ebPANLYNesw5h5JCMeHBWcF3riSy7xu/UvAEhBgInhMtqvZ
M7pWpssA+am4xJGZA++rAA7nHLs/p9Inu+FTZR/MmuAzysZMwyUeVr7cVfqpg0i9QcdkrkoRM8My
EBMjAbLVaiwm1nY+oW1DLTmRnIfYe4dkGErONazF+QzoU9M1+Snbmv+ctf7Ju6DlqOjhOOStgcWI
cHxFc/fs0YhOCAMs3kiRBWyRtWKp26PV8v0lM7DM4FQHdb3defk6PFnKE1DSjVw+Pjgn9NAmTozv
SehygokJyzp2p5WSQ8OHdb9eMNn8sNIbCzWf4sdsOcDqOJL4NQZ2YGqmcoexk74oSEDNfSL/w4Eq
w/8L09S+Ves7iNtdTbHiAJT1cyRp1oj3xbgMF+ef/CeFjKywt7aET04EWaRTLmdOVPdVN3rnB74t
L56VS0FIbgbnTmhyKo32s5VCpOKkZl05C4HSLT4ackVZyXoBCmVCyKn05E3zZBeFJIji3FwpbkT0
eSK8lMxRAi5QOtGbOIQow/ILch1j2fCtB0OqlrgPyk/g1TbqZTVue7gnwxB7L+Ye6cd4gAYzYlv7
viuttSbAuWs7v5wUF2LuSJLkRgEDb7PGpEpsgfT888zvQGbWTSqo++a8krctiooO9tHR1NAZIU8p
xehl2V55teY6DgcqTXiImzyHKcC6S3XXY1xwflZFHXZlijzt6I1Lrri4kGIHxlKyhvegfVLu0wSi
P/MRAIHdwbF7ZM7KP7NfuQO3z3rP5X1AUraZXJM+YB5ZfvUOtbIrEcVQnpLKBc6uJrI5PsH1gtn8
E06kFyfh338bROGRbxKNlb3MbY+TMdnEIsVHfzjtnL57vTxoSH2IrKKA/xUaV6mcvvHMYQFFI/Zd
SnAJ0f9s1/seTQy0oxi3rUwI7NRJmUgxcr2DTaTUG+HW+yu1cpIL9P/EVHyREfYbWwkBjq7thpuL
C6LsIm+nszxm3QI+jzWWO5QA5/u+HvBcHMNZOBEypQFHrxgbklWTrFTiVUeoM/VZgqMW5JXnkreA
7sKekYt1CeDP3dpUo6A/7y0Js6PVolt/MYE/bMTxqemCJsabICXyQze+UGm19AZTyNtAREW5iF00
5xpU70u+/YOZGvYE11ymztVnWrtyWVYzLR+0NwVULPeGEeavLS3mrVMClPqtL/NgTC29dSnfZgLh
4wes5wM5sCaOzpxpKUQfuT4Hde3pnkBupGAJWL2z6Zgh1jwyUxJ+VnGdVmi4RZqBwHWztqEVeY+y
HKUCVrgMqXFRPfyOFygju/LMpmDEnB0+ObotPnGx1iYFNEdA3QEY15H7aBwP70oZPDNIk7TrQTE/
+Fh6SHpFRg5X4xdtDAuFQnxAFBtd2WNXwt/K3SeExFnPGMMlwIY1Eq0n7wMjs5UBqI861UiQ3HNu
WCGzNQ6vkWk8DV4csFeA5FZWiDraPzyW7geh7tqxdVTaA/iGQwPyPNIXtdw9o2Q6kWJbk7s018Bv
zD8WKtPaU5xgCugcgY/vhpS0snZ91dOyfJQ/l/6WqASnrEBG31jYCTXd2jQm0fUYGDWNqsw2a1EM
F++WS6L8JhVHBLksodNUzoWuCCCfOdHz64bav2LhugXeZxpAga7iZ9cQZzbofueBbGX95kqCT7l4
TIrv1cAj7uleMBxnoDorwtx9IA09H6N6ussu5Mg1GH23F7Gz/qH1bdjIO3ZGdfpoF8kINuBA+f7w
GX4l5sGfTX97GDXZ7AKQ3kNsA10w9DtYNfdr/VmeG7h+7y+rRofVjy948cVkAsmLzxL9y/y3K5lO
3Qd1dAsHNC8PjJjqf5kS9eemSxBXSzsaAwsOoSJUYIhvaXUHozpvmBIoMiVY61u0U9n4/JvOF1Ld
ZVtuqjFWnXNnpzjAKx7+qJ3sE6fg6b5B/8nSz8B7EjmPJSCcl0ctPJwT9QmAxyRndXa1Iidmcg8u
pCYOWFhZjMOQMVD72HvxSEI07Pm+ke/bhfO4EV+enHb2rOyxQ7v0bkPMG4ApSYbAN6+ikoF4aUbw
oarNvhJ2ZEjXPm+/HAYXwJD/rl1MFQ21uLtSDceDt//STxkZZ7vv8kQ2yp9Vgb3xkMUHTOhy7KKu
kR48M8N/QsWn1nkDYBbky4dRQL0gEYo3fcowhS28QZDhOaBhVMOYEMbcqTL6ojXbdJAAscodYA7Y
+bv5plbZwlifxfjxxhQg4b5F/wrjDISxSjwab4nu7aRwiXT1FL38lIa63rcm7ZA9cnZB0t74VOwO
sI2Q9DV1IV/G8S4a/1JGzr4GMIKi0idLlH8GRMQ4//c12wfpYRTxo3+WVS5nQpWD1oqxpcOf6foW
+AuXT7AcKJNSeQf0JNPVikuqnDBaM+5Yr/1lr+4UOg4s/LnOOD9FMhVIeN4Fi+Zdq1W11PT02JLU
f1r+Z6W8/Llp2C/x26n2u2ckby5jM5mJmhYdob70iB8ICdLWG8Srd8bw9S0dg2AdVETFsDzhhS49
zFBdP5go7zsyvfs/dmYA9XcCRMknDFTW/TebOycQTsGwXInTz76tMIkAwJ92jKwHclJEIBkbrcLw
YJSzjpQgBveY4+iMzpmlUbjV/nrKTHEOrYLoPnfl5FdZDf5CR24tHg7IT7zpUXNCl2CSkFORTIm/
xcln/yezGyZUhxB4kQiyoHOxzWsuqjMprOhCyx1d/3E151wmb1j3d00f/6s6RT5mPHC59Vw6DJlf
L79iL3EMJNUVZr6dhfkqBdvgJ2R1DtxWfxtPrEZOQefGPvzvOAfP2lCxSzo8/zl2nNOVtBxav0bg
75lqj2E77Otk+eCuIldfywuo9eWkRM7GcKhl7A0AbrC4PNlq6efatamx7U2PPx3hiGujguv0r2ty
lUy8dBHSb+Nmo9zbguKW86BLgbIIrmZ+NqcVl8vaVeSyWRLDnd/TFvl8FxHp7WvHyB3EiabJioz9
SxO3qMOtEJi/lGVjoQR2Stp2Uzuaw7VZt0tV2l4be4CSp+kBs3qC1O3sOCnafBXsK0zOcfIZYby6
Ohk7JbSNjoXvyTlUu565+5mNz2+ph7LqIeBeP3Fy0WczXZOJ0wf8fU6hoaF9XNoCf8gk69FC5w8U
p2YKN0CcaRMFb91SnhuBNzvJOPJcf5RWE16EK5mDUsqwWpXlv63YusJULb2Z2Va0hrYNq8wFAbCb
l8j/EPoJj+YjTdZTD7BbnMb9LoBxnHS4gskmntkslOI8s3jeX0t+D7xHou7zt5MDwD1ZfK7PbEjK
9htmcb17GNfGHoXqInXADXMO2f23sgL/lJFvHKByPNHpIHcf28qxife8VBNVDc5lTlkG7T562y0P
Uikzn9TOUkya5Lz/MtrJmXZKm8zF7kV+HMmMwjKVlcb4GpFAtzkvUK8JOD9U1FOoMf4Lmx8+vCKn
w9gZaQfAfWrTe2x/yRByhlhoSDat0K04Ow0aTzbcAPKReIlRgQVELOfOkUiQe6mmvsZ87ADixTed
gSi7R/66EQQoUfApn+OLqkhcTlpaLJxrqmviR4K8CiGcVbk8UG16laJBPF5Nc8XP0KFxgmijio+X
8v7ca8RFSj5OujTy6ZzQ0E9+GTw7lqTZG5C96TfWT4PHBXEwl2h6i8HsXfVwGTANk1qGZQLRmrxz
DPKFhDrqGHd8VCyf7F/onqU0duMAxtEqLC++RyFCV8Awkh4PlcWLoj1gTbvtZQKOluTtnuzv2ASL
C2cAkgynQAtNl8zGLrtV6+z+DB22LvaMXTmKoIsxWzP4WFYre+ef5cIh4mAq8xs0Rabr6uTk8yln
pSOUGk4Sae0jAiDR36ZNHZ6GagVzndbLJHlAigYUwDiXnNPEh6CZybUIYpnx8TtSWY8aPCVAXulA
U3JW3X8YmU4PFxd26zNhIP27G4ZbuvHsJcOFEVn43pICvxjVUL+VaKeL0JnvoIHZsO8YFQH9O4aZ
cFmwbumcnQ2vRNX3OXEU1vwV0sbXFGOkKTAUIENkhmnGAYLsVSe4hX+a/BVmBrcd/ED29tFERBZl
DoU9yqbHyJlaWJ1ZJyuhh1b7YEG0QC886Dh0sOrsZuDXf9pjcadLO7cqbdeN94eK30D9ttr3F6np
9eACap9iK7bMXkusjBVsQnj8gQD9ddIwoOQ9bVeYA/tdFTOSwow5cmrPYAjGMdhxIxsVHQgB1xsg
MTmIwBFA5uSuxfpJoCyL3KjU6wJy3vuUM1UOceMpUAjoSGh+n14AAUzE67rEEYW1XUxMoCWFgW+A
awWn1mL4HPecaawSWhQVpdByIAwW+3ryEfRyKHXQo+NTr7/PSxOGOe1GPQlm/hI7jzEtFTau5ExO
WTEKRflKQgefu6fou1FxSZWrbWRU613HF1u8lYt0NLJ4h1mttgt2OBDHhlP7beK4G5R8dlLUSbUy
BrL+zDkgzKYxVJ+YwJgKL/en5zf1U8ySs0wzZfAoNeD5gkNd/oxEa0PS3xlaNupx8ZJnePKkt7Dq
Bd1m8zCutg3/U1koDcDjUkqWMMC4IcAZl7o5NgwdIh3h30FzKdbVZRxjzvz5MynKpGhYteuiki50
wT5PSMU5QYxY20qEFHHp8yypwjCN9L/FUVYUn9KJ8NEZ4u0BWypHhrdz2xJaK5YZCRUP4s3DVJnp
EtNA2+zRjkH/ifjBqFrNab7PP5QWLLfrksII2o60Rt1DbceXAMwmhY1d1pemDQocIE1vetCOOgcj
ZJ7a0UVaYLFYL4DhuGNjbF8QTxH9ojBf5zSnNiZm+sWtG3Gz5L6MuLrtU5bMQQXiCoBomGjLQDgW
bm2kBzdOLzqzjtMGzZuLfk2dDN638A+UfSN3VACT6P4kYdr1oJ7mQWZHyVAtgX/GQhQwKGbzDrvl
K3F0toEOwu/4z2UC3P3lsFSg1IAJOETbwZXAIOq1Gjoq2kh+89rzt+aHbtTU07C7XaeOQZskKVDf
eSXjeRpETI52gbV5P7araGSBuSk00vs/AU64RIx2Rnsmw8EIV/XzwDrXBRtVus3sKKKNnY/tO9/Z
IrRMGxQAsAuphS9PlkIITW2OiIP1htxU2WfymKRt6v+PwCZrxmpsE0zycAe5D2IAdc9ah87MgXHF
eBzr7ivdzaNn4R2nmpL0CLGn7R8RruecRdZYDlMPeaB0AeVht2qScJfob6wqqOeCRx9BSb+XF8Cz
neCF4nJov8yn4fSot4WRnE20SVSa1embbkx+3adbe5elrBya48w9pvQ90Il7pwncCUZ9c+DV3z5v
dN1P1uMPZ6id+94a73VMgC4jd7eom1SnrKiYseNRKWQpeAn/ccqnNwoQ6T/aOkdESwMeOpZtf/0b
uTRgphoz02zmIUiGxTOpQUcSWaVyRD84jxZEhIyFNuq76icHZZaGlUZMCzSLQEFmrxau/BMqYhPR
JhsgmyLMlG740I98WEjDnVp/qPluYdVjFATqNozuZW95VGC0mf0wQgkBARbAuJX1mNl5kufFr2PO
CQfZeMWpxawjX22KYlQ3dyqjPnoqF7OrTwPp8fPyBk33U4Id09uOv/Cz09MD9wwq2pwBwrsiff/y
n5NDWkVaq68exDB2HZVElIMVkWktjFIAunl0W916l2swZneFx+JSTW3UsRGF8pohhJgZM9ioumx3
prJ3TCjxgTUivHsNcXE5ygZ6fPgaj3IYkAxkpcflz4i2G8x2GP0ONwZpG/cSlIxQcuHRTSXDmLdh
NjnDZzvL7Utz3y00WTzrD2RxdBYz+m+JvSaPG9nKrhsgSn9WHOxslVVlUPvvpAN9jEmuenEyUgfB
J7DFE+Ivu77qd4wK9CiahXty2WrGcJnDIX+bvzms0FHfMRevczQJu+MXleX3YHCH9vcQVYG4z1zo
Z0Ste8grgL1htQ3+1UemDuT8/KDOl2Kbv6BlBA3Phjwxo+n0rJXWB1rkKaZJE/j6BHSzTfCaSbuk
kDqI6OTT3GNM4/6t/nM7y0HCd1+CGekUdNuMVr48EWzYAcKSqvw981wHaUHsLCXcxacBILxlbPN/
trMRdZdxshEnRDdAKQPflPbo62YlJ5MbYsNx6vMBhJ93vQqVLZjmxpRGsUIMb3W7tlLrOqnlypTV
U+4wgVfpm4irqEd8OqyOE/h4lBgnipTpIBNYdOxGNjyYusezUOCvqOSWX2+csMLvlE7gPdP7g9hA
Rk1eO0qwb/B28cZaolyPUTMFwZDdQVjrOaCMfLelQ+Qc3sP7yOmhYeS6xFEuFiu8MxkJ6FUSWHoU
jdSH/NliDaxy8aMpyCEDAOIhHDBf9aFNx9flo0Gan3SlLk2EFpAUDhrfQRqM0sieNlRnQscv1tGR
PBSWeHQ/M/vAr03v3v9pdllGpHSWVy9dmcXn6qWk0LLskkEYL2i2kpF/IhNu307wfxzV7Gfv8dyN
n+QYNAnQI94IerJEE0S/gI4th4wN1hCZgtTpZDyGWljoBrAbrOZwW2GowARALhglCvyDChnO9BMC
LPPJTeWufpdyIQmug7Pwyd89gugGueRUAypXdL6f/QVSl+5CAhH16F4H7YhLihO/qkebTjdmPf6j
KEaR7uRT9yzCHnQfYXZSW8SAMYxBhSlqhNZWvmmtPLdYJwyhFwK38J65LrpNNiBUCvU2ZYminzH2
0J6Pubsol4Cm8USdpyGMgGWjrTdKZJOl/2ilJPhU+2eeMsbYdQgArY99wC9PpLsE6nnTjSJPJpRl
vJpqbjFGXGaSy1c0cBOnY1MdgG0g69c3H/PtKs7CQ6DiyV+lk/3EmQehtsE3Q7hENDtdiZnMMNyF
L5GsQHdiFl+kT4tsIuvYQy6o8RWlp+JJYEUfl2MSkWDExCisgaunp1n72RSxb6BeMr/PMLzddjv1
8YEfBQZWo/oipTf3vueww/uG1FYhgvuJXw3cT3KPTzSx7Y6YbGCc5YVV2LaM6VV5kxofkHjN9TDY
SJ9HvJnfQ2NIWOOQnvtfuLOq417a8jAEdVuJ1dRBHVqLvgP8x+E63XGgHyYMgc2aVlx70D6I3nnQ
YkX1TQSXsKrEzku68sirQ/GF7Mar/TbXrz08EfyGcHWHtC+K5cAqxX1o78IxjNl7EKtOUuoMKnij
0008aNwFxORPuUE+dY7YJB9h3DWEEFCiYzIMAAEWpwWqxKn3Pbn5PrFUKq2gClDMDgxM4qXpjhmx
kFealXrLzt/PcM6lSzBQnhuuBB8ugjRag/A9eTxuILYj3+ZkURoF1mS1eU1RosKVXtXYPeEZOhdx
R+6sVYyGxjddvKfUIZhYqDdp3yvIdDaMriU2AXBmat3zEP3cO2xDUTnXFevmtyGo7hGeSfgno7oD
JDeLx3Gs1c6J9XY7TTiiXn0hH9uwmxkfNX0bWagUKf8Tj7LqT5lnBXIefSce0HuD2DUWId5oqK8V
PkaUGv0yUOH2drQWCFVd8HEMPDs29RUjEf/h+GujXxfH2xxDjUAz7f7HOJpcnMfPfrr/t7aFE2Xd
OWwvmjbtqLNrhlugRF6ZE1bD0boH7mG8298T+RNdC8gNwr4MhJ+oEiZetaL7ocAyp3Ph3Z1jvfYC
s82FFOmhXqY36QBoTTk8D7/y0XJMzArKsIyK7t5pj7hpYU2EGvQnPMgTx7lYM+wSBY+1Yu7RDFO7
qlYIZzqRF6eqDI9vCt6TZ+d3m5eHWQWvbRnKPhkrqbW2wAiCj7lKg5LS3Xcc1K4z7FHcnBMWJagt
mEBuaZYw6EdaoQb5PbyYqBZulEEfmjwP/kWYjATPZHX4ukR6unKD+2sizm6wCPlLtA5saOkhL50y
V8Kk+PVNQML3JQ5aPSkU53QEO+VXFO12VKpJ2sa6OtX7Lnv3Cl+p6K+f1dy0UbRQIBCo2STzg5Ey
7ZrOO2mBn3ixSu901JYXNrVenbBDiXhJxRTGdztDpq0gkjO2IV3SLc+s5oCfz7kcxQp16krnTwv4
5qI/nlVJ4AfbrGAPKMUO9t0EjXdfZp93QRrW1jvHUky1C7QBGqLph8pASOYbfCd/IfKG7d4Xr17T
jMCLoOfvPcIx5DftnN/o60CEpLdpKi/xugGPr3MLw0JXmYMELIKDlqNUn6XD1cAHu1h50u1szb+L
5uynqrOZsTq8VFuAd7Eok/K2/Mc3igMuhHoo6x/YNRyYm03JqWatuYa/48mcoUuzPzrDSu3PCpZC
shk135fWQBtn8fl0EyREslxgzqHU8Sz+o5/ZUWMc2uAmiL/1LHqHIQa3xGe8kt8sp8A9v5mzrwd0
Jlgj7IFNck8/QsQpjRMqJTE3C2bty9Cf4h5ljbTxH8cpw1hRQfAcGkmH3+RkO+TizKGzNvRbY60q
jdAlU327Zrj/mj1qWTXR+1lUeflkZTvg/yOpYJWtmVcN+dqAyYD5hZyrdHh+WwvtbXh1KaIIljtm
635+q1E4MenmmMzLnKE/e5m63Aq/l1IvUquNIIz+/YC+KA0m+5dCaswwJq3Z1RfRdwhWUobaFlO3
f4hTZHNxya29nxzjFYKvyEQTT6d9OIyaxWKic+V22OAW5T8Tn3N5GOCsYB7VSjIMRs56UO/ITyxm
G98QfUn/9P9AcY/DMUrNbXZ9mokBLSRlBhwXDvKTplaCHJQq2tiC7kvwkfV3U0iZHjBB/FyhuSfE
1S7rXLW1TKque8BOR6pjxdIZdgiC7pY3bd/VSUKvtvKt2EMVOLleCmRyoPysk+95HB0kD4r+dJRn
ooVf3P3jhp6t0oO8hwpmc9oTkaqNb7wAgEQZqFB4LZAWo4wGacOCgCuI0gVpd8W2aU7lwxWzc41P
Y55v2RHc6z965QOR5+egBwYC+AtCFGuUfR3/WMeRj3BDmJygVbwJNcVn9VUHYc608iyth1OVR/Zq
vjilTjF14zEwXrQ3uSIIDU0XeZ5a3S8TjLXveFUHP0oAQwCir37VCikM4OZpwra2bk5befNFQwB/
gLZyTBzwd02lQKhMejDuxrnOcbWU9qhdMWcV/X/quxFwzycD+8+PJsX9dDMlKSYXJDfsZTV2n16V
1DEOgCQTsNkXYL+jjF7bE9uGJUzG+Yk4yynFLz1k9dVQeA8Kxr1ppTOQGEWCEzpIhwtqdUzg1z2E
sZ63r7rC35EFemMQbp1l2z4e2OqUF+nnNrqtkSWSASE6kVOyKgkbIrWPs7VnWPsqKM3MDfmkAUPe
gzRVTayaSX7hbISaDFo6M1lIYLLMh5LP2erUAhpDtS/Y7w5EOyP1HnNOOCJnMDmMrMK89p8Fp7nW
XMqxQ7fyPc5bAnCZ2XFrL3Pz8PRbAJsTCpvIP+odEOqSVEVk2rT4MHZE4tqBj1XHZmmxWkJPxFW8
GA5GbO6TvzLaLLEXrRuzTn/wTLyOVTkap+rn8WiYESHr1eeeubRIpNzmchrnNd47+mkIRnVOVgQ2
2gYm/ToAxDE4dJDgh6O902yOD9+lLZK6xpadg2wjyakl5gRiYCOSgMOPuoK2FbQ+Y5VyKoZoMHy1
YEw8LHj6dCQUYPTWyg/dQYg/7fgRk8NyYNjBsczeic/U23Wx7XlVsWqWDDjpdZV4v5gnz8XGtElU
Jhr2D31lLWktZASexl7rjnV+5ByBulDZ5wI0O+jZFIufUX72pTBn/z23nlpbBBiyk/3rp257OPDc
FyX510F2I6obr9B9V6y0qPdoJkIAUQ+TYN4XK63pvqSgXrTqCaPdIL0yHKVQQR2ObOvjisn9r7ZQ
u253bGhI48h6SEg/0aRnfyQ5dA+VoFLgV7Vx7va4HjobjuS+oPd+H9RzOh5jwe0ECxG0qhzyZRk5
mBPN2c8SyT0pYBi5D6h/UCXMuBDdrQYUjkaK+2ds3gV79y+eRjjEWCgAceGHMQZDW4ZbuEjWmWAW
U2ETt0qGCUX65vBW3Nj0UkxU34Qj7sY3cTFrAeENbrj3HYONN7PkAUrg9IjOLqOCGgtvnkO+a+Ol
iFJL68ybEe3NXKKG4qSrxs743fhkg8fYD8wFxuJX7m7lRNq/j5c/MCuPNQYFRJftN4g1tKCi8hio
3u1zGRvozLV8GJ3VpwMvNGqczGR/2zdcZDbRgR5BbHalzAJUPXZh/dHGFRVujmWAJtFbCwHd4DSg
a0NBRRWHdYL+e0Cy2/3h2gBPJwRCAlxzCFkz4bhKNm6OImgFUThcrxEWsBcr763Ns4CDxeN7frNr
PfO81wLN3ot98ELAD+uC4tCIa92OC/HDHEh2ok5t25GeiZWC/6iYtkV7AzZs0jJLxppdtIJ94LeE
VaxVwhEnCZ0D9EGLFJAqLhd541nSPhlTDlQBY2VRDlTO0tx5SHIuxEkstXw/JJjMkQZSKdQ7m+rY
hRVVgftJa6iYKtdztgaQie9SumYojCg5lI8BDutt704RyCil27ZHGzoSMMeDxuuvLdY3PAzvhPYe
2wt7CFWcAXzjm+BFsnnVqWjY+25oydh7aH93D/JR5cWCgZwnL+QzqSbgYFQcg5Sn0c2ZgWM+MK5C
ZnfY4sQliXJAQazO0qp2QgrAT+VrK5g4PO/RRLy4JaAYbWS7jWlwrSMwIxN7Lzh3HYyIHbzF65eW
5g4JJzDYsDVg/774PxO3LiXE3K2wjhm13J5eCeE0qICPyWnyEI8BAFbGqBADKspfhHNocTqtNHjJ
llNYUVcoClHvD4NJz6pFsyU3RAXVnC07IKYIcUZJvPL0W+wWNRs7voJdWi5z/0/hFdaS5ovQEl3k
9KkHkmbk28IiIWoxs/1+Gf4OWestTAR247fFhUkBdB/EKvyq0/9EhvTbEENAU+FN+B/xwJtn2nX0
Bf8nQhiFuPkscFeVee0DprU25909TvU3iObBvfgk6eJnjzQiqGZGn96rwRt2Kw9dxIksUXUMmFOj
t8x+urqG7TbsHOnsGh3l4M/PB3S0/X3GYwWpYXRIBClxXPJK6JhjW2tVunTGkzy0yNhLMaWGtNuc
OxaBPypcmyN50ftW83CUwS1uEMGZV/lBvjKgGkmWrNQdJ821qp4Dpu3NH0FLYnP1dGHc9IJZgxew
VG8T+1u2Vn0uMRP0wK3eIPCXqhliVA5sQangEBdHJbqDal+P90zw133V8ggELJPpJqc5AA1KREln
87fWUtdg4qq0VctGFNwrTltyaQyFb65E7Q5BQsn8iCKJ23Pwgr6tYT9Xdnt6pgWiUczkMjfJYHFZ
ClHFqJYPI1Of4uVjfUtT14+rJfu6K57d6IKM1EUM59SREGu3nnmUwV0qS/lIP5wW+6N1jhNLUx0H
iOnbYdhujfGMjCWGEKHVV9/o0Pi1foUGvTiAyuxYLwqKzEWF/WbGVcAjd+1kPXH8uMsShShPp0bg
lTc/BZ5Me2+PvrQ7n2df2gtv+1rrQafUsQRKGclVL620AsSzKcpReH28hU/19MDsBAH9M51AKLWe
KKacfwtPuz2JqAxIt49PuHuuqADTDNntRaenZmcw86C2w5HQ0aQ3BQfm0t5FVG7+THfQXmtSKUNv
7HkwBEiPL4L8mqW62fp4B3hGGAx2p4wlQJhUYHKE5DvQ2pxT9xGL9ZR1+lN3ByAUe6OMMjhPqARV
Y9mpOde1zw+vVH19RkaAmH4W/POo8lqHoNqQI0x2WJ8eABvMRyZKKFGLQh9G/2bI+tPp/XAjqAIi
0cVMOAhaAvJy0lc8luvLhy6ZbKfXbixs1n+SwCc4lXM7V+W5wsoIVrgI7ZQqtyB7rn/r4Zp/TFaF
GJ91cHTO25g/IuVjgF+cuez1fw9HgjCBoUgL4+gcbsHJWQKGDtqrmyWYU+C1PIB9G8OUjwoohZBN
slGEVOzt+o7Wmy268+C0ADjJKMFOkmOm2tpoKyGO1eBoBGil/fSi0aCU4nCTAwMyW2R6fxWcZ4NQ
QqVJ4wAb/dQd9wYYSbiRiInetWZDRZvzK1afScQ8Avc0i+EgWq6MLynCjWPM6uUZfHTL+yumt1kf
G/N8wOhsu7oftmn+jIq7kAh0vREBcpEw4hvMtIeiQ2HM218+eNLGvkzjx+nGUrSGil/1qeHDnaZN
4KvJlCpeM/+Mb9zXazrhz3hw3pPFDPHN8+wWjcc0JdH5RrRKNS3a7Fuuo5WqTNIb7uAvCPBCqDlv
YRV48Th+olhTvzguF8ZMzxBv7vVIafJgoCez2f3WvWqvMX22FEFOtQapT5P8u5EZDCjF+CKEhOI/
oc1vss28xU54qsnLwwA7bR07y308xv8w8Get0LEBsCu7f+1f950hQeoFpvl2u3OvkXPJukyMwwxv
8EvtHv+VBxiCUbbKogmWdMFrjzrldq7RlKSsUIykG1APQOMo4p9NPFXvXQlo/nFAaU87zjm17Hsz
99FTg24QUAonzaZ+C+jrLGtPrcaIPUoimI5WYiujMdLjWD0Hhws9RshF9gxtho9x/AehdMlrNZHc
XEx5ChNE+XLjAbzWSu6EIFwIkGO9XHjowz05BGQUru81qjKmUXA69PfYJ9FWmbed9KeymzbyqE4T
I8x7aSZfTkVjC7C/EeV0i2AOPIf2LBgWMqXkxDVgWo6l5DsaoZ/hpS2w3aLTlIaLaqFGQ1Y5SRjz
Ynspki/CwBnsYeCSeaCKz9HxU1FJQFYS73d2yw3TWwDG2I10+lLVawZ8BfPdhlMCfuC8a1Ak4XKX
UyzDsc0zC8XQJdEIWydO4t23/CF2cTTALIoDP/tbM1HA8vpEuw45cboyj0tbwuXEEoSjbMrSHiQy
1qb8zJfx7IDUYmxj5r2VohvpQ4azajRapvy8q34UDchYcOte3R+ofqbc9cEF6EpLvVlK+NSs/oSb
Y6q8NYcN9z0uA1583ocw7kRGa29UEYC4gHGno2OMldOwAOwldxCOdFPq9wMAebkDR3fjMEGUls+N
1E1kuIuGynKif9BrrLEYTXqlpGxu4F7R/9r9ltQGO/dC5v/TtrYB44CCq+c4NkqFUV7ozcJu17qO
Yk8yYSsieKVixgAUFH7HKWF4Y2gJvUf7u6zA/uaGKo3+ZX3kdYIF2XtAZ2th0KlzNnTq1uOIVg2V
AY0uo/JlOhgaIuG3HwN1z/6TlfDeLyfz/qzmOdYZQCesXl7AcWTKSWkQ1cUFd3+JPSWimPNov/js
r0LLtghtYm03EADme4OuNrBUXG2wTivYMt/0QPtBQzH2N2Wv4aAyQqLaRZ6exv+H5hV4f4XkI7X/
eZyqH62NTQmsZcPR0lfSHxjG89Xask4zqXPuJjbOSs8gUh2OP4VLwtL+9x+Qrg2fOZ1dyeL4gi6D
H0I4cle1dYdDtrU9Ofpwf+Z22QdJqXMi1NduSx1PnxJuCIhY2LyU2YLGo9P15+0RiZeaTzznUdIG
+0dsuz/vCIi05aRn7bAMwj8+gnnDFlJSSsdGlag8ERWxyumXxu3QylU6lvqezKFSqsx+UB1dD/qF
hY/dJ1+aC7XNEAlwNxMYaZxoKy216ymfZe7sqylt9FCBJMspvJl24BwHDor6WG6WA7/xLw/JdJHq
Kr0l5WYqWHMO25MOGW5TjI+ywoRtfq/7O+21Od/IegxdrvnSM7eFtkx0MEFzQESdhWCRx6DfPGoK
mwaxUdhUUUyfqC0dCL2x5oH9K0YD3i7gCU332Eh8A6eAhL40pJOZrb41yHz5MyvHLY2Gk7Xpxyzx
rgejiS7Y+vLLnumfOQNCXzbXRwtUxlSUc8AhhFgAhCNL9CfUScm56mdiCjMXoPkKG6Il9fYCdck2
ZlHU3Ev82GNbfXgY+ZXANmXQBGY/qSAU+Www2VnRlM0nb8lIkYjH6mNGQAbueLXkGiApl1X1HX3y
nzs6ofqsIXpNWMmfTBKDsL0vU/G3oHUwAGutthK4TImr+zJBS3siqJ0B+NCRWMoZGZzQ3WcdhYQM
G8EzeuxQh/4tUMri6yxhu4BsbM0Swu3yQCGPfdscr+oZZXVgZpw6jYXuiNeLP/R/giQuXX4wffZe
RYYSZE+Tt+shmwWmz+77qZsISh0VDqYJWsv8Dw1qoCWyfDiyL3bW2xRGQ5U9Oj1OwvTWxPLZvoKR
N6t6ti7KW0JbcHOelMHXNSrd3/bqmjvk79J3AaDwZBQxm6SglefCd3f/xiQhjerCa0R0fWl1RdRk
/4Pcyq1MhTR3GnUkOOzD6TIEs4R6KQ3b7Xuo8lBa4q7W1L2aOdutcPiogFTegTWqmlSHCZz2Dbls
typmHqjhd6UO24UVNFePSWqFbf3cg4y6ocriRyv+/0JlNVe+sTuUYloyrgOalJNKJhEqv9dbF871
qvv4ld9EgfxHOiPMtz0bPH/UMqWxUmSUSmt/Se0NS54pKVjuGmK8OnQdsBGL+yVHu3F8R0FjIUj1
FXk6P5v0o0F56mod7lbXvwfJVlYrKOtWAPYJyTQl5j9fBx7IObwNBLG8JOsia7L35vgRKL+xcuaW
JHIyPHxgImo/nJzblOXrmGkXHsRizQ0PZrFFcSuyHr3ZFubIqc7c0NP7H+iJZu59VqfRiGy33T34
svsST8/+WV9/po2mFAQzHnutDFf7gKTNKf+4GvlCoxJ1YcELhokKZ5k++UxDXn5xThWL94yUV0U4
ttb5T5uX5mB8BTHXGhmWGkoULKpR1BYzwyy4z/eSFsqWrN7RD06E613oZzWvynR7d33omuHFAx50
X0P16PlOOJDcXM5pyXy6isf5+d/PpEOhQnDjyAnWBXcCbvXHVb3nOruCA0cS0iLz0SsxgCGCFt4q
e3mMbygbY2OncvOUlvTw7BEKgf1ZF6nGMrkIH5bEFXCT1e0BemHoTgwOjxeK9JAIMyI/QYnYY254
brXycTztsgsWlkaPoca3UoEWADoZ0QVCiaRkpF4wT7qIb0pabiNF5L+nO04U22GDPPAG0RDWES/r
aTTuGS+LntowAd9vYViAT7XomhQatGHMsPhbfQnZWULJ6cWLWFjlhQGoeXB50MtK0ueREex3ff/h
l3a2SJKYXlTteiiQolYAte2bFhSs23SfqMDMSdw8i1CRAWj8YQ6Up2s07uMf187vTnrbkb9oy1a0
Ft/jgVI+4NijiemWdD4twvf0PpvDbGpxaSkbRySlPhIto9TYvBwWDO8DMlQ77qzQ8gOIbIeA6iZy
S0AFGBgJJXVFuhOJlXLGth97d2RiBeB7j4WB6+DiatBmAycNv5N4dH7k46ssLTqke78vVu0R8zzT
q5X/c5B7hiKJnL/n/teWSjz+GU/xHan23B3J4nyAWcKjWVmSZWYpDvP4jZdMMr1rfC4iszrniRjP
F9ZQQXkDkXXBfw/rKOTWssw8pldiEv5KIyFcvxy39oXIzFLdBxV3/BxI/oK8NeNqFwclz7owQ7k0
nynHri598slNSz03OrIK6Ngo2FwPmO/12HBUtAkCzYh4MLa11Z42c+zQ2zp64B0G6EyCi3rtvxtL
ubklz1I6ziaX5meuY6kYBAxq4oaFuaE2iklZcgvF+Ix6M1/ALRPdnMnUfaeUF3Pr4gKY5mRMzdq5
LDGls+U8Px3KBC9URf9HgMo/VzpTIcXryc3C4hluHnFMvvpTk5xOiH8XWnlgESODQ+4yZ2t6hM6I
ozwvLum1Nr4FF5hmKvwmqq6c0Gzre/vQROELdrpQWaqT/rVy7t+STY9wVRvblnRh81pr6qutzxai
zWvcNIT03DbDjxXVtSLOIxTEjLeHDYmcZhPMWXTDLSdnNH2dCdXzySuAe+OxnnydTbWzyT59SBE9
DXunJfbSCEKWn4/TMoT5R81PmxGQcAzRzWfzgfpEnBFkJnOQnp9W6IzNoH3SHqhWRfSRXxF1g7aJ
VFh4mzzwNMkcefIpKJdCM+WLOjeysLnb+7D8IdT+lEDkjuKaGNX3qmGreKw1vRvMrVErr0xhmSa2
OXu5PpRMUB98iQyLlhpTG9unQHF00VgPtAuHI5CvWlHPVFmNPHvHHDA9/FLZgl52fASfJ2Q7F0tN
wbYMz7KT7Y8kx/9+gMc13JXyYy6ZgMrZmoDssalV47SuNuqos6ULr/bU2Gm1egqXtJOwcUeWSDrC
1o6C4VC20aed8ms7JSOA+Ldy9UClv8pJ3U+g9m/IWssvPBsI9yNlxkgSKeyj1msamnBr5HcAgMoW
9csc+Gd3ApWUCOpSGSgQCZJCO8XLXQIjzVlH4faQIzACfxmv6EqjO8n2lWNnokYQp5+FlgSxKdWE
J0rxX7rkmwnnbmhpd9z0aI5dNOSRIQ2OsA8CfHEcyPQ2nX+MF/3RZn1n0Xbpg+ulkmBQ4cC9SGxG
FCtB71dycQvmjdB9pw5Fto7lqSinQkt6Xw2ywOpIezTVZtpEq6AJ7rRPr9KfUjEFrxOhRQJLONze
0lmd2VvSNkPUD/SYLQx4X4zFDTwWi4/5NqMhHVmkRvCEdBQWbJCmQNS8MQ4RfIEAAgyPIERpPtAT
umBpU9Sm7uqQ27DrxPrmUzTorOzwP4RTz5S5p+afWB0SiS99uavm0csU+2vKSHoFngnwJ1zD9ZXD
cD2AwuRIVdeNA5iALVPgxHZt70YvGv3c8k0UtQUAHwK6cRqhK3av2YgV9ufnzi6Yysyj6uQ8YHrt
wpW05XlxzTckydUFisw/6TRQ5LdbXrEShgdOf829wrKpyxmMh4gixahoSbpp2v71pJ7GpNgAmYRf
94TXkYsC309PXLvkpAw3BEnxxXE0/g0qY4QTUzDKqG1G8zAvxoJRkBA4Saa4iR+gpgaaS36fReto
OXULeTcaYfTVNwG6BoN0i3VFhyBt+J+GvbeNWPWg+3BrBvoYBhb1aXrEyxJDTqgG0razWUefxoV0
RFVJ8qs8CrrT0eOArH3zHy0PuM7Gyu9tbCtKUwwES+B5ncTUXuZfEAJw2KlkJH0z5ctww/CFhCGo
tziFIyS2WwDdQYm9kWyE1O1m+ztc3eoxWeBdA7tbcEwR7hapdeyFmkU/o6y/H+E6tcjKuOR83XVK
NEl58V06RAxFia0tlKDcd7vXrxgeWoSrWFy/7KYAmeictUOKSRgZ7245nX8pXLcktciyaiS8r65q
Pul09CIZdXQ+vV8oky4XcmJh7SYaeKU/R4ygYgiYxHIzTz4M/5K9fakroLrM6JSfEuyjsVR6o9LW
NXf4uN5JiQ2fVtUlR2bZ20J6f+S29sc3qSlPLT8OgS1EsavEG6IPPOqJraS6CJft9NviwMCtD8NX
1zcT5dK7go3b5MjFSrA4DSr8EzoQ9AMTqxEiTK7jDZHs2wQnmic/3xWkTHncc7C3lPcSNh3dwVVe
0/Gh9hjOSfep712OpnZ2xtZMs7Ht3RQUmJWEfEovDR+tpiIPcAC9Dx4sh8I7GkvgZKIQJxxncnhY
/WxYHEt5uMMBuUJOpuctfOAFRJVBf8HQUBsC85VhmSIIo03XPry9W+dtQFxTGkfUsa0RShQKO0/G
tfiwXvUgdOVxk7a/S5EXuaWmSR/chvhKhhPh7FeOrqwcg7vtlEy7Z3zLqqLJRp82PARGLcv51Tai
DnMLt14ooYuIMHlJwlIymUO5J3c9hwo8B55FuGTyYgjyxvrnGeY/j1gh6kKjQMEjhvmb7b2XKaMY
FOjhqOntFLc/WR2FbfeJs84hzjsQpDHYWZTszAaFe+KUdLiNL/AbDaCzYKQPO+ZX3TERUTJbi0RC
ZGV9bTo1os3dQeHS5u4Q9DRqRASreYzA6D5U4Ky87Oiqv4ffLWptokUntvwU0eoNxxricmmBIj3s
Xx8upmLkHvh90J7dULd+KFuAfP/cawPGT4UkgwsWri9R1TS1NcfVsYXO8VwngiZnWTasl+uhLD7l
SYNtyJyJauJeB7vqYku1pMZyzXFranDzFRhXhJiyosCdlH5GCGo4oDDZBTP4hddqAFw9JCaLzh8j
ts+BJ8xNVZMGh2sZkbHMCrAB+YUsD6b9DRN59fnVigSd0ye89ORH9Bo3BUfW8tUfuT7fobvThWSa
/y9uINFWuWtFdWpVarYc4PHf4MQHP9AGEjIkG0UVPnwrYHePS110+ETBX0zVjCReSVgMAz9fluqt
Deedjf0/7JtxBAk6N2yOJanItQka26nawwayQm/S9NRhTy98y9A0PrX8hscKSYcxZoJC9y5965ev
/cGekN6Y5gFFWxicpDiAPmhQSmjPkC5iIX8KT06EvC9PO+8LyrarKQP/cxyF2Hy9YAgyaRimlxn3
Aa1qMbTVpKPdsyO/x1lPMbeBANDW0L0mFYby66eZ22j65/vdIh2c+/FKnZWZFp1Xmryp0t4kWW85
H4DWiYtb99bhvW5vhr1y7Hcne7Thu9tYW4hivv+ym0VMga/LJga4g6w3ygEetG72ZoGXIt6vq65a
8TjpY4M8nVd7Te28CJmYey65KN996rHE2UZLgPNwC47dWvje5YBoIErkkROZj11A7Tt2M1Nej8gx
61MkDgNzOTpLBo32Z5j2EIStbEcpUo/iWCsPA1MaWfSP0Tbhz0Fb3LUrfp38ls1W1FRPamaFVKHD
/ImVZ40xKuO5Lkb35X+lltdDDVDS5ihytn9tq7YpKGGr8X3bZEKXKc3q9SEG8+crAyX3GeF4iFp8
0KpuUwHflBUcgb2gSTfNB2kWlmi/mo1B9PylcWoHd2Bs6EewHRSEsl0+1hyj8WkBa4Rm6aDUuTGA
b5ok5iB07T8scwbS6ZncQbBpKoNvKjosZwzGn32SGwVfKuXUD6RyiJRE4mfBvGbJ3nEvbjBo0pr4
p7776CfeSfCu8KSqGW5OfsvPkOTyxyP6sgYVUQn23ufQY3tkpXTuiAB9D7eW8ulQkViwwS+B5uYn
kbtaUB1GAOWWiPuqY3HNrySwjUrrNFgWqnh3FxdWtU+PEk3hEXSvXtVa1EM6WgztQXOxVWSWZ5Xm
xxMSJTwm3+vwDEZr7EI6E+CcDHrv93R892f46HXo/y6nYOceCzXB/0jFJI9vU04Aa3dYGRNPMycZ
s6Ma/cH3t2DgiSnHzprTyEVOk+BV+OqrAxZb9QtpTBYEHiX6i6KGnVI48h3p9ZAKYXh8B+EeGBEJ
O/eITQIFgufHPihfAl18cRMJ1+HjCqE97+WbrFXZZDNsDyNjnB6jakdfNhV+qzqmFBGwz05RnIF6
hARcG0U9OTUSEQrFd+evHlZSMBZH1FFGAkTmaEKLLTG0Ctl1ACbC5h9dEpyoXc1biztjrL48TYgf
eI9OL1yR+2RphJvDLIryH8V6T8cM8uztZ7wYKJBq+sTlXRXs3QfdpSvANvwNLHMpJdso/tGTSxYF
Jvn0YykgoHDwT1SXJgnMfk1mgibKmi5TxUqqWB+U69DCQKIVhVnd0n+CY6Gv6sOexQoTKM1Kev41
9A0qFE6d3+cVETVNTAyGtZDuT0WYvEM2Ai6xRDIGA/BJwNdF86dfS8IQfzpJnz1vTHKnWl//IKQG
71M8rEPXMg0XBhxTqa2lrKcw9TOgGGfw9JeHEtAcJMWnfLdv0Y2v7T/wC5lNwP/nHEch+rFW6z7z
0BRYYNQ7L2YPJmfcpwj4dUK1j1xnmYZu7abWG8XKK71oCqOXx21rM7ErXuDTP+fZT8lRa50fbCkw
iPgJYY2K+A5FkguLk9TgQuCX5HGdqhBEi+XTIgEXe2HRt+Z7H9HRiinI1J0828VeaI8pLVphWAU4
cMZmH0fDsAwL1VyRdvQONOzFo3u7BLfmYY7RNJ+oNGc71/tWSkMVeX+gfOwdOGqx1D7SuwUUt5hM
VFP9plECdxklpY603oCcOWFjTMEA6qR5DmRz8whgeeBGjSXhZrYO08lEZC2/mAoYQNMdF6vPo7/b
VwNS09EwvgtxyUZMYmr+teASWf5GICzE1EIVo3gBz5jldsFsgBGrtG6lwuyo+SJUSls6IyE5Lt22
lIRh/2/iK2GshwN8pULmqA7trFVWwFc8pTCkrFJOEpdsRG8jIBmBG9bLqMNf1YE04/cmJsTtgk3x
nGe5vBlf1ab24il0Vv7JtbPzg4K0XxMb37qCaPwnqbRHfHdBjXb6Mi+vI6WMCJ5nFHCQfHpSmdt6
zPxnVAHiUBq6C5O5McCyv1VwZ5EqDj7Mvef7JDiV4p5j1mkgEWjrclmQUYE1TR7DbmPvD7zCRWGK
wymC+90eaPpcUCFCtambPPlgkNMnDmjNOAawBc0qS7KUGye3XV/99pIP/Bl8kTMZDGpF2w77GysO
NymNvReUvPXuQEfoXr5cnPQjsStgOLbMpsoskSI30ZOmB9kwVMzakrq7+BwpnSIOaFhX5th7PK/m
7JDbBBLvkmSXGuAIkP3fa3TZ/fEq/x7yDBiWxZDp+l2WzOlUcUvdbZ6dejDNrzvKzdE4h1Ymeupe
m6uk2vdTBKHgKYf3aqTH4Pevok1hX/IBEYcr9bOnHpWLhm7hhLQUygbq+e55hPtYHKbB8yIQARVb
aEF6dWN3qWjwLKT0QSee/YbYCtcKFg895OBHEnJJQ4igbwQpty4qMcxngrEZqE771E3JFe/wtOvt
4m4aoIxxwDVmdVlyPiftO1mcmkQDC/StquEj9hwldo315uYwwjrPBm+/ZRvIIylFGun4nKrI6k65
d3lTzXoiEyWnXEqmNYxmNfccZBsPS6Hf6Zcm9XXrbVXHkvMHpEH+f0c+exK8rLvdVx6Ciq8w/CFA
FMWSMwhIgG+aDjEiTpw/Qn7zFUKuxZDdnFFLDbFsxer3x/ChmU/YHZFAqOW0bEAwilt6rwhqMPh7
56ZcGuHe7rWxwZxn1rHE0K66gTYpbpm1h6ZofCfklzDDut1qAk5HbWppV3XoQnOO6hLs4WY4V/8C
nTqrZN7nwy71f3veZ+cUfFM0jHEdMPHFHl4T81pzlb4py+KYl8Hu/fAfaKyItGpJRXvHt1PUu5yD
84jJkMsA7j+YQSFGZexwU0mZNPcmCcizqe9ddBHz5YaPdXMw8whlspalqXnKxJ1nGjlv/XjQLhHz
O+puRiBjB07S7EAZ+3snpDz/D3DOZGLP6fSE9O7ikclomD/EsCUAlUfd10F9ORKfM6b2qq5oJTxG
wOdEXW7iCwFEW1tBC+UCX+z41RyRdqg+zxs3JHlEFyWT5k19jinWXKvWoYBAe12t/SAsDT/mwF7+
QOGVS1RGdNYtleSZ/Wmdo0oCYcBzKeSxyybMMr2mntcTEVAavijEgLQUney/hRDgnf32hI+YXpWq
shRP7ThVxRzJn2CrFhqZ+gDGFhGR6ipW35cUma/Kz0kmmcI1Q74p6mUHwaUY35nZuvmGoP1sGfwZ
dkd+wOguKVH62kilZoSIpS4BHqtMS3umwRgT3LAC+AFiwPRWWXLeN7tBQoQPlA27cqIoZwSDqaUh
qnIHUva3JpCbuBMukXW/vrN0JXhjOUq9DD6OcMV+WNSyu+7EI0ZtHTvUaE2ie2wE94RoMkRnjU7Y
X+IocHYxWsEOZu0SgWHXJ7cowvlrEoQOsVtegDl9CsUhfPgvX4UiGBnO0PsjyA0LYSV7i8WecJvy
jxgPBTi7+qF/nt2+VIPWjVkZ6e3P8XatSDJfZxYpb1dkzyw0Rl3eVFC9UH3Qby3L7tDu8X8IPoGE
Yvh6vXb882xHupzgvIE5Oqv4vxnkGBj3NJdhqfaUkgWaDrmJOgNgd9ge6kRx30zXAqcLXVsAhBYk
t5Bb29RdosF6sGPnPatNNxmhdQkjIsCCYoCdAJoNhR1IF/VP2n130nfBZLTdooXr3GMLMkyvsBHS
3xnw+wiYIZrtfpHDu+oWJt6Ym+X+NgS4CO0eeQ+tMxVsCcJOC4pX1e0od43scXH2bA3AD1iRRmkq
CQkrmsOUNPDeOKVhfnJ9RhawditlfRHglDqjzz5JzFpqqgag6MCTuz+oYpmeLG5I7GK+xSY9gcx7
LHpXwLsbArQDFAkjrKeVFk32iXsnCOOKeHxypz65RFCkKATlRU9r1SYs6fHuUg8pZQGHGzMLz0Vq
3Zl4QCoPG8I5aE61IWf2BkVRZ6Ing/NIGbpJnNOyJIsWrIHh0n0vKGP+rn9Mh25LKmAViu+b4gg4
knA1/13u9J2zib+1MFl/ohlgDHCK17MoBVLcI0MHrSmt6dy8b4yliuw9/RCNRRTZacDNxBN6jCxs
QcnWexbUpI1AXUopkvNliGsDCKBd/TJReoUuR2D9xz+tHqk7vSo8WC2J/h488eWQJmb4cPzgmHpw
madud0NY5tWVFlxaWk3DvDDZ8fUW7nCTtY+t6dPxYU5x4qJXYYirMZRNtjx8awA+Ygc6N5y8SlBt
PDbw7QAfZB+GA7lt5JkCNJSeYr833SgLgvFj9TzqNH+p+dH5bTuFTMmZh4LCZ10t4jTnEZa+dJ3Z
NYNw5khnxAgKrw9c5y6oAy0x6zRhbBJN0DZyRdAC6fvNXziYeD3xVCEcpQoZOO9Mtmb9k1VgQxZs
QTeBPURGoEI6eEKcrA+gcOOaKY5L4mB60U33r0q/rqUExPDePM0saV2mT/419qv9dQcCCQrN1WYN
kGUU377xO0nX/xIe+DElM0SQoywfsKpDfXtyPU4F7YuuOkay5s2NPNbNGWoz3w3EcbJPoOb3kmYu
SHevkzdLOp6CeZw0g5XD5wB3Z0YodsR4H9mLW8fivxsi2K8LzdJpywEYGAHs9/6mZct/wD2p506D
y8xAH6OV4QcIWj0zb03mOem04/uXF+jOIxqo1UPUqJBIqUY2Cz9d/tMFe3yYEJZRZBvJiqpbaQio
zHe5eS+KrdvuQxiPUx8GpR1AWqBkMEQ2QNgfQ7BngtNaKD8ZttDe3QCztjPVORQI9B0vVdMnVWlX
1Jo+1KAdL5Fwq8bPcnXXQNsXoOqLup3+MdkYntnKx69ctZgJaa/3wMagvrRVF6WUqHfWVCUASs/n
cAscZhIRWCw1CndCODlla9/Ez7KjqLpgyeS2UU1SXM7kc1vivrTxxtua3YRww5it2m2Kw5hWLZ1d
BMr3TxcjmXTrje2U8cwje6Fedi7vSJMuS8rkRMUkov4kPGZvmIfTZ8ut8TClK06q8VA6q2klJm3k
ER4DAbi9EMqz+Ya2fBrtp4s+l/yiyExhP+4x75rzml7h7/LMdxs2aZkkKdPwCPlHYnCRVG5YlKmZ
p/5mvL/pNUoidQEdeLs81wevckuBIT23kqu2bFy+ijRU3vhKxNVqOT2VAQB7CZcfXEvLuMagEeKu
wVlk0llWAMRUCLrS0NuK0cohlFTOlvTqw0P2NlWVgzO48ZEvlMYBwb8/+s2kQ9khu/6WZF0EtZ8A
1Q6vX+Q2gYeJcy0YH+jATrWQu7e2djdHL/YJnj2AOSNJwxXFLMvrB8VcROYK+K7a+LMFxqex+Dd2
OCdjYu+gUZLgrBkeQvBdh6LbJzNvvL8uTschXFDj3nUelb7EOTa3XgYGH34GvnwYWzOLxEja9P3K
12CjbIirYgJNRNEdgFUyWVD+jXLkyysGciauzMOAGeLEyWcnkKY5MM4xz07EfVdnp24DYacO6u72
sgztnrsYgXdhZSVXGFk1da/rmHlyplvkKN6lNGEO6DvjEEJqrdC1HC49EQ7dFxRrxhbDiZodG0MJ
q7ZGc0xS4+FKaWSVWJTNxVGJcROuwi63HWctoOqHkM/DVCJKRqeVwg9EEaW5m+4J4KZ2QlVUzHQk
nZyqYJo7uGrTkr7HEAA6MY9/VghWnBTOdRg2Jh+B7VcCNdKK74H/YR0yQkm+aCdhpf6It7Ch/sAN
LOURU+gMrcfsJEIo09EarMCelBLtMPAYJCaQzrUSmFe0RD9sRuRuIGg2q2wk0+1LU+ttk4WYadT2
jo2WpaqfmqlvuyKfpiCYyhYLencVLSJX+1Heiskf4EGjAFtuf+bg4/5swu6P/+1kbrCrw/kZ8svk
AdR+HmRPFfG4bO+Da7ZbGEk9DNBDiFQz7MVS2EAIuUXBJM4p+LfsfxPORG+A2cYIYnG1MvmzkYRt
yS/FSeCGHiIxz7muRF7N2lftwBsh4qPX7gWTJ2tWt6dKJUoBKQ3ookSKbieHLQiNnbnWDfB+i0UC
W0c3iZZ6QaG0c3sTgIytLhNaz//QRxoILJ0Y8PrPi5vpwHJrLgy5uzB4ol70pRl4uVL5uXqC78xe
eoSScClYTMn8DJiD8A7ZXRrlB5w4SprVK10AsBP7C6okldFrAMAZgChUzdLYQaBXkKtXWeQOzrOT
ZGWq/Wj4jl5FqOZvmM3EGjGR12mknrOHVKjxdxQCD1IIBbTdVOPEfxhRHxl8KwNWaB4wQDqxLNc+
knDXrUH7/RdMBkL+IHCajLesk/W28SZdAxe5CGIDBet+DZ8j5x/hgc0roQa1V6x6yz26HP/IA0hJ
vUCCxBld96Kif70mDct0NN5DD19bmSG5ufREH/8kee0jhkxW8QzvLwwUW3cEPOnzXiQcLu9E5xUQ
n+w69VwJPZ6DTrUqktHsCLtZoQuBsuZPYWV7mcJ+Op4f8LFhrJoK/2kf4IhaakaZUf8Bvrk+ZB+B
wN0mJK02CugObum7E0Uvr5vTW8C8s9OAze0+WM+TAMIH7hlkd3OE9FmvuKmhjV1Kkmrr5YewI+DX
ccMubAPXQnkWBpLjQ7bMmj+V93/AgHpFpgId+9vySzYtcRQ3zP+7Kzd9Deue/lbZoGuJgWFtSRMl
IezXvUQ+BUJ4MHFSmK/javkzdyuCKkaRNpm3wUdN5aJS1sEpSyUa+sb9DLCuHeUe0svThoDF6Ylw
aKlVc2/MnGyfI6X40NwkUJ7Yc10ca+zgZC4FBDABr5/7LX7v9Ikb/Ygms+8qWpw+EJp8xMYbj+XY
abCADwymsNh6UG+KQrR1IbqS+j/y1Ssrf/PIP5muwF0CCQ752bGXNLbm22szM4fF8AQ/6qd7l30i
cFux7AEB8q27iEgMU/HPhcmPyC92mye1Ov/fwCMDkSeo7ZxOIz50YpPubTJ5lZ6M9B+RnvD/0Ybk
K9MPP7urMbats4k37BPeQxMdlsSjP3ooq7OOqlzxDpmRFRJyVzN/4OZrWVpL/O4SxBriD6A4w+OV
/EK3Ti+pia93G+v4VySun1eBhArLqniSdDVvoMM/sRYw5YDRqQpzs51yOPgMEp324gJJCteyVDep
hXLm2+wWAJb/mGzA6rqp9OVUv1yEyTA4wgeW64eIo3TNyOedErwEF4AZXXREIpG2ZhkneyQsKJ+6
AYoOb9wWtIEuKZLUiAHKKz46fV5842Yp2bysfczhPxF7Er7Pko38R6+wV1mo8Wjk7Zve9ijwykKv
9EM6P3ksI+BADmDELoM3mHcd98UWcCtiOzZ0QTCsST3m+WAckHSrYVpJ4Gt/EuMa3blUUHR8LxAS
XsP/FetEF/DlqwitXjbMixPh1yzBQRv1uW2XU1Y9BYag64gAeuhnRnWSvj2p7nnvqCmwonEzttld
/O5sv7JqlgHOQqpyLy52yrDt8vqhLRCk8BLb7q2AcQudasC+8Szllzune+tEUkhSyUW8+plfAZ/P
TrJ/surzJ7mpn74+GxAmWerfkxLIV/LqY6kTcJBB/em6I1xqW8EYAipwc2AZZ1WgHId+9SxPtBVI
uSKIVriBimr2XFnh5+M2l/iWDIFlx5hDzqgl6OHStylkPcJXxJ1idKC64vKhRPvqrmDeUuGuldt+
33mabG4KS2WghZrJPSs5W/7ia5UR3yRN43KSXM0dMWpfxTKOQkgT5jzkNFfMr1AQaRAcDk7HnLWO
WGXWUrMGu5XvaJMdfw+q18vgoK2+n8bhx4/OVm6dBvxt9qb1PF+JZ2STpQjkxo22nOHo9XeZk2wx
JF3aUW1UxaTPYFjn6BcHJc3mgf4PbHkzCLprzAyShm2kmlcT/KwwBd7X7AjuaWilFqZJs7dK8IZK
L4lDgsgK+pgb5QaRDb6t7XYpsCSbysh6wO97tcb2gh6r87uhMVlQXTvPliMtYgG1nSF1fJf/z0qN
xR3W2/p/xLkpwAT5U+HrSuxiJBy47btWBdfT2Qhri2LyUTxAB66/GoxrpzGj6KPbPNzA4A1h2r4h
anVRFYO70/m/xCx/42CpyfEoZPJQZR6U1YyU9PtGaW66PiAp4ll2aZmvZcyL8McgFbyCpTyC4yov
eZaZdDLstrhlv2eKg74LP87KebsfIZSrSMAemg3zW4owGFfMJMGrmWq6cZ3WQuathIF09jEqcJne
jwzDiC+xDcg4p1bvAxt2L0WcPkCwRU0aB5YOH9rRGmMHE9ZUXzVuTwYj64Yc57C2ONp1r0j++YV0
5lFL4P/8tslAIOg5FzVX7A10EMcyGe3EtM50Mb4zs+NMhogooschrFDB7Y+4DK4dy9aP29bODXQs
gNUHKWgrkWCDxWKZxrnAGaOb7f+cXAnxZSyMRORqppOPxtuabNWsb7EA66yNpWQLUjP96Q53/KdA
I9MAXIoNidSHtcipfecQbL5m4IqL4fmolVwYGjoYLUyM1pYMIJP/py75kh1a7ZGQsyCF7dnprD04
Elok7CeCIdHkYk8M6iSilfUW+tmlBspnqdYqMl+j/kGQU83aC80IHaKESZn1Fysc8hYThvb2k7pQ
Wa5OvvJhGI4xqiW/ENaFdBzYe2LM6pMQPY0SwJplI6Nhs3aTeGnwjs5mdN/ydAhA4NkcxPrA9Oti
ZMfZ4GsJUiRtiooVjDOLDvR68UX24e1SUFsK7kiBMdfE59uTQgBf5xPR5ojQ+1ZZVKGwyqlXfA4S
0/uDQKznQzoEiQfFWq0pedg0NL1ii8LI2AfVbhGmXv60t05qPM778/xH3ynZ6KKMd4qKY2WHDUMq
2fqrAxiy99xYc2LyfSgSOEQiWH4qZUim7phgkBcMQHS59KltKHonoPQB+tHcPgKIiZEVWAXYqW11
3mOge69oUAx2lST80IMOOAV3R2s5VIrxNITqKyi7P+2n3M1g8NULswnaftqu1ma3DHhhKV3sn1XU
Z088yJ04JjHVzpreVbeyPKkD6aCaGztZ3reBpb7Q+X84x+VkPbH+eixCn3LKoGXN1H3UfPf2u1mt
LnZ9kFSVDinrmrjXk2mW2m9c628JDt6zgQFV4xr6DJ4KueQcor6ZE0wF9VIWMfF/HSEtPW/XyzbL
Epo//Ji92pcdsZWwA/IOinFYoWJ3GN+2eIahcJIHb4bRXBT6YPZ/m+qlFblKH25jqL3GnQnm5zHg
WjXAPaBGTlMMnnmLwF96rlY+H32w2/P99usII/xyEZb8ROv5A+f2hnAio0zpLUB1Jw3HqP5YQ4u9
BJMghpQZ3wy3M0MZNEeGgkom29UMfgfUtb1uhxoSj2dQTbzz7wu3DfFGsYGvWLdEIGI4fz6eZMwI
QRCPedSPGMZCkQBL4XcjM+9DW6rQNA+8Dh9xmp8D/RKcXZWgO8rI7Rm//925XWQlGRMH8rdwSBuI
VStj3nztkZk0LXNOzTqnZqFz0tUcsn8tLJa06u3oM/yrmK8Fp+2jyl12/7valWDpJOz53nhthpdf
Ku19FRj+t2ulv+9jm50oEPK6yjZ57pvlu9ADgK4YScjLO1jikQu+e4hyrm5Ga4QH7fsQF9Z0xRb8
1xVegynwQRD1IMku7JWh5KCbiujF/KGrnHFt/tkjlFkHUIG55vOupRldnvB7BoQwz+hcPP9xSNHL
Go91r1NBck6m+qnczLVRgq2yf4AcFHBJJUi0918HBvLc6W1lrFUbZLl0n+V2ilscswoL5GrxQmIF
7FzJTxaDhJ5b1gUKdkFnUNBN3rIFpp172m2uLJR+6TUhNF8dJq7eUXXo1wCQ/jFnzD67tBKh1jy+
mP/To0bFQ7q0j9BjlFk27z8xjwaMXAARyqXvGyKJRLAIBTB13uu+mQ+jMRuA0Rj+ACEOx05AFmok
nKQ/+HggukLWmJfV4li+qPK/RebVfZ4GpXoOKuW8J68RAbH3/7MCREsGd6hL1AJdN+KNvAfkZEBg
UxtmkXtHT5hdS644X9yCf+DNuOdPI3YEMJFZBBVfNyu5/SS1NGo6hz29roP1ZXOtULn3y4dtCpKd
ffLGSR0c33iRxY/GFJu5SAwaPUQTw1IVOcsk6EyYNAF/4+/6GPt6lk1+LueyIwwthfQMyj6WfYIF
gQD+6kUVH/Ek7BZffUg7t6OYeC7xcnIolQf87pBjNCrDZh1q2m5gopr9AyJmHEIWiod3MovKrUTq
5U5+f3+KQlKW06w/uymYomluY/rtMCF3syyUfuFVGcU6hBTISLSzQiCiQSn+Rtfbw0+Pe5eO5YsG
Z0UvLwaiTKrXwVdSdlvlXkAw6KDOoOHZnwCxVCKCDvK8yrvLl0RXj/SDcnqTWMxeqEACUwFs8cly
2aDr1jnTFdMkBixzl/tIrZ5OaCa22sIoxrXOJ7oH/czgLvZjlrTH9xl9/ecADDzXPZScQIsg521v
Vyd0K5HrLbF43xr24X/QR+C14QO+GTVlIvomPvY/cmB+wLCdJHnkzF/wJwiviRcJivqtNRfVh9Lb
28m3YFN1VEclJfSUgKoK5pE1w6qnT089RzSDpgP2ucF57Jd9J1vUjDpEpC63nNntQnbx9m80UVzU
dy9uY5iwqvi5WQf/Zz/cvR9G14ZbGfuPphztFKrrptzDqWNesPHDtT9+kPynFNTcLRREtNlOlBS0
QrW8MEq/lM6IlXCSnH48SdfcG6FZ1eLWe8ZGmbnSrfewd/ex6G63rl84hB4Skq643y1qiKfrRCQC
UNQkjFUPwLP4f3KVrU25PmHKtPaC0A8oHbjpWZyy5MTwxa7d5TXayk2Vn35VlnjQedaVPsMlVQGM
QACC7CNw1L8TBjXEfbXkD6m5YtxqUn8WVpqW+lWbz/iULiuQxAiYHRPsmXJUMvSHyHR72x8MPB3m
GMc3k0jRRpIUmdDSLaeJWIepdlyUFCkexEi8UrBF85528xxO9IO+WXedfUckfGN0B7nePsHhapXS
pdPJCwwuQnyc3qROLdHN6wHgnCNE/MGOfUR3WoE3R6zDgb0RC1B2+JsjVR7uEPTNn8GLUs3W9JwP
BZI2EzncdYrAnPr8Ng+lepBH3a6BPPvBBK4PjPnFtJtfbdy7Udb8kT8KPx/o8ylsLcpV0YmJ1PoW
IFAYPtvL+xIojNrWOpeZsOBSFzYq4iQCBGeBayf9n46QooEqnv/uVYTN4boPEUuSLlRd81qmcuZ7
r6s6pZ853LVGdqcc+PQ2SjjCZoxJykH89hdwTLRmj6+NRgg2DK4aNSvAx3mWr2N+vzTWpZxeZAcp
Qyo9Mw3A4b0hBi5rGBwc52DiyBIA0iCaBEwVJn9oAu0bq4thQHpKB7iKqmbo6CTAOnn5OlO2chVn
te48OzxyZKEPjNesbjXI7cjVOWi0gdXc5+yKylg/UffD0DkPZrHbSTyWQA93viOLUJJup6YjOYP+
rCJOQ3cAi/v6mkYkQ7ZB0xNIr658gPCAWkM6aROhwOCDDsAmNzRhYxbRgz8ufwi1/XBbwe9Zv3V9
J5SbeV2V3alvClB5652tu4Vuo7yB9ANzG1JplFcP/f258aRbuTA8QkIkX4VzX0SXsLl6ekVDJdR8
Qmf6FwHMTfw3/m3RCBXE/6vs9gY/XtqCMUAuivtg6I2E2iDEhvxQpApx01vIoOqqdjHVPitB65FL
U0VooWkZDulrImn6Dmr6cIRQvnZr0cv6fAVTEpwbBUD8xd82djQUL4YPfZ7bS/MBjjQiqHIWGc7v
b95pGfun8Kzxa/H+EyctorrkWcL9s1LsZyPFMMoG7PBJDlzQIRJ8Be8RxBobofohVYMpcSHGXxhq
BKXTSpt7lt/D6iys8lHZR+wBDt7Gn4NMYvFHhnJH0wCob02xl4mLntm+yXrtx5SMxVSXwkfdxGOT
IK7+hyrSvw79TOzcf/B5pMVK0u7rzy7Rz6d3SQFyOJLSu1clmYn0mWF5CHDcvE07jVR7mSok/uqo
TBQLeW6qP7LBPYqgOfqwYbCZBi7nZwUBxqakg7tm62tL1qw5j3PXyWJHfnRuicDHigO7aJraGa2f
TmxBQ81NJjmsgKLoMTjHX/KlgCOPM1+x3FwFq6mZ9vEaMA68XlekC6c906Dpd+AT9d8ag2fbtlaq
BhyVUTwmwd+Po/r+oAGJdVqgJDnaHt+4OagU8nl4usEsg7L3GfTIZIM5cNlKkE/AEg/YNmgCRgPD
vhNSXq3S92ABJHBXOz9YfBEKQO1YWeD9ADCKcKHbZqo5LRmsQpAeoaPL+0A4V+c6+QGhdENCvQe7
kXvsvxZ0+9U793XuF+FSsKjEHxBwYjhtBCWbpSneQfMNsvHs95HvDbWAEu4IqfYk030qcngPNt9N
aT0RlOBGCsBT2PMisUkpZbQWRyB3cn9IJVjglIwbRfTEjj6CGQ73h3QPMK8wCF4v6JPd4iQHTl9+
WOKpCQmE/wQZBy3H7yA0a9Ym00gmpD4hEAF/JZdNtl1rRROtl/yV5dv0f3+lnbyLT29sAsPhmUq5
UgjT4wnmDyEJNINYSCHTWOT4itf1Uj6J6nEeA4TEe3PNuoVZZepBBcmQbjdqwS1A7k4b+E6LTk3F
0K+84zvEBmCYFK651BWk803APfFJb/FBdrC4xihiIfb65+xQi3OSX0bRiP0V2F6EKBYCnxCZFAG0
m/zfKwaU2tD9FqXtwBGKxUreve2mufuI+0Hcx4mOUSh5/RHOCqmz/PSWxuXgu9U6bZQUMoI1m1Vo
gUhTUHYFB2sPg0w4j7grfkZCi91ckWdxMa9GWpI80mqGH3v0hab8yu9O9GwX1mRZ61Jgj7JmORcA
j8OQXuV37NhCKapGr6r2s4+fqQOS10EvsnMgqdXxdQKecpZDae5eTuwjRuNBfQX6Asp135GbgfwY
nfbCGSDvXKoxDmMg87snhQ1vHL2TJp2QjoSwlwDIhRr9+BO3oKI6zaQ8/sz2fPxoQJJ4UkSKIVUo
cDnZVA8cM18cs0FSaW8icWf3wiAlu60gJ68jSltwmuIiQDZf38XH5xrIng3XmqYicYOi4gjjuO7Z
v29oekZlUNNLH9TXFHbvCl0meRn6yhfeiVQaHb4sTCVe1nf5Lc1f552kOaxLmXJYDFTSmwIBMJes
QRp93NCXL8fPWTnP8WuYgZEacruPWhIGLjzzzr999H7bO2dXoHurpWKISESxiE8BIwev5H1kMqUX
gQ4E5HPlafTJlnshi3pAUP4dybLyBZijiG+hCzLdjETnKxojxBE61/tknE5QzGz2M4jmo7FKoqGI
vXSUIBXka1rzLWhIg9M0sQMvT68n01v0XIXU1dC9zs94597HyPBloUOheJT9Mg3RvHE2Kum+My8o
ZCgocTLUA34g1ur6NL2xV+qA+8ek1hXWF7UclREETf2ao/0tjQlSlWkfDUtvzrH3BOWPsuM8n3jA
st90BUJU4Bo+NN2sfn82iUeQa0Zgg2GHaxRP1HOtf7FB66D/lg4cBEIWB/+zm4owfVlZf3PyZiY+
uPQsQ5ZHwfe/hVLbCOCSiGu35a1VLFHr/p+xOIqtMb7Zjg3s4Yaw5/K1fcTZhnkkUzAQkHjz1erW
T8GR764/q1kJe3RGuwEQkoXEhGYtTyDy240U7SOAI/IhC66yQz9mFHG3P0KVNzHMjC7+J/am1S72
GWwIRdmM89LxBEt+PXXjXVvRhb2aVT46ccLJyz7tzXY3V+xH5DCF5azz1ZVftxbJo0PAk/u84y3j
ecIob2KvEIHAvA2bXacMRnd96UKXWVBBo8qPRApT/WNasxsxlm8naFCNhqjVvwhcFTGpSCd1q8pV
22d5aIKMFbHIPvQSSxoZm0NTNAhe8N5qBF5D6aCLikOBMBEDLNkNk3KBOcFEI8eLnFa0GeLFNq20
gjzeQR+sXWpn0LxfAgy0UCqyHXVKc/+t6rWn5Y/ibI9kPUAyTEbCj72nklXLyW10BHqzeRvUMitn
NFHTozzze45XGKvupQ9RvzCMDL96B6h+DYG3Ba2A5+zzwxHmKvZqM/78qZn7uEsmioEM+Jva418H
8G8rn49p6oISG5/FCdlmQT4oYr1X3Gc1GUlRXKJavU/hV49cYddaR+VhrAP3ceb5ZxfpwT6b2TVS
PgElUhlPoqXwGwAhvSbSG5lpMGLNSN/aah4BAtVZ15IjRt/QXhQ7Zn5tygh/BjtMR5MoHNDS/4vd
nD5cWju0voX43h8qgRphTVM0XPy1B2qxM9FderjnUeWaNBbGEfHrqr1YxCz/WvvNQywgEOWb6FZi
i1izXeacooRNkFNwkLMJbjKGtXW+f96okrCvbWZaUtu4tpObugzRmrRTIk4ZoOwcACjh9P5WqFe2
LeNGNWMjonLuPv32bTO4pqxBrbusTbNfbmG+KSGaD/0v1EtIopcjD7uk0tpbyHiHVFHHmkwRLQd2
OTDKoNtPqiEVRPuJrPF+CkvccqWdkDNt9vdSlMvN1UO20b+twKYhfjmM0rLVuT1vRIbM+YUmvOsB
ZXmeNoLDepte7ckRR91skqU50KbSLSM1+Ge7+ITkuV65gFrNvMX4OIZ3S8th7zgjISKhBZ+Cx/lC
pPPBKD/DkMeD+05PzGSyycm9NAyJqYkLvc5RiiN9+lMEGm11ab5rbhrk5TR5q6r02GwEgD1VEc4x
akbo4ey7SAWU1cO7oEe2tmJVBpbP07XNnlknNlHBUVTfSenhPezI6FyFQubJJF60IRPJ/vqXBDWc
qLRLL471CZiJahNKPplOZVVcOJD6o82VhFmIsQwdM5rVoV2z+LswAx1niiNhVtl3KK9ng2a9hmFY
XmbQ+8bxcjtOCdVWjTUyYWhx8rpqMPQ9gyQ+d0D644WqEdfF62lWoGBo/RKNm9bmgUHxPTCtM1ks
WCCMU0SFBzTdCKWokyw5iCRP23ICunswLobX7XgcdjhvO+dJaVG4yDAbTo5ba2xnJALdR8ZFyTG3
XAJDJEmvOCJwIuLghA16GdWK/At49EVpc+TJpj1rZ4w9RkHDq9uF3XBwkMdU+PCziSucTkZvETMG
uFhl+Im4fieV0MumV4rgWWE+ryqXIaA+EPkA96XkbLWyYOpWXMvAZbAQYD1XHtyjm4BO2XruewWq
FL+Z7din9sGtAgDIRNNqhSgVxklDQkvUhxsSnh423KlUbfMxgfiaLw8ognf0WR6sHJMRuDVmB957
vaY+J3774peuMcbZzGaeks2/r8ZDTJrLhkNbeDIkXSEn59HdfOXaXLKLe7jrEMjdsGVAGk5bLNd6
TNwkW0OZTAEU/tsQYiKQ2jwFo3946TA11yGmry28g+InTKOeTobl3vZBDrnkFJ6fJbmflclPYjfk
1yhx64b8oKqH4MCvFlLfAzF4U/xSNKaaDNUJZtdfZWo0qHSG2kOoS15298oRvUEJvP40OBdQNHno
RKFJ0Wjeps61Hd0ejkzayvleSboE/JSIKjXFja5pPw3Dk926P7tA808Ky/Bhx74TtN6WEo+IgSzF
R3ADVZ347HJgOTYNKTBUfO8NBLFTcnupvu8sn3VFMpKLHV8EFd4tL+Kk8GZb1eTeQ5AfCSOw8Ofm
Szb5gmmTZDHssjO/AdwucXORENgEgALjTa8z6mL19HPHeGda7SnrLkmmuiUU+/xsFUDL7/4UvNp6
5Q+rWDnGLtNW1jquuhBCmS3G8DiPktakupXjTQ9za/hHXIC5sx4CzLqREgi6v8ZNfMBx+uJNzrfD
UqaU3PKJnIO+aKCD5tYoUYmHG+7dudXYQvgdKDIswPlui417XF5641EErIYwc+6R8nMZ15bSFOUk
SmuT3bmN3UVMGSWW433qqT74MXLzxaMg7DFfiPJy6156WSwpPm0EWrup6AqE1uKeI5dXmvpJSKUT
h2KRR42YnHvoF7Lg5jSH07IZnk2dcC+8U3epOkAeqAuO6XYpHi4L8ut2PukOUXA2NEsqLaNypJ3+
oZiWSY7i8nWuI+nlZXC5RpIMlrbuxeqbq1D1lm2M7CV/J6SridyxbMYmjrZNcC/LvBP9cdKbt7w/
AEi6/CZTwToG0iOHlvDvREJiR4VNHjhVm508igrluFI/HcPpHF0TyDrNRCVvzkYxoXlHllVgUYtg
G3LUaOrDcA3FNNi5suo8IhULFmlyhPWfGTCDND9dsO6xBcWuNKrLPyV4NoZnCfhINQHUBl/NC+U9
i1XWzzSSsHKO4U8WFUVBLvcecrhYmBzkEd5rBuyh2BrUhAGL2hey4YtEKTvJP5j6APbcchlo4dFD
JBeJ7DxCyDAXmGp564ycs6qfHWjLWTF06Mq+UdhA0LOG9mnUO6vnoIqWdbewJEEI3gqIBjNkrll2
TQKKnxdxbPpt+W2t+AyWgOdckgdOavMl5M4YcY4gjVMrkAneua5BiSL8JF0O2gVZix+cMeh3pWnX
UDBwM+qfjIr33wIx0ynVJK1E/Re1L3sFEtFKDzy1XbzpEMCaFG5B2IdWfrY4n+cY+L0qIkbFttNy
Ilib4xsxqFffat11OpCRxobIOhtSeDfZV5baXwqfadAhyTXAfhTX8vwDRF/WHc0aiaQdsdtlqqr9
6A6mLaKtVLwcUiMtY/3yD70c+kjQHkzc5ZyznQNYDWwIW1ZxJgY5tD3sLD9vdgjxYiluqbsF4lBZ
ZALb/9O8IbQ8CqEK9qV/+lZSI6ErKu9GYswoSCPMqZjcyKP7oSJpPi2EcZmuSQ5qgKOpVCfBaNzN
j+yrnZ+L6es/Pbr2hK/TRSIP+IoDeP6g6hluHEgIpkJPij4uQ1u71VjgJhsaJ4il6422pAphKwlP
VOLlO/PNPcwIarsZl6zGXrTVCGzQXqROxqbinWeIZ0DFgy9YIyT6f8p6Ws/482TAgGwFbUj1lr4W
wqrRVWo9xzObl+FbohgHxQrauB7XYQbZECDRzmvdKdu9XliINFzMjwG4JhjFa4ZnqsZOyqGaIiPy
a7eLlST6hvJIaD8uYaYujTT66ZwO2b4KJMwL7yyDdewmZB7AJt0O27WKjQXp2NVdQKhdc/HaSOOI
bdnu275wwV813pE3tgwGePVywm0iMiLqMfVhjopPMGReqIXAvAqQSuQkYI7ja0v1ODIuxpUPlJMA
rHVBCIF0eqlMkv4/dxCfPjfBCOOIQ16bnzjvtIsC4A9jmr8FIIV/S8IiCVAMkepXV+lBm6Xd+stu
dsBuyd6v4hnYAO8g4ry5IdyB8CbU54gxE0R/r25/F/z/8NgDnshEsDWJcMQOUb6pZEgvjBj2i2NX
oQYdDG3WXY8SesNCPKHtpp9Pz/BbPkxN8hbbWwmN5VOOpt/7VAS6i+msmvpEOsGtpWCqwxtPe0jE
jTzP29ytZ1BxS6kpFLQmX3iypoXUx8fSuSqq+m+QDHGhGpWMpzsD8IKyZeT8jZ4QOlNHa/4+w4Je
QA51WC/8W7pZa3iifnuzRGKN+gvfip5hI+hUgjdK5JG/Og1bYpGiWeo8Gs/mbi4ZkQO0vsyy3cQp
C9Yvzse+cSVS37h2/ihUYHhyBsQCgTNgfg8Xv28pc2Zlz+bMO8uKcPqo7Zj3DQf+JAKErD9DYvQe
lKxDqyv10tH3Ls2ydH++x6zurnC2PNBgwut1lMdGGxPkP0Fyn/L+vElMSNkxzMWxLiSUU43Y0kdB
+ijsX6k3ubDOsABpNRz2tLESMQ5M45E8pEufUT9oCWcyhkk+2YJnUIsyU9aSnKp60HsYewa+prpg
BrT5ao0H74Mq0c0gmqOMcVrlPBbrSFvB+MK8dwGFsQCCaIoz//xTNJcmGs6lgDbeu15EzZMqliHJ
4LqDpPpvn11gECWPZj6gyhYLRyQiMNR9R+vUmukzz96wab4tdcC1v6bq71jmeyaDwmL7yLdbLzIu
DgawALfwMzWlXqlAaMFC4JowjRJpZesm49rr1TKVz/TscyY/PLPN4Kxq4KGHDqJCL5jlTApaCBwq
l8t7C0fFdFGk/+0sAODXMYpB83uljGQfUwnZGBd/iPRyurK5A02pEkRCpEjgBIj/wXLdIm8CKmCl
o5gksDRhJGjPM41aXGoJYKH9tFGxzdV6MzsBSNzebKxRO8x9t0tImNUYonZ03CEw2Y7M1+70kLrM
ZQ+jbIJNSrxSQTr8chRtprvaG5uCPeVQMnYgVGYBpLm1nUoUikv/F4ipFBovVtRexb1iK7wys8DU
ipU1Tsy4qJxje4uErUKnUnuxcMg9bYKsrgJ9rwuRhmcRcZqMjj6wvvgOXAepHHngNpJulz/PH1vp
LtteupTTTLtqQGWKBIaUd4JS9XRVOyycs5hFhEaCP9sYa5sfRmts7KaRxSe07z/nWVKp1w94EtIA
oHgcsOUsjCDXUO/0Qu/3dF2f/7eclAwigzndtuKLTm3eXNUIDD1YICWU1wwwDHjFv7xwgYZ1m5/5
57AfoesrOXL7vq5dS6o4vMvU2QkTm0hmAmr74iurgxQlOK/feRkuETE57pgJNLutRVEIKSerF3hm
FT21Vtgy5Qt4pFR5dNK1lg8FJy+Y/OMCGvK/Ku/lgmYpeU3f/qItJ1XL6khhOXc9Zq9YAGZxVPZC
sTWA1IXLu0Lmd7Lhm4AZ4BtTBy13Eu1KtKfoQWTuooL/QHF8aU+s1Mw9VLl3/wfBJWeGX04t0xh9
6wMi60bWwJD5ep2OEG4UKZxk+8sMRWYpv3mct3NdieNO21JBos8hzBqJGhv9SFIj7pp3cCRuhzjL
qBWQ8gcSwp0j+a77sxHK7gOnudKGBaNdIGjrLkOBf5SlemAsiw17qFN5CiOyJjJSRvGtocOb0rRh
oWLW7WFvUksQ+2PDZEHXJTyFfC+n75xr6oxrYfMQezH8RhoZOs7RrXw+m9RoiIf+1PaWFB+odA6O
U1fw3KGLsisEbPNtWj22vYK6eFD4M0qOoSHd7HxC34HsM35Dq6L9oFtIVL35uBv1pwpueVbF44XK
TeUqjNkO6aty/MvEcLWVq+h0c9gdGAhZ0u1xvtPjEGZmHEJmz6hU9717KYQVW2rLGRu3ofnLDMZ8
B9Tw7ZBHwalqMd/2/n9wW5KYEqzelZqNxyLJcQH2h5SUnR8Ju0Bu9dpPMegJMoMx4NPCLxsiPBrW
lJcbjloI95edWVgRCn7TVqyZXp02hN6GE47Wdq8eKBYIuUxlpA1BU6gfqId0xQRuoTJILoCf7ATu
uyFaKh4RS+MFvvR+jBJU7nrOv58oUQx8yopX4GQqqE22MEHk5ZO5BbBx63iaDKIOQA1HngqKisA/
XAGDZx8/8p/k/0jvNdYp+WKR8rDmvVFjolv6bPhJuxF56FdJAY/F5+JQozOQ1ngd3xdMR/qxS2LE
2fbj+tBIr69BgwBKlxoE1qaALV+6CvFncKXDdwJpyahIG46AfwiLd4A4RBRQCaIR1jeF3RNFrDLO
INtXuyGHq87r+bYQRPB/8B/EF0vNZCv0R47aLfbNh4xtjKq3xxF0ukzFieNt3q1JGyP6bJuveICB
2e+4Xg9DaQcgZs2vbogP2Zkyz5HWph+YBfYuQi8ulXrFYbSVYTC/QJM2L8dZItn3q9uSayDohq4S
wagMzQpxtAkMWaTGmj/d1vTh0kR6ryE5wDNJivPzOF/yzyxfhrYr88KhieVPuSciMtRMf5/O/qTS
TXN3+QlMV0NyyR+AV01HSzRf6fbNmu3R/ooBqw/hn0bcaCGau3MWnap9DQekVRkr3UgXs9QOFSvU
z96ywd9BLy4WQKO8vBrPaToAvu+5+2LU+J9oN00Pl7TKNHfQK5Wp/yYvm6bYbOV457yyHitnwM4/
KxHwxKwL6SlM9wJ3EMGLwZIk/uAYhn4ldi3SZNgghrtxJGx9UMUuAt1bm/EHbSySNJyZmBrJr5Zi
61hBhnMGMcgp26fMZa6NOjlU9+oOi0YHWwtp9F8nSMn5351Kng+xqQVWR/U/LgGAJALrHTDvfUBC
AygMndwFQ3j7ZAKBEpbYrcQ2ZQjZnP29Jxc5UFxYa+qNzget0kdrVdDKZD0yqawrOPWS6yT4dlLL
qq1qhV8wzMYNmpwlyAcAOuqoeWG8VzIyA/e897YIQw5CmGiuZsTbUhjtcJ4quxWLBPeeipV3mKyb
yoe3AEWLP5EowlAlgh6mLVuWqigOqja0gjSX6kTjy1WWtpL1NCOT16sceo8mdF+khA7yiNLo0qgn
HUDX5cvxR9bPBmoRFXpwvP0NzCVkrqhHKOdXKn+ev3FY4tI5LpjKzDpP0P8GeG6MqBxSqui7l4wk
WpGmwa1PccKZSKqf7MB0bxAdU0I+hn8+KArgFmP+qU6oejOAlvYFigSG05rtUFiVunXGle8f/sXB
QwPZGLy40Om5Aq10nAHS4gSxFv0qS88DMGMfqjxyyzy3MF6KNBIDlBivlriUqOGeDHUZeWHwY9cW
vtUW9x64U+mGioCntOSXlxe2YoTdR4dpgy0BOwHL6nmMGsSENfxtg6jeEp67DgXFE8y+bv2vEQg0
YeSHsPVrcP04mnWruCjUiMOwjtPaGbVXI6Ov1PC2TDmeFxsszZoldLkrHpMtHy8dsjv8gQgNLQ5F
UAvayaC57heYfVT4lHnTmoGdYXWAqNCm5+svuVjZSIY9vCMBure4g9txjsRYcaLwrBbFG/lvv/rr
fzFltk9SEL1HNviprhDP6HxFt+WnEk6aCdo3ZGNcw0c9+lStHgco7duEZeGqgw+XDsEgaq1hwEqP
Knf+HbEaglFPkwwQQ+uhY12vNQBN+D1gJuwjgcX1wnnISMmnVO3Ng5iyxbJaU4jWguC10KHojuPb
0nDJ+Odr2/fBbz7XpypW74G7YZnStb8/wZayjSq0OR8+Q57jcIFxf6NxEv6Q9dSgXARsOZQJjyLc
uRwHECW84F8AUt0Uo2aUq0+30NYl9sX+prTJ/jkMv9Dc30xeIEiM20RBb2AgVMYIcLUgucj55UCb
U1u97lg6+07auPPq2Y3hCsWZljL+LEw5flzq/KvOpqhS3GXBq9oZLZpDez+sp56L2xqj4I/XNFxc
2lBhEsLJZ8ksZTtk0uRpFcRZbuWt9MmiMTgZpyNfX0bsnYVW2nOT3IudUSUrLtfB+0muHbWvtQ51
zmZf26Uu5MszVjnlaSgxJTcJwJ89hjKEreEJd4BnhqLZMgwHSzzQTLG4gHRkBOEbJiplgCcrz/9/
4cf+nVRsrUBvnJ921rqr9Hyyh7lMkzYfOdy6AHbzo5uu2hFXfhbRZZQQTSRhJW62GF8zLldocJoU
wKlZUpNTuheSoH01mgxvYIcQyjdAb3DmwEtz+K9nhbHF4QaGyoXZDS11yKmAG2wL1mTtsFWtwvHg
Dw/Mm3Fy0gDyK+UK3gwW5fa9QoeaMHBYxx2xAcv47KEMZ2glkPHsryrNWdUp8Xghjg0JZ5oioMsv
YQMP0c/Zd85AU9u22841eRqUXQiAQjD7xarYzkGpuveEZPN2b5aKSaLRTzkOtTOQJhhoweA3r/1P
/gm+Yq8qCQE7C1+ndMD/VN6wnCGQZ+YAhI7a0c57Xgt0y0d+Ow13l5jZgfHgFLp/LtLppyXMdEnP
5xKufUZWbBQ0X9+mYNuEo8wKL3JjuRreo6vy+1v3lQGsyQjAmgGywRg9P61jJOST/I/dQSyOk+0l
g4FkF9THBKUHsgHPHkLbLT6XEU05sFuA8+/6sjKY58taJRiB5bLWQFZ+fZUBmDfG2MtPhe70TKH5
Jw89SUcSslE6vQdusXkbL4rHp7Vl0YKsSZRPIp5gY4dN1hjZtUPlk6G8UyIedv38X8qeESOxrcag
x5312jLMwiSiwUVtIFRH+Fl1FGQXxLgvQS7+XTl5RhhKoP3C8KLLWiDqFyAy2+EN65rvg3+FRt6m
LoNlVFv0LV1QVDZMLSkSX2IPVHfU7N4yZTYhrMAUVlrx42+0vSu3YkqYDk7jax69ZWZ612a9PdeT
KNP/MS0ppU0F/H/qABnrYudn70qcjCPq9JtsHUNvqCSEdYzZuANpCJ2+Nk+9hP9E/suNCWToHfJa
XN4GfSwlVz39pcQok9KzIefmlAzLmTfLpo4rlWvtZUOnRQbQSRwlPewqlAdKuM/WPZ3GYMZTWCh9
WZ4VWvv/0X5e8cmQwW+Y2FduGPb60Ax0JxmcAY793X2JMN7nUAw2HevJiYJVEKwm/hBnD0Tj1jOS
tx5e1KDKIv0JIZmn5/x71iimKUR3H9jj0yMGfvWJ5u58gsQsIna9XzP0xrQKEJY+mbX+4bzMyP1j
ja4Jaen8GGl0rwGPybuUmavcw8/meebIfPSa9nFynMzak+66TU8mRqsQj2+K3TG9IpKzftsUOfp1
9H+85ikbWQvnuALypJZ16pKdQIG8Y3KpsIwb6YQIxon0ZJU7CKdke5QIgKk5XxigR9O0dilFecPd
+n7g9JmqI1mNc2cO3WacBj8TIJA3R46RricDi8SzcPBTbJT2wIw9WMDcFgAzbnXl1hnsIsh+iCvk
KiEuZaJzQ3Mjce2JKqp3wQPDOtAwAV4wTWZu5BuzzLDHaP/IpHmoId5uvgTdBxSNU1S5W2fPHmnt
mtzjvl2Ajuy22iW3Wvxo1dyqzI9lyQhVZhtxLwyUhkqvA5CRhk7THK84EtIoQtFRD67BcvlS0HjA
zGiaVhD+Jq4MEKYvbqUqHGoTyrn9d8vOU/2a+65VrIRn8/EpN5YZ4y6pnECFj4jh+sHJMbMFPLW7
4eHz681U8e1qVJNyMrwRdvPGTkfKlqaToDC3WR7nCzwR2pMFkMtLSJSV1J9lfQR/9sAUhmTrtpw6
vHadoGnInL3fEB5MZ/wRjU4+w4e7dQU2WTdrTxlXUxC9L6g9ogzPyFNsGhvr6oDni9yTcPru0Azz
YAr7uKpeleVprkmKOalMzOSXy8zwUAwfPPJ2E1N9n0t7i2CoslzPYtBk73duxKYZ/oESgnkBI+yH
X/nwZswr8sBhV9JI5gFce+2+7b/MarcBHNkXsupkTUijXyBEQHHRRBnYACnk0AsUNwUWDjgGyHWE
TO06/IsujF8HjE5WjEcsbqZzHcBEsmCgh3HjKmw3AYdHVcw4e9I2TF7RQaOudR9QqeO6Pe+9jLfk
tdhdBtX7EoAD05pPGsyHltbxF56nJjaOzJ3P60sgNzMISoOeTPljMlbwfwLVP3ph9vTmUJOTyTyV
y0EYgABk4Ld3dmT6CTIiQZNUD7PVQdJlidhK/uVsiYVZtoAIzcu7o9RDO2fwLCUamAG8t9wLAmMR
pZXJl/Z1RVY7clsJttW8HzSx5sy8a/clz9ogaEEgcBSDDkJqy9Dm9MKywPgPnwKHBDZkyQF0NTSM
n9k+NJlONqhYCWezcBxIvpkG/rFefWy4lpQ9FC+tq4s7VVXdtIrn3Zltcje4GhomOtKUnnUqWPc0
KwplPetcZfJj+/O8pl8nJjS29GACTK47ZBaejKzbGB4W/IqYe9nOs3YZU0xCHGuAu5goX4XOYaz8
+otDBLfZrVsS4HDwdwg1IsotBP2oaTMGqg9L9YSW1RZn7gmYU7XjRxRM7JIRCk9gvIcbEPXfh0Iw
XCzv2gMm6UMcvZIsleyvxeR2iDQsfQ/emw8C5T5fhVf95/szNyLRVfUfAEwVGnzGDGEw9WMCSibv
HGh21xSQjp8cavKoAAm5GEiT7eTdxE1Vtdh/BnpRayI5Dru2Oo0x/3czuVrakMZIhAbGGeSaR28b
cLphWkqR3H4QgECeuxylS6lDONUgEfew8+Vr05A5qQ0zXE1txACKwUnTvPqOfCsFOLQNO1PYZ9nA
Yq8ZC20ipyYV+c2Fuscbasz5XFY7SHgM/WkSJdOOAMSdgqn09l1U+3ZfwtUJrmi4dhx7+9GS6v/J
uKKvEWq7zybvtoisRlA4d0MWrICGr7vCcAB0GCPaJWr1zntYLQTXSZ3SRTLRiAC7S7VGXrpzFMXO
Pbte3rSqyQbIwtkUIrDqiRobUYlHRm1hfrtxLC1HdIfWW7KAm5OBmfgQvn5cWYYC5x5dQZZ2CKZE
LXXf03UOsRuAu50iFXGOhUwKBAPQpOmu0J0MbXAtFq5r7rcdMDQ6DvClggwDNokU6IDSWJ8lZWCX
cT1TaeKTLl50E/jWJgq4UiKkr+NHuzBSywhRqS4cZzPnOUfHULvmNRzO3FzVJXVuUGPdSpc6vAMm
ta8yQEfncBxKaFACPiq8rUiFw6nACwNeacR/jCVSKGmlV5mZ2dwG0A2fPSQUe/tZ4DmPoh/Kc2Rz
I1Xm39wstvP8R9CNTUMV6fmY5bof6WtWzx4OBC070xVk/fNqIA5s6gy0ySeKW+zc8uIysmQw2CwO
XvWYbDu87X8BgWe3Bo0t0JKGyyMgJ12HZQq/92VkR38bK5CjxS43YyC1ZMOK5ebwGXx0N9ghzQ0G
EIWNEg8kWyMmRQlKjr0eXrvU3719Gjvqn+bxCxhEMXpwuuGAI8rwPG44iIzJoErkTlLt35a7J4kR
54y/HDE8kZ9C1wzyIic+bZUg04HjZA8/ybhhjXJws7CHR4uVgoLHYi83ZOot8ka7yH+U+ezZ9V3G
sLfdsTV1Rp+3sF9BFjlNM7fdzrawZrBxYbHv8lHnIXGeGe/ndRyHezFUSSVQ0UiiD5Q19oHSxItu
HlomINmmbR4Z97fLfi8WJYtUvUnwp6UnGZHEQayXlPxMMeGGP7j1r7FkFeOFMqObBPkl3WUCEizo
HHezCGSJiIq7BfKLJ7LSqP0ch0Ln5UrGg51GW3tF3nFdneMm+y7PCKUP3gIkwHDceN1ED7Lo1xjj
R4Qpw77dEWqv3gtRKZF/ldzErVA5xX3nczP2nJ9EMngoj/9ddRXkSqVKi8N5puBwR9lOwOlB4DwY
UVOBmFrOS0aSMpgaHTxAdu/9jyb56qS8SfuBXfPLtAjXNRK/7eyxB22pZPy/ujOtz+jAhaVxU4Ol
wfGvCOE0ob4GHaF+wzPbOB8Jh1xDPTF0OUpghi92L3bzfXEu6PvZuPTtPu25PuVeH5UbcXWXXvPE
lFdem8rMbpY1c0DynKfWHr58GMHrjY79nrSfK/fyF+lH8bAimVyZcCzIdO+1CCCbBsrOHKnpLu29
vgsXFO3eolZ2Fmds54KaTv8lX6xDEjQSPF9Bpg+/urNs4dxVaHaTjEg8OyCBVZ92FMSQ4IhGHLMx
jMABo8qLNhsBORt5GE4Jf69rwCYX5XRC7HMu0dPwcVnNZW7/4Cg7EL1fl+6s7UczGHghHuCGFNHM
4Zu2qVzg3dhsptKNj6+QmZsqEh32ylfLLi1UNhmPBsU1qkwArCDZIJtWxh4EHH4YW4POIbT/o+f1
fQMmcl3vVfdn5ANynnccmJl323YTi00keTsR+GgxgqGxtb93pwfdQTmPmSmQIk4BH0FYb6XVdS3e
l5WuxnEsJgLfVxZsum1K18sdz32tfi+oZ5YeTAKcrkZlJImCx5V+tcq+Noo25eZE3ZN249OCLuYm
O08IJcU+NXYgdZ4rKIqu0FQYoFuHc03v0WP/u1cgIWibQse2536nxYoSECBxDtn0sRd5xKYhvLXu
A6wsQagcV3cgl8XBzmhAhLbXSfDtr6eN6ax75VI4ej/79CbXgX8MhiL80aiJN+HARGGBfWJ4zwBg
bMfL4GB0zGq/jNAFLq1u083tDtUVF3I1aNabGHpUA0BpbEKnbOj+SqB43gFr5/w3DAKUCp7W0VMB
gu88U6qs0f+HeRNGMm2y0doAoi3d4o+Pr8MEtouxQ2ofkRZUXcUAKhSrXvwGiGOWWkSBZChFNPLI
3RfO6B+UrccjAosR9RS41vIQDpkXuGn7ph6S4xB1Gs0sbAysy2HIzizGy0oBQ8XrPv7t7+5jvZ+x
F4Rfq7Ifw8NfCze+w9iorc8Y1eDrXBWkhA/H+SJEKAlJ4eRC0RkBdrBVk9/4ayvP0lSjUl5NXs7m
OtcKV9j9yfa7b07t+qhOLc2h/YX2RdcNMawT7brNZZDqe9tzUs5da0ALQxJ9crPpBNSgoZnXzfQ0
jcYZSLfqMbeJSV8Xtrdlqr2kgZWgMro3zkPY0YBg23LoMOXahCpZKkYwQgWce9p8j6zvkIbnJEaT
uc6jLBa6uzySDUd8jH7OGAbeKw8vvt76uWDFtCnv5ohtE5B0U1qhQR/prnAhZ9delzDFehA9xvAX
UWE8a70VbV+BlqnRCS3TKNywBHsV4G1FqueQYp5CCcJYfACg6YReQ1XhnJhhgad8DXnJ7Fx+TycO
bLAQ8FWX3NbFF4CbZnahleIiPR+A3Q0/KWftxiGTPMkW8Lct1KgEcKjKJwvf/HXV1nBDUV+ub3Fc
3qNqBtHcdfSk5WPpYeSSgePpdyIKqg9K+OCA9Ik3WRW1JQ6hNtdgqLub7dP7o9lz0THwRwM9moJ1
VXQP+gjNZ8fdJHsP62qMgS2ps6miRYUpi+UddRnpnMvqTqT+CdCQS8QAC5US1Rnzne5BQVneQ3+M
CW0EcUA2dRRXIgLwOk+wlnwtMnpvCxRSIEhjAR2WzGQ5qhskrQRizkhlcdxPoH7oX4+z7wFo+cqB
YXf7Cv19UBjY/OK22jCYUuP3Tv6lXY0uKBhDjHMi56SP9EGe3gpS0y+otuwPER2bgaX8awsnPgAQ
vhHCwlwlqSVoX2sJ8wWQJWrKpz7JlOlzOZjtHeaJjSgQrRYjdLtzbNZFGRoGKkeQ0m8enMMHGqLW
yz/UN5G0uB+oAZz2uiWBN/fEh4huEql9EqI8VeVXhKE7AecBThljnXttqRrUrjtHOL3a29v/y6NQ
6d5CK5mrjEck6/nFmV9WkbA9IudSG7hiizFlD6fdXeNgY0k9daVu0/UAtGskaeaygnwKSceJHYnb
b+8DhlU+F/tKZfOA4ste4lUhxJtz797e1JvCyUjC2lXEqBUQCDWcEQgAy39tqzw0iCJ4fpbfrzP5
jrskrJoxgINLSTwzJpXk20KUaAdMxKpQ2WQHho2lGO+zJBDBrIbW/XLE4d+kpxB5zpOrRrtiimf0
3amb0LBC4yvEzKer2HofK88Zif/O3uTH3sBHDkl3WIXCA6rtcqldvzQ+28Plhy3prU0zTdVP+mNI
6QSE9b4IEHheXP/MY1WRim8ykiASilj7HseNfTNCjA2/k2Enaqw9yGdpjlCe5eu4TkPF3RrjMDJd
43PZXtbH7s4MauPEcXORfOXMiB/pGMsFWatsUUPkjSLjswVftsTY9412t99UFLI9psvEBmvLjHtZ
l1l4qfFzEjYXqcTpHcCkTc7q2dc2NWcmhg7ox34sS9kh+Cuj+QYFNTTWEe+IYu8nDGAGTi3zSuc4
FrD16x3C5p/WgCGypiTwmbW473BNQo40HliQ3d71EaROYXiASXeTa+//zr0rrB+PtIeREmCTKTyO
S5hdztL/C1kzH8Cra8JECxRusKKXLHy5DT1ZNiT6tJySKcQkLSaLBQwRVyEt+5F9SiWZHnxx7Io+
HXXtywhviUSym2nVAOoKw7YWNIFaqyvTsrK7hvL3255wUetgxYdKJWMYggO1j17L1iOapjbrGmvX
UCbHIE9/YqqP6DPTMlDzfkVUMPPji/l+mEG935LjmroPkfquC4EHrF6pMpUZT8k+eyRJbjCr/i/X
th58/2LI2cUjifY3ZzTK/r5PMYuOFlXwRhEX1WUl2aL7KQe5KDqivBysIWtxPFn9Kh5IPbO4b8VJ
YLViJ5+z5Tu8F9MejKPXCtit6V8vgC+277oG5FSEEqS0owRmmo1gwWQ9Hiq3UbXzUtOkreI3BSmo
biqjUK3eDY6cWKTme4MRYou4UKIKFfqSsjxAnsyoa7ktTHRzyPInBQ/GHq5CyW3SOHBI+Bv0eFnx
Ks+qaKk63g8Jp1dD9GttUDp/8w+Wkh+0PqigDoiXG9637yI0brR1jR3uGbrd99f3ywDm8qB5DHUK
uroWM1iYPhqY3LJ/q037S3O9ld6511AB2g32O96HRRvJ5evv4sl7oYGClFGrlNkir8wEo8ASCcHV
C6DI0hUx5Nji92/LXfuKyCrmwb2fa4YiLl+4MdAv4IqN0BG694JCdbFXeADvX7Yh5Gw0eucq2uxG
SPFibZF3vqGMWBWaIwIz/gHawF1ewc6rCB3v7AU950LQ+OqidqfyPBHfxxZlGaVD2zBUHmP8WqMC
CIe9X1nla/OmZx9zr6IuJMp44qcKXZRVmQnVCCVGLt6/HvBi4rRJa3OuNjD54x7kJo4NpxYx5hJu
UE2HzixK+QGe/NLbgaBzETO40TRR0pOglqYBrv0iRhWTMRF5Yl2pmOVkovCKUK4sMd9ExuoqUu+V
jAu/Awts+F2gVRMctUWmljmiTn/x8YYvbDMZUcMHHzYBNd2ACg1uLqnwtIWR4N+hnX9KzKuQUTMF
RGqoidfefKb7BLIIGpu1SIG9OYHJkDuO/RO/Iqs7CVk5/clCvbZgzTnEQM2UDonnkdNjBVEMe3Rj
uXfct8Q8g3cCme+DSboJxNYoiw2Rxy10sHyTwS+ZyfbMi4DuBaXc4mQyVBEmuwClbHT8bhkhLava
GZmv9MZPu/OXQ6fQiZqQnzLrNz2mx/SdH+RX7Z5JI+DSYEva11IUrqQ5/B7eFRDiSKo560aN3WBB
Nupv7OgZZTd0fW/ky2AbSH8y6xTFeoQNes9RUR70RV4ynXxY2MPADAHN0X8nTPV2f9AzSwkHHvxc
t54SiyhyN+/JNfOhUIGN6jf7zABknuApd9pqNwc4PLqIdqjAvVuoG5SIQYQ5pgr8hV+sKWHFWE4v
37X6iLOwJn+jG/1xHlwnsrpllDL5US7euya+mTaOooGKT2u3SW+jveVST4Cxg3EnlShEdHXYc+/D
CKbbUfSSWg8UUx3kltzJt+wWAy1HNyLiKK2w74ky2qePGPWJji+AoQATSblt1loTSetDZuNXEMON
QlOOV+JCz7DBrCaF/FqNY9HcF7n6l+O76g6PxHWe4taxA8Q+nUymHXN4iM4SAMnV3cDJXE4w4DgZ
/Z/cWLQUw4yT337HO/jiaCgvUEjpqPvsW1I8U4FXSfnMknNmKwotqro/+nnUq8PfYjbg8Y56RP6W
GFF+ttnV+7rkMEJWfoseLX5ilJY07CJ1i2QMnB/oY/RauVh5t8k9oY4p3LTO+MinaEP8cXPykoWX
/YAqZS1xm9ehy4fThIbow3TR7WqMDQafVvdXAtVFWKuAZU/iQX+V0qIsngu+YOz/Au3RfoNP+4/C
hDQpytqavwyYsVvaZ3ZCKpHQY1bwZIStdsDF6jLUKlpuTlVoWrSDoMzjCV96Z4qX+KwoeXrqvN70
rsEJMyd+ONivm01W03aIdvs1vuc2JVtC7pxq1OeGQcie1cVBKfX5nXpjQIZQxvyoP8zDpFzF760/
6jqRFdMIxPTxgCzkqs6ZjF3eX1Mi+AZg/glFLnN/5Np1j2Z6nilDxKEwSaLhN6gwe8+tsArF5dEb
yURZscanPCdQmE1+Cu7hKXAuxeWMk7vwVA5Ab9BtzWak5RigwlTf3PrKKwvgoXB8gM81wyBfr2t2
kEkML9fMyDSyQWRKYD5k3Ncvh1g20RB6GzhEL4NXtiSVKPj8Jq5nMLwfZXbdI808yXbvJrZ8sZkg
YB7U2XDtoDkXEm3Nhr56j6asI/MRI57ZISPmNIAzI2ZxEdw7vRs1GpY+JINwEPtJO/uB/iS3fCur
fxBMbVRU9OSFwzOGaZxumToogHxEthIBH2BpuA9TrfXPjtm7BMtaZFI/BmKtqZydxHrrIUz6d/zp
+ayNRIFKM8gFnQzH3PkqnDlBmbho/730qWuWaVfU9VTLg6BwBsxayZDs2PQ9T0dx9zz34rl3e4kB
yfC8WdsU8JmHrMzcF3GQhUP16Fv652n7VR4vnwQ7QFrLm31nAjgNqGpGJC3P2LK9lFFpnEOh5clB
nwzNp8VdNTyAKu1gNl5g3H0T47/FsXOFf0QxSb88MgpgbeDG8QEZLzqRX4JVurY3JTHjSVcmON5m
wn70cdRr2kfItShVFc6W3mDJsBoQNiH3UZLardQvTzs5SgMtf9QrA8O4f90011VtYZSOKriYdH3F
h49ZQ/q8e8qgU9VjQtcy8vnM5KHSCC/w6TYiKX4175+lCYV3x3JYjnPzkC3HtE1XkJdclXCfwPZH
SvTHV+Jj66Kc1HbltsyeplProUlQUXZF3FU2g5D7vk8HYsX/A/tzUdGLgbAIvZznXYdPyhnLWwHG
6oDuUekFeziR9JSnfAPE1AIU0FMi7kAIKOnCr6TcxyIr1cElP1EpaFW87sxggsFP4goKITVgmcfO
tpjkvISxTmY/f7E3GByl8drRYs7qliafZaqCGapR/0nyuSTWjalGOdLkrsnL5NNgNbh/bthThUmA
7W5UnY1CO4O03t6uoeS++l1lVTeS7XNyF6uMtu2lFNBhz7vK/x9ZkMh4Bat3zjTaNxpAhxdMfc5/
UYaQ74FRPJGZNkR+UwJ8fr7xcnxwrUa+mXu7//Oj0vinNiFC4v+owr3mYDnrEb0Qtu1FRmPtIRUP
cCwCvbiSjMn40Gtxpe5cSFboTwQJuQ3PeJzyuSxrjoTUpJ5X6+JTf7WdfWbhSE2qMNX2SM1CnJAA
WfoyG0dfgbvAbRlSW+c9A8sxxdJiFmB+bZqQdjy+OxPPocxK1hC3SS+1wdYShN6XioM9RhOK0/KX
w7QfKRVdlu0pGnSJKn6zHSKsb3EkaS5DQWuj9L5HuT48Igsva545pUfvJ6msk72doALyVdYRgiKi
QewIPIpssy8gpk4Ntj2QZ6/d+UDg0ago+SuUJ/PY6emqv4CFAzOB5pEZkHXNCmghq8RoMvi3okG/
uu6oZWFZGXCLaepczMOyRXFpgaPDHfCHmfvCTtwyDafZ7y1fvVx0twS4+OuSqZ6pB1cYduS/hkpD
6Xeoa0kXAK1Pg3uQCMtmxouUs19YUgblvxHAduLMfaEPkvsO9iL1PRepaSih8sYK7ozrySUBRscg
ad3XzzafhuSckr+X9nGQ0hOXQ9aaAOVqB995W+mX5hm1q47rkY3L4sS0oHB1vxecl2SjYVdAPJPB
2bPrEWxOTpOHrQhkdyswxA2avtjIFmuYWfYw8nnEq7d36QpsZFjcuHXMqVYUJNzO73OXePns9mJ8
pX0D8uYWArNKmLnij7Z8M3ffwnSnXcerSochD3BB9L7eRqTQFyNabShvV18ry7lX4buz+GKFgFfr
95yndIrTILpF6X8uPiPuLMX2kLtj84c3XOJ4ruZkYhK970LoTeEtYE0bzUmf1zKa9UiigAk0n1lE
e4ocrsVMaSQOYiqlcmm8Mu/ADow5yFGkqHKCaC1Y70AQrHDmwyblm8uP5BJ7j3baM+PpmBCYfedD
rWNBbeamlF6PAazz5fleoDUH0se0U1CLFGSVttwMm27uSC7g6e8AbjXK9B5p5pHNmAAjdO43gRZi
bibAzs/PYvwtDJtB7lGTvziFfkdOxX14+zp1gxG8iB3KzVf77Oltu1u5HJwAVal3CdplI6BHGlkT
uM7Kps3JN+445cnc+/gdbYLtcGei8XldY4LnkWSmeaWC7oZW4W+WHSkjkV7LDCJBu8XoDedgX+qK
4WK6lZ3rwveKSPHfe3BcvlaWznEkahs10IG9Hu8NQnQswye2NKDr0RSFMwJprefVrt4AZK4v8XiG
y2at0s3iW8nNk0bl6DddmFrh5CxvIGorG15ZRXZnZgIFHh6P770vC3k+n+ZMe1E4KcN7HGORL2s1
yEcADkZVkyJ5/cnJJ9ZPc/INaqb0eKrExEZbCZ0EsCoAxrg+4idz7LfwEMSXIDNWoyJxt9MKeleU
WhYVC0zZziAM7Jrqar6pcDK+JUrriwOjCOLYZH284EVkYIZPBJ3TXEDVBLOS2WlbvqjGhQe7a8kk
BFu9y1zGQbRfy8S357APS1LMjP9sJwQGg9kZtipZfnFjmIqC9AB7NKlaFFgEGYVrk+DvDeMRvakG
juSHbFryx8m9QUtmufj6ALLskC5NxsOwhBlosLdjOudCYd/83WbS5LiJuXEzAy20BJOtjy9ELDcs
wDGKDRoIQ6yjXzKZu8m1IP4wHVjrouBzXXVhL7/V3XTWarXXAdVBC5esxPfx9o9kl1e9LUjbPhih
WbMn/o+QE4+aUj6YRaiQlMaN/+tGPhokBoHU2hmLkzREQ6ByHG5ymR/IPsr18I68LePvNkbG2FUY
4dyDYd0hc8NuLGdfwRCrW6/z0zeLtGqp91jYyy+LOU/rNjMsni5hXH72NwVaev9aqrefHUeciM+E
TDHUpBPAoAE3Y6GELIkA+IPr5Vcx38cM4CtarY1rhOW7XmahkhYz5KTOHdqcLngmExfupEcGHlH9
d27R75u3MSSDSGv+KTUMlaVwFobZcY9+lGhBzenKvAJ0yTQVC6rf2OI2uXujsWipFLYFSRNBglsW
5WlBQP9iWlrItuueuONafB52mAP7Svwvsv20C2MscBa0aSxaHU9BCppZBoVMu0UMwWxeqI86AyB8
wHQe26lwi52JP5eS0AqgQCaVkwpoAFjLCZubWC6ZuPH0kIsiGEtPXWD/ULSsTEw5k1BxbWqamSpX
dLs2q7pbY+r1Qdka3kbrtZHb92HIjcn8f430XTdWk4PZL1MkySiG/vUvgAyBM0MBd1VCJOAmk3IA
Lt1bkgVX1wrGT+9Bk84BL41BfY0znJKp8/LdwdY+Z8v0qmyjJomEeBr3rxrWdmfRY38v3eubj4uw
Q4/SicIc5tX1qq+2MDzUAC3T6+jZh5KTSHNev2b5Kfud2tsOiZsEL40WR2sfyQO7GoqHqDIeUQgF
OHOlfUmImLUUySF/k/Ab2MEMYjJOmPQNksL/I0DAcyWiWiEnGGxoKRZIcKbcMsOND8ulq7gQP5ZX
BauA05zOlZDP+qqQn9zQDcU4JWxtth6nhNmxqVF3/bitvbvSkLkuilqUI2FhEKB/EmOaY6clGcdQ
nV9yG6wifBYR2oA2evk7Er5d8NutudEc+T1XxeRg3zLbG+7xC6JI6gw8lEgkCcgOpc/1XsMnRPp8
UHxUrgZXgUov3XnmNYtDnYUivX01PjiRkUotEyEHmZlG87b9vcI8sm25SN8aoYhSI3ueE/qQf5U6
ENFPn8JWGecGJoJOi2LHdXwBHmCbaKOOHHc+GM2ZorldtpNo3YZ++NhBIeuOaJ/k9HXty3DIsWqG
k2cvBLoQsL6v+dmrVv79fKBDlnVwcWZTY6Oet66TeOXZKI8Eq+EAmFcVSUtFPkfDOfOl9ZJtAl5r
3svsWgQKN47+KpBXCZq0uJEcDU7wE8VvYiqVzdTglsbed/2OEroH305cDdpERMBUsgTsgKY/6rsP
Co8tYLpEAvKGg9+UG6h2pP8YuZfA6nUhdghRI1GcsszNNtXQvKKCNlcLN1x8kMfaIY3ZY+86FRWn
lFkcW/SztAzmECTIHvcncLQh+aj566oPoTkury5mNnmQdBZZShraztM3ndwlSWu9EZjRRZMmnyBU
KrTvF6BU6c2nM5CFKi0psH1gIvyoxREsyPWmG7Y4YiC/KUs4iA/HsLce1A9y8k2i3Y7awrIpG/OU
grUyR1hzBZiLkpzXvs+Ow0MAmF+j0ljJNvvd8YqeRwvyP+t5buLEwfvEiHy2aB1NZ7RI4jjgUOai
4e4Vn3nIvt7hvBWDX0bBfFBlTPcb7kHuAFS1d4oUmKejgDR5wiz6dFlnPMrRRFNssRtdITc4ffza
O6IbRSNzgm5MwWMwrjw73qeFKCyl5hKvZ+BB/V9gtHn8pTHxy6p1aHT1e84grIhx7v4bUzsy46Ta
dMlpqhvrcqyJlv+O0IkVyDmidM1dK3KHJbXUFXZOTY6aHwE5sbh0DlOXw+XuN/aNVMmJPGOFZhNL
d8PjAOVel442MfkdwTqwhWmY3Vj6J+RL7cmIL1VB1qLFewfIOTo1K7gNsPfyMNeds52aQq5OvDfq
OowRO1G2Otnf0PaMNFdnrq64bSgz0iGcqmEzFzscUA2EPnOrvlmDUD8nuh2TEn0fCXCgypIl+Ml3
NYYIzLoN7awpft7mC77oD1Fu5ROo9eyiM4kkqIcCQoYg/UPPK3n8PTuIE2FclxXjqlh5AdNfDCtf
ce7azQddI6YuXqJG4CiSxk3U3F1eH5eCaXH4HYT52/3m7NJ9+qw7JjJjzNRQ7RINA5kG33qx2dKy
8R8fKdkwNXzFimcu+P6SveDUxJ5Jvj9glZqeNu58AFAONVZ/uZBegd2rK9N+OwZclIJm0wzeVGTM
xyCXTH+LFJh8kfpXum8EXp4eeAqKQKHt0rZnrbZH30k4/qiKRiJ5pn4qmOrXdrja2jj3s7Pp157L
9+YGkmS5NLjfg4OieZEH8rj0fJmZsczoPehyxJ0JhUxeV2jixdSRJLPjKigFlmL3zT37YUPvqcvS
0LWmpDAUU6rAKMXQxwE41Sj6gKdBefLCP0oqq/9KDuU2CXWsVmCKbIF/rQnvuGcov/nPY/w2anea
xC56PcS0a4Igz+FLfZH9aHssuDSFnGV8yNqaM1n0J6DvthJjnF5Mtpsj00Q0w41JBy/NLzggytdK
JNbruzr0K8zLpmhPHShoZ+dwBThfpjH+pNJlk5La88UdR4WWJv1v1SF0LEXtutCiFcpfIVzYlw78
7MKmclSBlhQYzXuiVvbtAWJKFcaisFoXTb5bjDaCBCYRnkqfUlbASz8Bif7UDcn1pwOXGIgFyQbz
S0OkuQUX5KDEw2qJ3wqdc4r4zk8aQod3EDXYHl925sNjxG19EFMvwCdZvqfniXwk2+BnNdz8gMz0
VMxr4MCB7X1MD47JEIfFrY0eAJymfsNdcEZ0+PKT59b/FAgq5k3nntj8MW665ZLuuLmv4MgQH7ae
U9gql+vEEyWohy5pFJT1we5gZXV3k/+o1O+XX3WR1WLkFjwfWko7Ku/8FDEUipudTp4ooKRzYtU0
9eF90fiDMpjaZEYqiPjDgjtSjUw4LmGj7A+Iq/iDdKouKBR7wIXvnn8lvL1OobyT2bCnxBpRiWsA
67eeoH49EmjkSgWsYZNhMsGVPOGW1fYCdqfLOZh+kRXIw30LQVsrFN7h2GN1ACROe9w6sN3om7Wm
4uxP9CbAObhJltqtxlDVgJewhOQwCcnDGBYARTLZxVJPyYSt7jtRzCcapO8K/AVatIGq5IOL44gB
lAzZFKzO4EM2VYEOe671JeTwVGbDyoDJ5usN60w9UmYT7XI7Pu9FXfESGhFj76akL6aa5Z6bQmpj
SOEb/S33pwPpkpvyU792qQaWeuOwldLp2H00HlLO7EXYdsHIyj6jfSRVLgxCWApT0+6I9M0CCSgi
hXML3Hv7pYQ4QJV8OXwbdBsl7REYCSmg8j4T8pbLIdowfLpNqTYEGrQ2Vv9nKEIp2h/TnkLTnuht
WU5ZJK8dVRMtYor3xyZcPtqxBLg7AdAgIOoG/8oyKGV0K5buAOoK23KnkBBDFoN6gXMydZbGefWA
NFl3Ez5n5O1c8sGQYd6yD1wMRJt2+0LN2oLpPzUSxf2XVwMOVaa9MxVxsL+eKOggCTyz9Tg6TI42
adNbXbta0IYlezi1FBLUUYiry2W3fRkeSzoHtutiI7Jw06ZAMqpWCqgBzG68U+vYIKe1cdWQLZg+
I/IAvVedbPmeODfNqvKd9YdgAKSkK+LKt2ifgPYVxlzL4aI5JEncGauk25yfYCD/s/IIzVK4v6Ks
yW0hfdFqnD9Ux0AVk+goo/j22UlwvDghHbkPtDyp2dYq47LRvmze+IjgBt8iKKU1cCr5W/iJh9b8
tR3lWoA06IMAaSnCZorvZJcwTit5EBzuvT2tyP76iBj+stjAQz+rK0SiWk23hKRRUS+Nhxc1+Q5E
8uF7NEjdZ9MYGdodm2dlBurWdbF9nYZn4UOu5/hMI3V9OUiaqsl+f8aTnFXPeUGG/ydL+vE1ImhM
xvEZ9rhqMJakI91T9ytUGjUE3W6J5VF4hrWHUvjDqTD5CAu4SCKYdv2Lvi4mF+BuS5+Es+Q7LrAh
DD3CeF5HXJnqr7N2l0SBUQfFVBovEIS4vPi7WQmC0UQuV76kC7FRAynoakuNUZ4YkviCSAZwn26p
ZZpIHSXoGpBkRl0AbNvMQ77lEv8bQL1XjcnQzVzlCWU7/ZwEpW8IRTSyTnQ4grehC6A8qW8EtiSl
JNgv7FwJfynjeOrY4YFn8ptnA/7svamg36dhemidNYZVdw5KJg0mLlRqORBUEk+BN5C8Uz3pNo0x
nlDi0GFSlLdW/mhMdLjfFBqqs96mCjNKWa3DuA9AVeJdZgLz5Pj1+hYZT1ahGNAmFxcivX0Dkbqk
U7rsLtZ/2xGUD+NRaUAQjlz049uG9UfzG67zsUYRxAfTJp4V8H+i2SPLV20dG0nV/vRm5WJ+NB2N
SJMi9wfRls+T6kHUss4sIHBzRIHXmJa17TWTJIu1t6F+2J0siLQG1Nevp28pTHpB8z7UAU34Lt+n
h+5eM8jbZ83vaKPe4nygCWb/RXmO5XgTEGWTvHd25Mw99D3rXqdl6/j7FaTEQmA7nvl7lp7a0dD+
4NTWRINQLmofTyrfyMxjSHoQcGXlLC2mPFTn3aHjOr+J8aCwDkh+Z9IgzyUCy4b0Dvamgz95VWxF
qake2jc1MxmPLd1uHhKKQ/PgBuz6lGfMI6mmBEeAMS9QLvnW8jUyq/gqAJ05+t5b62fcIqDtkCQV
2MB/84+gvUqkgrLl3sZvEfJ0hxeIXXvkULPe5HAWBTQ9VQKI9QCmj764WD6yN1CiwsHwR5GxwZRd
EnHPjnz2SmeBKweKZ7YzkYEdUMKfQEAbl4/Q3BUm7YInsg9sSJYO8d0kmIe5ao70r35fdDF1bShN
5nYMJGbOOp839BTjcwFrDyMef6pqxdmRcSP3OJG+s+ErRxUNgLVANutFeRC81g8isJClHFj5cgR5
ZoZIHGOdMtbz0A+AkZBlZN6jQclskYj9//qwaMK6sEcVFmUpWtZT7zvunG2k+qth0h5CxCrvrUBf
iJ7vYW/Zw6q9Ijsd1uPRHZOBYDnW6GwueZkzPlT6Nl0yrbRj06+cPeGr/LqN16Y95NIqdJDRFcUr
3otObyUtdA5erwQFWyOj+KrXjZdDGGLu2/7FQrdtBfKaK0nWBRICwtlon4he4rgIpPIspoy6XOiX
fYTWeNAShQphBZGHjqHVNyMmnl/FCYaGtcgN1wsoKGL4pL+Gq4vjI6PF3X3NtoF4dxQXbCGVzUKt
n5ftbXFNpb+0u+cYZLKadhPA4tASOBneGarJsOZN9URzLFCtRKqrPrf309Ytiv5+O4InytZJ0kM8
n6RubdaGi0OkAu9FXzhOiAdPBf6U/pT3BaxWccQ/Au6g4XUoAm1jsn7nXbMkkj5Zr9/wa53bRh3t
kId3kO9vU2XRo94ZaoNKuQd1756FEWVQTtrqKfGuR4rqIzPBhdQSLwGmZduEJhwC1Hz8+hxh4+5O
4grErHxgEbQEP07EoAgkNqP+EBVHrKF8lTAtwU9ZLcJKewciPJKUfQhxKujmy1w4GireQ+/mBRgi
SXIjXMXWt/pWjrjnIopuP4crheJ839+OaTKtIEonLBkYt/9i3LPzs7S+gaK+YieoXCrg+tkaJZMi
iignq8G1BRi525OmcmNvG6to+dX5OvD9rVMJJotfz+WBaWBIS2Zi5YoFQr8RKXpbHU/JFYIaysvi
l9DjchCA1YKcML/O8RLoHX8WAhsAmyclE4JvyDTGoZp6H4H6RYCLMxDVzQD4Y2HgTup9xBLv7kAv
2syppE0bK+Lc07Ga6xFwkl7Pjkt8jzSLWeYahnEWm6+AJGxvbqcBNk7ZDuMUp8MMAS7Sh99wa+ND
QS7rAHoZNrO7AtORxQnMBf4GdAgg6kUs35gO5PjoV6UwsQlcACG1tfd+iitfWrCh9aNtW12KxHOE
xzZ50TMknI4D8sFvWABHiMVuZZ7mzPyGOAYrJ44367YGmRFFXIzYLdzH2dynn6H6U3mYFF42NZt9
hET0s6qcEi/9DSeF/oZ9xNffmEICJlgIT5d0sqmiXc4zGVfKbiPVI7d0ujjOkRfHgLihTEfm5Uls
nTQGVAvCUqqAG+WuWo9l2ZnXPjThBmzrpFKHk5xKbQwjEYq2a9iprbMugnSYVAqDbx8OAApyNN71
24cr2pALsvPwd6IXWbVjOp5mvcCH6L1poidciQAgJospHCKBECVWumYxBUqt09OiPM+kSFZQbzLL
LSQQeI9lqUOXIX2tL6LmyhtmJcqPFEIWICIss9CCohCE3EERpZ5n4KwGle8W07BcfVomYLcLjC82
tJFPzagroN5OSg3yPQVZgSdsPkg0TaChB1CXGVvRWWnmgFMxRrJaGajC3X8SuYcLxT/YWLoGsHlu
cSRUWzeC01xyQU15t8AAp9RQBPN1lNDTDfUXoGEZ3FIJR9Q12hPbmIjkMuirVhnGlPBoKJgSThcv
55ftp1vukNEnNAE4yuhHY4K5kNHxrjAJZrGLKLxeY3mhzXZsayAK6bEdQ3Mufi/zAsY6ByeD6F66
nC0Onum6U1YBPrCaLez4bXRwqS8kUKE+sRIDhVOFrGoVgtaciJ64bmepw9KvIi5mtZE583RCIEBl
yg1ar6LkX+KSSI8N102CEykVQv7EeDcT6iy8hXgfftvAL67gtuIx8NJX5eFyI913fb4Jqp596QWC
q6uLFTt6WUhRMLOVMY1/l5ydmgj/vHLJB/3qOPLQtxa0eHFEbVC3HQ4yR0zQlitn4MBwTxXt6IaY
L43lqEcbCEAWVvgJL08QOlC0wT7ah3QpcRhvKFa4qbDFML7LU5Lqt9bOoH6M7WxrZppJsG7ig473
hyRVR3uu9Q25OrjlNTM8ySg/gkTDldeZbwzu+AfYR5G9ftuM0x+5nR1hjoiATGI4SATo04YhhzUU
1QE4G32FXYFSWiwPYCD3912/vmmQE+jHPCGB80uICyRwJoAVIV85N0v8A6FsyMtWpprNFBAb/wU8
tVyhRIThI8+MWv8INAVhW+jS3+WVhfBvSWNZuTsHq0B0+6LtpY1ukyPs4dPPfHcmANZ9Db73ooE3
2kZN7pZ7eGp2xXbIZmC+sFBEmrSFWwPoGlvlub6rlR3Fub2GU3lQw6kfaEVSmkDt7O/BfAp5deG8
fqJb1kR+CgJCvsLVovuHKuPzANUKpc5zvYri2K9ytkt0JR2+8yGmA+neWLnH3lSTq7Y6dO9RZp0e
7TeU85e7okM+yG+7FF79bVeVYOgbfSxtpKK/WcKZiedY7hanCdpOPYkTkKDauU2qpJ84P/mtoFEx
oZk465YrP7NshYhIh/qgHq/nAVAoiQ6wIwzdZzjBysp6PHXkvmq8s7SROIbshddtWSgkTFa9VzEf
4V9Je87WyfDTcF84f3TY3G/FazIOAPgqwkehPQ6UlIyxETwbN1rFcWEbgqZmq4gwSDApzKUiAV9F
0qa9la336ShjKuDFClNBMenhG/iM26lcS+++YpcrFNcWiBonEAq6tfnOJaMxMO6UDcakN3MtLP2b
ULWY/ZvcAbqfgIvrs0Ifa00g7L+sjbySubCKindiOPoEGqTjwttyHj2TMJHnCy9fBv1LSvdXZ6eG
qm/rJNTfHF9oGgjPEbAEz0PSM4XrbhSurfroBPEgBsb2OqjP9ufTygHgigqRw61acadYDasUyIoR
tW+TDCBR+UvfIXGIRNaq6Um3HpgtwEULa+e7fBfasV03HI26sbzvBUEPkYngmIrRfNyN8wtlBeyY
rF0aIHPZTiTtnn1AqspYbZ0dJAPVoDa77maAub76KeW7i/OWAAPEWJyc1r45HWIR03FlthA4xAop
P6wogUKAzrO332FYuDXlMr+pUnjwjBvwG0mXX5Otn46z2jTDIdJlh5owO5uMavKQKRDQwf7MO7d6
p1p/QMKLg83+VR7SatFl40fi4RJPszZvEC8JwlQINQuh/ohfdh/56hecxnRSHrD/FleFGacqXzJN
ejhl9KQcluEBzGLvl0FDi+SV80rxn9kKOIp+Ep972FCqDhKwTlylJMpWiMMogB3hRsawPbXDHSyp
r3vOYKQoZ/a9oCLWXXofUfrDWPUaxgO0PkSeeSlRgxpHRZxbVui/5SN9gtpetJYjxKFOEewi/YfQ
wM3NmyFcVddYDgsoSdsd7yljz031e13Rqr6bqDYX2jM/M5vLM6bdG3SzRR7Zw7IidqB+4YKFIjfc
F5yaDmoxRS3N19qEy9i4Fhs8mmGISs1u7FmqvDlbHyTeuPtyHwZld5+Fw/bm95DUiDe6EMR6eG+V
hgE3eUlZcTFbYxVlpffazejbfD1ii3FTGi8fF6KFLmGqoqKhxg9/Lpqscd7ckOH206Y8oI37semi
eNsFJofNlNQSTHmrADvlCrc/YFkt0KzxgWCkONciKNaYOPFyBDYCQhek5STN/gNgm5bAJW4xMmyJ
SKArn9QR/EnorrtVPKnSR8VRdUIBqCB+f7/KoZXjjYESBTps+Ng0WiCeW/p3kSoj2ebRHfys+f2g
hax0JyKFPKbuJrwzmImI4BaERxpTyDIt4CQcuDW0EU1jsX7c5HUtkcgMJBJGOlqs4iIyHjcOBDx1
8IBIqLrXETZ6OZhg1easZrzPoZOqEHrPasQ0yFgyvKAiNiHkHIfVgmhGJW9bJ7ot1QkE9vOq7fUm
7pSFHv2mDy4/KZ0XBK7FkNGSiAk1jd9zwyvgKLcwFa6BRBAAKRnePgKQA9GJd0CN+yFMCv9waPX3
TqxAPAfucz6R0+IAcn4z+Jwuan2Q3e62KqUjZL7kXFI0SntT+MRXFsB1sv28cESKTaBJuLfA4VJo
jUm4nxHlmzNs79UxouL72Z0rPHJw7vL6ls6i4oivLmjte1V2bgG87/c8PXfM1lXaZJB9S2XNY+ZU
keu5+2Q20/qkZVsmM1orADhd5AalcOFZlxF8lCwND2vnfVZZWKGyzFT9Qd2skGmAIVSH3aWS2uq1
Y8Dfas+43zNXkhJs4K6XG8bAq4y6iPOWm3KPNCxX5SLz2VhlPJK3qkDkTloStzoXnr+cLlOSQ4Hm
adtRQiBj0PGwzO4wCOfT/pnzJSTzrn48BWYoxibihiTFnhCNbTc7TH0fHMkeZpK+VrGytM+68O1e
re/QbdhexZG4N0zWKNSUimtnhOXFFnVkYrurzXwAiZPr3bWBQgxbbBEcXlNZhhcG18EzRNP7gAsT
NaXd/Tkfonmrr5BEV5X3xRga3wqvoQVaPZzhCJukpbG42cm52AIsKrhzzFbMeRY6OUCoMFr25i/4
Gjo0XDgGAr38zzbPjKTt/vkT7Cj1KKZWDCTtgj5sFu9Q2WalhQPKuh21rhDCN+V5SwNXuny+ZMFN
Bp55iYofNCl+2/I4P5SxkYbqpZCOgIpqDemq4ySDcR32IKmIyG1aRC02ZB3/kEu7Gt9bNEkNbp+V
V2nFsx/PjlTT0BKfpGpmsQt+xYyfJ7L/5ieQEsqrWyjJIhC3C0wdDSUJ6ZjLZK7+Pm0PFboqMYmx
kMCeGyBtWaFcfVnW1XgmzxOaVVa+9NzszokIfD07VTLH3yAj08SFY4UXY1YaoU2fKSZAUNFUToob
eI6sF5VvejgEUjqDoQVBntZ+fBAJcvdj/a4YZ3v43XvgjRntL0W+LrlePKvk7p95GVGT8TZrQ1+I
eom0N8uKGI6052Q+fOSHpeXWnJjNxh2pF9fBxQkPkNYD32S9q1P1OOzxC4+2QzboDerGQDoBOBRA
V7ZSxdGg0WdvYAHewm+jnautHRW+Q7fELY3bMtuwcrMz9jxNFaDiHVD+3Yq902dIL3UNnupuHt4f
+sGUtB/5fx2phVmI46i+lR3MnSzsZJ9/QsGs7JLJ5Xwk5YGNacscgMVq2bbLdVUbuPybOpfF3xiV
qHZabSSRXvxDlU6u5gpjzDZ2AqJHBD74deoZZ4EhOTcvXbcFCYQIBZg9bBxajl2Gqmo6vnQLZpdO
fNeEUvj7qA2agwRag6aZFtcvYvZgvffeByo10jMfYuklj0crNemjCAhwn2XCJbmhyKzHCkm4STFM
BCu2qArZPLcMuVY92MshiJh+FAjjAS1QsVW7UceoalD41rbG7kpw8NzQk0hpFkH196ppOjNhhBqi
Zqo2qerN0sYfAtPUtlst/usxBM06mdpuADA68LHCnVp+SvnlIQz0ne+sh5Gr12njr7ZrUEKrP48L
BNHvUfnwYuycs/lM5vX8ns1sU9zPEUFtYpNFzuAWeaLnDO620kLYnVZWlI9HeBDDiWVad8lPSclr
a/uioRVLiAcrzSIYQ/oKWM9CQKJyf5a4r5D8YR670zdD2/J+jqjYyoJGRwfWCVoLTs+BSBd2GrN5
nY0/DBdJE2FnrtcDtq787cQCcIvJPso0vgrr7MJqLcsgnGY7wzz1a6csubIc2VY8buTC7xuh6vz5
qyigHViqRcjHVz6tCjAh246iF5C/zC3PjZN9bjSwIeE9uT6uQwgKcgKiz5Swz8uY3TWrmUpNrDOu
C47Fc08bh8F+ipG/lFRsdXwPZikdS6LxZCp4yHp8aO2zmqRwCAlPG9QA+gW7LukluLJL+XP8FUbr
IbZXG9+/Ritki8P8luI7fXAcap3adl1cVYjlveczETt/z33kQhePNA3lCzs6N73V2LA0g1pVZwYT
g9fvQHC6bOy07dAdiWy5sul+sOmflziSjheJLNOI6vEVWty134jxI042ejCr0rrLiyi9gHK251sq
uff4lcWh1PgPRdUr1F5xcNvyd2LD6srOA8elJ57/K8a1WrAwPUpY4cz/wThmEKLdPBYkfyix+peG
tsa9LRRfr+lPEZCtZh8qiDEhIcUXvHvQuotxpsHcD1u78MJbzSTZBv9rhNK/dSMQZx3CZUbOokPQ
3xyG9foQjcsBim6aajdtuBp7hEJSMqS6+vadIBYxeTNN8X+pj4/MHEerMoumBUd9San/tk+Yti7w
K0unN4Nao/baIWtgmXgZSghZkOTrXpASoueHpRJvR+dEkwK4eij4Pq56e3U37V8e5IPaVmNofY5p
nEYbu0FxoCvHvqOgQ5sNTzjxKCRzTyv80ma/zqjS2JchEwZx+nH56FlJT6WbDEiSQ5SNtNYbM0Cv
3Ljd43ePg8j3uvDpg2neUYepg2sJBY+fEifgv0G0W8w3/wYDQ+sJm6AIilf+E8JANdNpABqvzuPa
y3ZCif+SO/aGk1UGUn5y6E4R72wmFLdEpALrqeRiFxV/Xwm3p4f8R4JwQ52VJfjYD2SnG6rZzFPb
njxQEnaoPpG55fhtvXgTUBHpfg6WRQWdvNEXaG8mPPnXS8XWZoXOn4dHFw3Q9SuVmzVoVm3YVkvN
lfOYGlWjgOsjVkHHVYVALJDMC+EhKC0h0xP7c412ojS1YmhzP/XM1u2Uivms69XsgnJxom8K0/BV
zwGUyNkPZZ5f9MQuJYl++yztoym/diRa1mHVlmMtCbv1+KSWnwbUgPRAgEseL6H4KojPXzrP3zJn
DBkb6snegNx3ZPyMtYpB4avxYwqpiTrfwkdlUIBDVAIo2a0HH82TvHGMrt1uG+oV2dAATeuOb4su
oAFzKmtAvFbp6XotoQ/35UtTtEp1GRw1VY3wDvojCZSHXwKZ5A0az9MXunhDmFpj2zv/QJ3d+hix
8t3vxaHmoIBIuW3oxz3bMHszFQOk56OoaRoJYBoB5ylkOSgvISA5y3T/rsHtOqKNyxKj3ZW/ZlHo
zCufD6xlmAnJGbw5fTxBFIegIJrLqgL1U8BqH+69kwzRnMM9txnMRYqsEe49gDBbc3bOkNJAeybS
+47PEZfAWJfvMsYbKLWX1CsHOsaHgyG9/ngiPjpS/+hljCpTyW42isAbT7LGd84K9vKoDeP/X6dQ
LGPKwvt037nSQp1RlaNj7yJDa7ZPUtCYVVD6dG+/PnjQdqoLyEHEFikTCY1JkB3xFIe8M8tjeRgV
aMcSpfgOFh/6StGwpG1w35rwd/shBuMO8Cvvj4bYMrJHtU+JV60VAz8s7mZ4HHyuVweVsFKxW6sz
TgWIKrjc9JWHKMbh4fGdqA8qjuOZBzoysy/CBNBrxaQsCBRt+rDpjmcNs9PrmKsPhYqChQtMTkuR
zGPyZdbIPpyn8ZP40S1KcL7VSL3Qjant3gKZj6zSlMmZ7DOgo/5vbXmFN4YkY6iCxFZlCas+8pZC
Y351m6ra87nJR8MahYRcBAav99aIrfYyTYsjqpI2ngZxJdbs0CTHpy02Rx7V7bJGi3HTsCmWjHxs
IdvvN18aBjWloTHPNfQWt1nH2KxI9Rq/Nm41+P2GPhheOkAI5jgWQDZhwdtGgKfWfJUtgH24bw9z
4pCC/SrOy1hrKHOMnf0KYuhPx2vT+YRrEMkuxInKiNOnhTKdwhmhZKCFdfgH/54V9NyfHP7yuyXL
j+kEkF9uuCnH5p51kRirF2GKuvgT5+M/rTN8SmxkiJZJA0AiHxieUE6Ph/c5vaFfDgTFvGIsKNAf
aDjaXqYYqCYoYwlB77Ij4ThEdQKrH/yv3fzPWE3LSrPVbrzMY+JaiPmmTfZOKwMcAzkErGDVrb0V
T2xwbskXSwW4eRZpj8VNEASm/Ns0lGHFnrZi9cW4qhO6DVNKlhO8DNyKTH7b/wdqVSF7Y527o1av
NQLiycOZxCVHdTddRhuyAwA6UY9HhTf4nlG+r1UiVhelLl+0PzXsv2HRsMs5jmP/2ffDGGAA/ahZ
JWd3ib27axrhqR1Z0ExSuA0xm18hAP5Hhufb4YExfeOPhJES2d0bEzBTnKcN3q5jBRdm2EjASTWG
Y/jyUzcb9ecYif+yITF6lApzxikNQAmFOsPEVxXKBdTJcA+Al5nw0ade6CMlJKaLoovIsrkniP/P
7NmFO124eb5aQhmWNF6jFSnlFO6Qq6dKngPon6IokuqQVJ1okQbBNHFhYHfTBHrUtcfrwjQO5B+r
4EWPYsTZf+DZl/LgGTSxqOxyVBbZ0Yqr4DcGktoZ0hE0KlYMC0z+EZ8/91Wrzh1U9Fixg1HUb6TJ
7uWCZt2NamLXr4BqTOjsUB+JprOhloo6uPqy/rXKx86uBqfyaSQZL76YPy9eMQB1L26fmxQQIZ4c
rpptHm/7AKO1+G/OiubvhTQW2C57fgkZ9VS76e/N3unM1ZF37Owxrce2tzfeAnAo+ybebgCq0iPN
8o5SVSItjnHo/8kvtxrcYOWqtsDlnNbOM386eqD+uv1qJXHBjKT1AdmxqPJBLFR0MBOsAPRiYdtA
KMPOyXO/X3x9iShiQxmBzkkEzPUijJUdqrfITsjKQUihbeXOEK1b9TMesBMELwOIppbuCk+YTCpi
prSijqVuAU4BQ9nDf+A7ZtWq9JOJ6/xTtMvv9h7ukSFss2noAKgJbGutP+kbtR/PrMnTV8BnoWuF
Y/78iYGrtxq8x38m/Pk4+XgsiOOeT/LIunJiIyY/SRDT1GcmWMgqh4Ox4hDiJvQaV6Rn4LvnjTqg
7NbVN9mtZhuqZObMVUt2F/qo0H4cM3GUJLEcBJgXMoXzm2vbci4sBTPJa8QTs/d5r9bUpfmR+MG/
e0/tT0UQTZ6q8pBAn+B87YRhcj2bDCvu2mv5khpdWd4t91TDhQe5m7TQdFPbF4+6ZusA+tPsGj5K
FM1H8KAqODnud/Ay9j6AcY4TJ8KGWr+I9aKjx4adpPQ+7Uq44kTVUsx/+QKl3EQjvn2CMTUe1aqe
BXHGlDVur1vkl1J2pV0wA82aa8htdyuAxLoa7DjbosAkYNwRZWPjzy2WTy0hHX2+TjwGLmu2otGN
9wxe89SvTvQNa32xAQU3/HQn65IN5Zmex7sFQqwyFNG2a+0YpTL89pI5sg+CS/tlXzx6Iuy2VADO
r2HNEBFdaFN5JTRZJQnsx2zSFqreJ7Z76oSJt47VZ7KkN7b2/hQijcTZoJph9Ts/EOHytZLxol4r
297q7P8brolUnkcT/mljs38wNtgphEP+QD0YZi8wNWjpfEb/o/d9PNGx34oNIK7oesp9BUvjWawW
/HFK9VBGoE2QwlTOqktNMhBDYQuMK88vr00vObWiyByWSRv9mLUTE/jbOLUvFEqvKCICzcV9Nhcu
xyVxlu96HdZKHgRcJArVppVAcSHXx9BZ0HfGrLCYHDG3IyhsKQH7dSQYI+jF+/jLtoucUyD3FCel
0w+//DdHQg6qTV9OdTgkH+J6zc5CQbJWZrZnVaFJcgdDypkBfeRwONVcO4eNg2LegLakQ7cX7Y+x
M2Lq+yhS8OCMDoCLUffC4efj0wSKF14hK8HxtlgFbVU2M7lPILc72svUC/FuTOZUSE/AHNxmJf2C
bwo0xOovPZi/z3QxJJ5bpTMYIvZL2Ra0O6cOB21LX+mAqGFD1FG9Cs7C8jWqdhdqemsGmxb6PhWM
iq5MtqZmUJDnEJ4bg0Mp7ur360fRtUTAAiWx+C26jqKDYhTZgKY8CCS+Wa67AYhSKnw3au63X0xt
tInKytpv87wnmRoGr2wuvPCfJeaCOHKOWBdbG31Hzdjt906tQUW/i1zaMQqdoXSNIYENggNxbEyK
QfmOXKfJOUwgn+tLhdO5Ejd1KKhDSfd0MCYjniZnofNQVenV/xVpxAWFl58TmIVJ4VaFMx5NCm9V
e7q5yfGhZiUvmji3idHYiboeuDnFORVMbnwvnnZCKWXuAdLDexuysLqvrmWgBdKzZk6hd8lhGDEg
z3YJd4fMRnFogVcgesN1ZltR+xw6N3QF61W9lC0fQojU+hptFmFuPsXo9mZ53m/rKkWuXqzKbPyI
RQ9vtYRYH5i5uxM8XfHi0buxN8Ly6e44qRkM6SxHvcx4t+c3zSPfEZOWPRLYyiDutNMCLCBatNVa
fO2c0WZQ69N7EAk8EzUPWxG06SiLWYRkdXWNbMytjqC77UBJWHMSnXknmq4bGieEu95QyfC5JlpX
td1lKsDjeL2EdA90+Z8uff08B+gCbsd86qVcqjdI9M6vodKX89VUyOMXtXyAvFa5SOXhgJGWr/YK
PKuBZEJIqhH2JGgryeG1Xbxb0ajqs/Mvj+CInlIZkRtFlTBZRO1ZiUwX+4+i98swW1s1ANQdXEi2
2plSW0hzGPw9Bd2NQpaDSvrb7qAnwLrwFjqAq99jKs6aeJH7JtQxjFV0ibButG+JAGmVFl0JB0bB
CggBQCLNOOwuWNdhLfTKQ08bi8IdVONwcadl++Qzw3vemhC3Rq3xmcrwc3MpNO8WkTSxtZmTT7gi
AdPn+d3/kvVuGhHshW8S6m1ieOjjpEnifQuxAVfdeItOUoZZImQRZ/X9lc1hJib0z95JPtgjLLh6
CSHJXWjwTwZjfL1lG/IGtqfHvVyIAOE/kUg/XvLEx2dPKJ+01CfgpY9TIAtuP0qnnsiaT37B2MzT
pBqsSViE8OdhiPpaVQDi/o8jjtICWs645r4lgccppErspfpgM1Tp5YFxJc5tJAHRtBPbdW2wSH5s
VUr7rEBpdlki4kdWaMCzPtMpgm0G4KgBQB1JLTnP0dYIaSl/uc2r2S83GzieOKljBleeVt7RMI5y
h22NkWE1X92CKA/8HU+hcELU4pKvyhOc3zQHs/XbNyUoKHItV7SwkWK77AVakdx/DHElpkgkUbn/
xQINlQGvlzmPNAHraOhEkV7P2SQKiSzTdRsFOtP7nytswi/IjyTfAr3BhXpu+Gu0UnUl6i5sQzbl
YXc6dqlbA+bbx3aBzqz+nTOGMovue0+yo3VQf0/VgOr5vZC+fjxZIxlrB3FD3FS6gN5XHDgzmZfm
UyU9iBLjzrYVzanzlcx8FZ4IwmLq0cA2G6Cq7seeBdkPa2aR/Kiz7mXolj+bqM8elQxDbXvckruL
SqLZv5v7Q4jTOorI6pk+VR6H4HNDitWkpI/J3HNKaV2nlXAOq+mfwWmlJQbMCo9gp7CLY2sgLrBv
DPHi4fdMyrmKBjeZtNtfK0KgyxauN9U9ufusbQquMXbXrUb6BsfGmj7BqUs8zP3+9aOS+W7Z4S9x
SII8cONRk0Z00nlMKn0Uz3B9NaDTiRp5bwuyD2azDNuUbi8mlTT84Vh2AG1isQV22hwR5jOMB4Ay
C0ehHjWrjin8Z2F6/f2PVN6/QulZaSkswQUbqs4cfSZQYDzFWkip7hAi66Vhjo6gsuCUrIHGDsZk
pF6s9f53SDdaih1kD1dwnfuhTjoO7Z/1qcTzOZL1Kqh+zombWscPDWLmE81n8mDHT7mm+lmc+dR0
p3KgdQRh39fQWJKY1HnxsXU5r5yuv7G7BDUzvVFBKbgyVhbc+2vREQKAziu9/J1bqHVFkDoAOuh4
QlrhjJhGuFBtxe1aF66mCul6BwLOvlYayToSlDgB4wKCSzFgmgT6eCgI2md0k9KpqlJB/PB/LqQt
gMHA5rBaMOrBsyMIF2MRNSDjZ/KP8Wnproc1mPSX5/EqR0PVXzrhutg/o2TLlM0CaC4hgLm5w3NM
0bU2qXE+kTSCZTL0VfXmhYTb4Wg9MtrQ2c2c193thbq/ejBJFAbRxFWrfzIPwoAYvRbpDYleqXVW
GGNDV00NmVzG+1hvoteqCM0ymFBmb+WrjbGMIsAQSlu+xgrDbt8z4e4GGFeDdwtO9mMVQv5NxMNm
+CRR3adYu4IqhuyTkz90c/pMtID/3Ogvcwo5CwrtQMxgoDfQHPc9DtYIjzT4UvN1BD4eN1HkRiQQ
A5QYVNyvhK9jD91jZdEcPmS45G2duwWkJTSVUqm8PPdb2xZIIV2EbXm/QJe69U5Wecem2QV83IVi
rSejYuzwwT+d7DZ+k7ymKvP0SR5MxwlefnYGl73yz3+bj4ENQpz8S5FL8pey2yCUljW1FANIlFtl
HOZCL5zWC0Rek5+gzmbLR01LSYj+oOtLbJVY7sivUgQ7MBiEEARMmtanzN3JUWFpRHLPadSRrdwL
C01YXaXnl71W1lJ2ySNXe5ElylQKmVYjoAE970ycVjsyAQG1j7tGiS718wWaTSeHAqWyJ08hi+UA
JIG6QWpdNyqnweu5uBbNtFBojZRvk4cIXufPJhNM7Azm/v0CQ+seziu5y/FLDnEctZgdhorKYRpF
p8zvFwegpyEmPrCsCIL/qh6k/RSZocyW7vDbYpkuwt1hxNvbbfDc71rZskkEWP/z8rcFGFSpeShE
Mc41oaViTu/KNcA2SQhYuVnQ/aK12ZYQR29WKenCcxxfKR0wSy1ifNFlVCMPOR3BExVHcbzDq3CF
/anPg2kw2tFLrHGVahl4OCoW+yy/iySSi54OntN+2MENfL0Kn6PTI1BvzL7j8Bx1r8x7m9A3QNAW
LapX//z+Up6hGuXwYYo40KrU3rDC2FKhpWJl6F9uQKs2WRpV92fL0yE2m4OV741vWhDr16MLvK7N
75ORxI7wNYt3ruFsQAQxVoA6AM9VueRUWTxvl0XaWeehDigxOWKeZWIpCkmqkzixRDmsDZ+X6+eQ
EdtRdB8cUrUmqG6Nhz9T3rl9DReSfwWnh74GfeHCFmUwcqjwVHJrOmqUnPAeUdynDS0PNj6NAas/
XTCIGG85X1orRh0IEyb6Qki0hoXUsebsHStcG2e4DfWpHVgadXdDfKV0xstp3n3i6IP5og0SOSiZ
UlUJ1Vu7dlrmzqmrRoKgQMnCRS2IUI92WZ2dkmQmHzMQAL/F2P01wo/ifqFrVe3Jj86pbxpeE3pm
gsupPJmPzL3XRySb2h/IbdA53pJluHC3cHQKt6VMLMwZIE7NxTpX84nzRy1z6O06erQAS25pHmVo
CRgghE/y4WlFZnSEg3BvOMU3b/rOx3O+hZbi2cHWsS68LOTkEIYqgia5NfhXEDdABy9P1Qk5cdTr
ZKjr1Razt0NObcqcjZ2KFTv/+xeOL8RqhgCnUKPECKWWr+S6E5ovokx/1HFqcjoe2jAPrmWzF4zY
OA57EVM4aKeo1hJdof3qkRPRl36KfK4ZyUrrb0YAYD+sxSdxsIiCaLXeSIIOBkRGFwSewaAQtHZc
M9yol5lficib2jMTL9Yn7cvhQkmTYB5T+7SfVrcGMAR+fRbREmXg6rm8JBrrubUc+EptZTpM+TqZ
KBAu3Cd1bBbo6lERr3Fstntdaq+gM78NvXUATrGy4ptH9/FnvOYEW+AF9pPCWgX75xh4/PplhPKU
A2JBkJtR6CV9zs+WZIu3p6B5EUBjXRfhIZH6NkPctmiKPY4wA6CcoEVAEY9fZyubp/HKDLxg40Ra
3Lc00ck74OAXjEZ6W17zn662b+oMU0xYMA59rwKqgvyBXju0jydfdPTw2te8jFCheAU2yTBJKh2J
ePF+sRYVC0AKhrAj99pgrsWKwu1oYzbeaU33mKYq7522YjLLRjgB1Mlgz6QcUXy9ihYxftsrowH+
GHZ5WAyyhIbRc1HMYZUh0cH2a7AamTWyqXt7l9ZfNM/OS3mkLb3eaPQMvnNmj/t3pSW+UTcxSQUd
FDs5dTw+6ZP1KLlnK/K9uXsxbq/5xTC54WAml94mJvVyZnWGtk2JfgYcRDxnRww3AORJr4E3qXbO
gNspresYSjOgCBnmRLznFytb4b39WmYNQQw3KH8N35lkrDtU0BYmU0V/fACJJzV8H19H6BivoQUx
3RkQ9mxnrcIRolB8jWWkqXtAKDx+giWrT4PyBi3kTurk1e3W9AphYmWKHy44y3qzcpxyx7Fs6ZJp
vEVDJYw71m+k/Ba9MT3SyizITuHT5N0/2UZrO5agqH0Xq08UA2GcZMYb8uIeupg1wGjimSVzZd15
iP/FTyGOkn0mUfnc4/HOwy5mUmtMnNxiKSppitJhrmxq64lFkkFLVYAg8nqazvPDW7FxJ/8fMasd
gfpeAXcZmnTGG4heqXiuhASTzOkPjlg3iTmLns2NBXjNpxggrTshjWlUPQDLCqcbC6UducPgi0nu
bMR9wAoDqUZ2o0Lj+m8gJqE0Z/B6GZatqLmnrwEgDtzaPBlMLgshkC4sEUzS0QLjszDSFbtxP8Yi
VxcBOUtaZTLfuPttzQJHX088q40Rx+ZHS5wbdmTX9rR7voig91LC0Jr/35+K33eBo32rQC8HbuG0
IzuNXBID8FCdUJ/gdhMbPMBx6PJm8hqEoR8S3l8ybaHvsfxUivVbdvfVcNJlU4L12IR1f3hLuQT/
c2mz7knCHzilzaPLnQVRnpBa++2Isa9JlO8lvhtlOPcT4A26WdCov8wKojpDmd3ahonQAoSTNiBF
P+pXlUo3QH+Ui1DW0+6jYc1iuhS4T34YP2Qj3dGklUDWwUcDLINSYOLJi2W1KU6zW/64l5mH0yZ7
sPNcDrVoemHW3cC9JXO5YCKUGXuZmdge49m0ckfoaj8V8iJzqBL2J96yC+f8jeaT79iDSwxncKkg
TgdPlGMlPGsEAKtujB/Ku3KdryIedwscif5cSLm7v/4vMZgi9+w9sXSZGJWMRgu753BBqJ2oqRjX
h6m9gWYUsZjJ4XXAS5wOE88oWw3QHrkpFd6fxBnZLhffnB3+ojpHyJBy2hlIixHWNWu1P0ZgMrFP
SvJn56m2htxFvptoXjV0FOQSZ/IhWIeQ1mk7fqr+6J1aaEqH8Ddcugb/W/X2JB+Pds1hK2EQogvX
YEW7OnrK3rUzoac2p+xI6pSIg4YxM/mAH4WkGIXQRdaDBa/vUXkX0FoMUlkav+bj6xMn1iSeME4a
YyncG65IcaMRV+vt2OZENUFbVe8bFZIZ5SegbQ2lYGkSQMy8PCKZeYjg+rlv4UNuBlA9KyuxdVg5
G53pTq41t4VX3fd+/koYSZKjUYl/uxd7+zhkT8pBB6iRETfGSNyz4P7gQri6cTi9xHHjb5Ytu34K
VJ3IXWeIXgY6L4rg3OA4Z8RRioETZCuHSgWp4/c8vEa7WfULTkk/XRyf02EDpMD6lc8gNx8ihzLg
XNm+tNG5A/+gVIvTBtSLdyp84U7PcACkWaGJ63r5U8n3YJZkPSBS31SDlyhCoLbVbePeMyEpomBe
tOWv9YMRhIUprxJhNmMiWgXtw+ky4jX2rFU7UqMuw5pIbGa4z6qiWkY/BSLIGRH6V7Y+j7MvLHTc
ZASlvlgzsQY/Bj9zIi6H27HEkXoX1lRJmwOQBpyH4nsfGRkd9Jlhu+6K6Ye01ap5N2tf58x6F1mb
kzIuWqLl9IT5dEyapLKLENmEvxfNPXtM7ZXw/6Yxdws+tLGsVG/y4qAa2PAkidnmLmsxrVKSWiVz
AW5S+xAE3KTd3GJ019Y9M8JgFKjVIgi1DSMFREOrcuyw3qEroZsY6kLN9EvCHh6kobCz0nwUEQOg
C3Skg4mEJyzph5vqhYejFMRXjOxYm/xLM6KUiPor+BN1PUdHB9ImN0nVcuov5nNpvIMX+zLS0B0c
IeTb2q9r5yUi3xv0SErjnpA7DrWlZJOYu4UC4NM0vKvc+LpbObbI97S9QMW7JtT9gGbhIdXMbjqW
nxNd6ALZbRQFARdAYqWz4OTLDtWABFdcUrORpwnz7rtDGIP5wTOOwFG8t+O+wHznI2YeNWJ3oJlv
NFjYxEyvLJvecuh+CUwh0+t6xhEmG+jYQjHHOa2sBUCm/r7GzM2uaI0Dji4ruCBH3SZJjgTJyRwB
hUhUOwVPq7UHKcram1gYNH9O4vr2W+qA6PT4vJ0elAL8c60eDQsTqsP8ycM7Bin1/+jUHSNp2cYW
OI8tTceTu3Jfpk/KySFGn9n8dQ9l7AuEnGbZZr4csd1AifzNQmYAW7eeF47VsF0KNCR/uyuy3DoS
qnGvdWANxey8GGcPzNYyvQ2ZksA/w0/OB7OTFKkJUGDcp/iKRyWz807zqAWDPYIsU3+aQvB5Lry3
j1rQORHjahE8uowHFEKWjQjAxKQrbbiPzyzPRq2R9RxhmIxgO7NBvAKIeuL6BcF4P+RXQNnuAGEF
eWkADOaNw3ViDD97ZHVuut8cujb+VFehAMCEw8F3IcP7oc3Dld5840fvwFXqv3ORPDCZnvggBFtA
0SpAwe7fxCPH/v4R8AKD7EZz8qxgmjsxlGTeHF8jq+UGA6PorADCtfuiGDzMBqtm9vnamd4oIr9S
ZADLlyAv55ORwdw4K84ST7cloIjRa+/5OezN7J8cRmdowt7jQW0Op7rF08QevWLCKjIHqNvcSB3F
fotdMxrjyTVOGMNyhpfyPIEUfr4gUtDDsYaNk+6iwR/sGGLd4ZRpht/JL8BziUZc0Izl7UqMRIO/
jfVUEDDEyepHDshDOU7AofrfiSiUMBkq4OcoMdbGDZj2D7PYTwjIqgUX5NO/6LjAziBE1vMB7E/z
8zTUIgL51VgbAklkzIpkPKPbAgcnjq7j+WjEmqqBH++Sfwisg2WbbIo2HwWlBNz4Anpv6i1ke9k4
jgx1pQLGCUDMzc7wxuRFzkIxEk2KF9KBR9AdBnTq/UHJ22r0s+SKf6FnZFCWUQZRaVSbrMNjF7SA
DLP4Uxt+jFdTJJMEZO8RT7cD/W0t+Mg2dP1D0Y7MIYH1T3IP1qYY3HXXEOpBTQ8UAcZ31JbRJIFB
FEkRCpKrwXqW4dh+oe4/KqlMsjuJME3isTkwwX986lF5azskPilbMUnE/8D/jyj8JeoFPVrFmJnQ
3enfIFXSjeoBcW9dUBEbNrcjVDWDMmEMmsVwlGB50y9yJXET9dS4lte/KcjpdKJzUD4A+ijK4EmW
jYq3gEy6J6k0w3RhcCScvA+wDji4yaGC7tKKJ2fPCExya6DJtxr1BnFPHZEQoP1j8rP6jpVGwsnR
/SkOksXzEwP0cTxrlpf9XNz10wAelTGmvpQzb2QdpZ82rEqJsb8foEyefkdFrI3fUUjAgInYcC0d
H+Mpd8gPTbuJu9DInnjMRdzdhpFY5u9XNYDzw3OMxEah0yxpJyUCQ21GhPCQsDiIz7CyIkKCu5TY
cH5aXYdez+/KxOGyHD4jE81qUeULJmIOikQKQw/IoWK2/n52YpjOkxTRaZsNnNKzShQnYqBWXvvr
ZO+Ve1o133qn3JwkBm8wJUWicOVwtyZs97ovjNV5qUcq69+rZG+7GE5uyUPRc8y15XQ68EeKMynb
ZQuT72uXgOBy4JEM799UMug7tl5NaWal3e2yuaK0w03/qU26NUjUvmy8tczdhWRBdgWkTfSVTTJF
PaKKmBwNGYZP/MtII59Q9cA9Tnqrn2qz6/xkTYKTvLyVpzi5nvidftWEm4DThyHr1BGmZIhMI8/I
ykYphXmYZ6KiM9KazwN2W9BUMiSlijB8DRx+Zlnbv2sNDbmO5LJupkbTLS/VBhVsiUAZabGL6gbb
NeugmaXGC4yNr+ydKo/p6gUHOYbF7GIZIJEOQkuWSxD621A1Zib0e20kQOXWqnXuDHd9nrI+7gV7
p2WjoTYiMDGUM+dXx1MQGHJ38i8c86KIB8LDMFztsk41FA9J0zvPdz1v7R1p3k51yg03iLsgXoGU
TrPxiXsrRmgOOFFHsml6Qyeh6lnOL5wLQG4a0x1J4MPDuFGjFHnEgw/O1RMpGoXD4cK6qXzurMYe
0JG/NuTnr+lheZ28PYsa1aJHbtv9RiQNLxfDk9Xs4oIIW+zyvwDMLrdYivBpCruOB1TMFnNuiQ83
zMZjYLWQNDDwnGckdbFaejPCnrHT2JS6P4QHsG8iZsByxgF0SLzJ9zDe35lCxmqfMUcD56cGCUK0
SXsiyk2Qfq8z+N4Kbk5hrlCU+6wjAVvMEnJlwiqRKWVWA3b8uTZYlt/q8869BeVbVqoNn9nPHInx
oIi6nyJBIiEF4plEcjPClFclT1hUKigdG257mFAG6pZagcHH2v1+rGKfP64TOMI2zm+7REWilWqy
RUGjrp2p/CXCbz1NPqQEle36EzAal8ptcdg6+iZJcHtkPnoTmuPomCFshu7FwHAeij9Hnvp5KvGv
wFgErhk0Vcj3zea99ugEPzsNUDMouUKnw73FkJ3gdxYNw7ZyisEYJ+dvl2XfMtW7ZjaQtpe7CZpL
GJQ4RLJ+qgupIC2pxVKHgv0H4UtPgc7l6j+phynE0pCqcRsh+7/Qr2os6Lj/5IvMopBqWN3Rg4Q6
5jVqz9zB1ALA41Xpj1eoNRfoUX8y4/oQsfY760O6G37jLodrc1HDvhMldIxqnJ4M3a3NFg7OtRql
mKcF+GlhXeAon6X21Gxk2Jyztr9ODO4GiltzViMLCxJgWxoxHn9dhRM0jXlpHkRJ9Bq/bl3uPd6O
ghrgOtDE7AqVOuZjiC3LbyW1zAL3Tw1k/Le1mAuZpUtMYl82OZ9mzjQZyjfzasrLlXSk6zV9M4lQ
w8ZKvbsy1NnGfreDgYg0nKkjvWJgZyaRpzEg8pfwTkhqY3prAyyWhFvGSMjicN8qTDgabTRvHgkf
TilGlePGjF6MOjJjbAm+x05wmQB/kTnPslx65PuiGP9DFrALMQ2EwTQCYLHgay7SuBw4xgOeXjUU
6iqRv5C7yTwJ6AnbwCpmpLx3lY/boPw+Lq5j+MTHZidXspZPY6VyeAOSRAwVY6ap4dEUW5qNBsxn
AwkFEsSDMzq5ZEDcLWlnQ7SL2oDD1el5F5Prkb7zm8U9wRbx5D1ufur64Qt3E2dkmnP0smzgFXAb
Hd7kP8PFRKXsV826lqBCQkm/30RHv8U0grK+85YHCKfy+cDFpiNgBD3Y9cRd1Bzv1B0eVMoI1nRo
54YrNzyk9wAn3bWpOprKbOtlwFhA16UEj1V/otQd/IbfTqy65JJD+AdsXViLUrdDHFvKcb6YeWZI
lZvY6Y/lNtKegK8km/bwAeEH6XFpWG6VYXqNfSLm/UpH1nCKV6lpq9/IHpQXI0YyoeEhun23uY99
NtWaNa2hcjSINZI3bPP0t1s303eHZbHbwukF7vPw24+a6vYlK302OBtU/6fSEjxR1K9QjkC1I9FX
qaqfpXUeJRMoD61rZlpQ9hcauFAyqHC+IQr/KFPbkb/2kmv/QGf8WwR8wH8DFT82R/XkikPe+mIl
EvfN+OnzzJKLrh2YcMWrWJZj+mo45I1z/veQQ0TfYDjVkPJn3dEISrYPo83/EJvrnQ47KOPvbGTT
F8yOmQ37UdIT1r+Pc5MeXh7xsrwPW9oud9qiBRACKlSSAIvyQHPzW9AUmOT8YA/+z/kfOiId8Rrz
8rLvXBM0OQh4ww8EnKF+d22EpvgDLr8F4PippPSGN5497vGZ/jTmWhV9DtAmnwS89ppsisK6y0OU
7qp5QAjwcyZiKB9ZtyyHw/6DgXx0XFskQHb+rHBogMBRMISqK1pX43aQDNHtFzh9m3gP1LrzEVo7
j3B3h0vu7G3PI2G+Y7t4wZPjGo0NUuQGV06plgCajJRq4barJxLpmeEdT2qwJAjq7AiM7Pi5m4yP
lbQ5Yg5jSxPEPPNnhk3ZB12RL/jdAqgkSg6zquUo/ZceZyzA7HFEXb9b3TxHBiZuS3L1p3mq2ib3
CGcwO2EJ8bsVzZ/3inci3hCS5OgKkKkzPeBZGW9ww7e82RY2Ibvvbbn5XJQptEK+DzgEzQUZu/ih
Ul/1BR7STbPNkEEN6n9V9uFMKpLE5ocwCE6AciCh+CyaPLXcxh+SRSNVD+lJUzOFBxtJpoeu8FPQ
av75/EGTVPuup0xaOOumjrrr3oOewhmeC/GGZdHbNReCDkB+HPn3d+bUuMG8lwTH1WCn/uTgWJXV
nANn7ODAsc2jX85sELiF4RS7psS9qWXOOPqLQyC3+TLbtEFg0N47UoSn7/Fmd78SfXr33F0sfIf2
Tr0YvvWxCB+XVYFdmWLttFV4uR4Sqp09gDM+2wQTT6T6CGwoLcLWkWsip7qJZ5ixyOH7hwQOmgVK
BdEjlj7M/8cZHufmjsxP4gh4N+gfuCUI411A9Qt3s6r0vigRPF9+fbPnHbfLjgqihV1X5Cx/+l+P
89zoab9hhP3xFduSrl7GMPgt3pcAyGRxSVQBmYZlWjgP/2qDaC6uvROixLRO5K7Iz8GDY5Hlam24
Ebxb/NlCJiNCCkmJxloiYrz78PnYqdrUhSkDN0FT0W2c7xw74D7BC67FEGcRs1uMjEAXpWlFlGPF
VySh4AfbV3+hnn8FaWgILSBS+HakqEG2JfxoFVosq0+UJEml4grTSS3DKJN/9UHeaI9UBVsbNAC6
A0PjFM5IdrMGsxSYnGCcD85rED1+vY4+mNCuANj3veiXQPoj9+jQCMYV0GsjRSvq+wXu8HrOjcWV
CHnCh2GMdk5W/et/MHj7B2dNwwEW+LpCj9wNvrcfn7QxT9TUwWVi3yaoRJnMfzCyX/3/3uxuV36M
/r9zkzDLvj3vsjx4WZxke6v+9sM0+h/XG9HdwHePr0TSJbwcwOuIYWrt9OPz4AcfyaCfQEK7uS9+
7d6Yky7zatRyA6opfQ2Wku4QV88YodxNuHC8igsFCFRlrycDmds0YS9UITof1VjUhqmWJx+PO91Q
3QG/aZ0pDrIbYi+49yqcZco/IhJ/xmzNRcGmWq1+lvtaUh8YHU/82g/rBoi6NYxWiT5RToKeqtBQ
VLqRa6UuMNorFddOWg8de2m/z6UkmQoGogyOBfbkytV94kNVpPCUOVKYYhB6Wxy+rhR7ND5O8JZx
BOOGlToPJJSSG3pAGfehqF5ZE7qqiEIDtas7BFD7dvmc6nX3YTj24bLuGPtP8hPxQP0l4fSW0Qn5
qJ6tNpkcaDciUkQcAotZrUBh91kB/I0PepKppY8R2rl8CxR7OVU4tCkqNHkSOLxskIF7PkLzH31c
94OGRrJ7960p09kGmZi/aq41rcMGTuqEiI0mCCBbtiIme3Y4hoI4PS3iepLB0HXckBu4D8WNq4Kw
huLr3kvSvDuCO/Lp5koDcB+WgLWqppxdB8onZDqurP7HQwFIx41uDlocO7uZMH4ArBdWytKyLWHx
ynfo/XF5lqGg7OFKjmZ6FzoecIhgIo/K+Qx1YfoVlgH6CDejfl7hyUTDrTT2mFCnXxu1FVJNWOYt
3TgHsTLSuVT4/qoleAdDNBaCh9VevrruvPYfaVqxIuF1njnsc5N9utw0ja55OyVwtF0jthSEKJFZ
psz09VijLtpj8JsxHHlFaEDM4D8I0SwS/FQkKEwhDpH2//LHje/yVhf0JSoyUXpZy+uS2NYUUxdv
mfnmnarbKqk64TCKSc/hpPiswhwbxwhVjxDHfxo8Qq3TtQVvIpPZe5OIK5Hf14L2h6u1bkGI41lc
DjJpQHOYz3QRgGSQm8sLZVjXxDCbI3Islq6kFQwSOjfTl/R1GTBi7t6fypcRDpcct5zac2gdzQVm
tKEScQb49NJeqOuLVF6G0OABKKB++yXsjXp9ct40ag89z1lsqL7wsMy6GZsKDu383nb0yi5sPrPw
B6oUPfxNUjHo93ffQcxIhue2avsGokLXGK/61pAdsob8bB6gxtGL8JseYHRHhEnKyuo3QmUzK53f
uppCQMv66sw8E2eaegKO2HBWc2eDNBhz06q3p11L85Pw0qb/LoscU84lhUIGg58g2D2tlN5TPBWo
8w9xHnM1c5LFsOFXxg3NFz85j8hyyNZHxwmkcYNgnZMARMgssM5/VTJ12CJkvALaNpcVIYZszNsS
EOQ00pRilZtxiyjlV3jgAZgm96MbDzIPiqor9i8CyZ9DnWj2hP2/jXFgBN9ZMpuHxT6DsltGGvJ8
5pE7eXv/5wg0X5fP7np0YiB98+bVbC15H7IW3Lzg7/7wcVsGeI0sNvo7jTBwD7xnbTJhNNGt9cav
n4bpFxB4eTvimxl6n+TM/yI3yd2Szr+uudGf9b8iAw0dl942eXGcGoiAQhA5e1qNtmEop8RVMkL9
MigHu6/Ht3Ne2cETpWDOPACNalpgmN5XFktUXiXro4dc6SYRoRA/T1XTEUEy9wVzn5aJfOFi/Ghv
5p/ny5RcVyR7voOYyrSksf+u+k+9343/tKyNCxOeBtEG/55XO1QLMizkAr3i0Ib4mSTiq6Xzi5f2
Ig8q/rQTMt7N9Qf5X8GxXp9Yk0NuQhDRFQC9BCPg4QE9y2imnuQ/JoSYpWgTXk63YOB/ECSs23gm
FucYEVxCIW+ALD7rxU9cCbklIHb1Guzh11Imsst2meVJcqfR8sjRISUI0rnppc93cDWLbyP1+8j0
qwKwXX7sMra3ZaUJLiCL0Qam5CR+Fhxhgpa08RFmd1dKmIffU2evAi4zmnK51Iq+GvzYyBpBoRW6
Yeer7pzWetTeSigs5qmjXqZlErzrxgYoM8UvDRSOuKrQ4roBSZRzaRfx2PJRP/ALu9y7UdZi5Y9i
g3VZ4pAuv4cNfSeZ6sBOplOeOtzknJ8izciT23ext3xaofMto1pIs9aIzvRv2JHui3H9vMWENHP8
pcWYKvHknpTS6heHIeYjFDEat/MwfTuufNl/2+N2BmcRV5cFjKc4nbOL3eHTdNff1dW0EOfLB6Di
DFQ3aQRJsmoZqEi10/aQlV778vFE2JSsithjf8BElABk0IjJ+jA39aE9shWv7vlqOZ6XkSGMSqiC
xuLsCV5cHYWzECHzbgwN5GPT/iq23vbiCTIpgcEGj2mfQYCVVmmNsWOm8om9FA9qs3cqyZT5dp8H
IqZJPchkwTXoCduvP/JobtZNykFgSSr/L5RGwDkK1MoaCwsBNaVr87/CdN23jSunOHhrZTQONIgW
ZxeUqGGiH7bjtUQOTtLNQBeYKo/M9apqrdz0hU2rEHL93BpKgEbLF6qMcAzJvXuJe7XanENYUioA
6fFNSXNHTeh5K6IcDgqxYlxw/pcIE9gJVbGfHQkKjKcFtavIL3RuGNB8mIHAOBXrBMKFyKOxAjZU
ViFMP7TtGxWEsHi2/KkScjdBwO0en0PiqSTCyVC5eEizeQzc3WYzajtvXHVrY/tGckeYr+N4uJHG
D9eVEXpC4M3Dd+WsyR6xmuhS7n7+0S2fYPRtxoTyFL34y4rHpH038TQtGwch5Wbw/OiOw612L0/c
GoYoWfVuUM0uFvuQ8TfAIqORu/n/7zB053Cv19wFZDmY5rxniDD2lgB893VhFPL36AMwPa8uwjzJ
OCWpnGF/pnXzHgSNk4XPY0cj8H22g+6ybhfopS2oFfUzVCvYpVBUGIC96ibZZpZoHBvlWZXx4Syp
CtAothFRtR+jrttjOvxdpYxVAb8K0e5rO8NuYseRqTBGIz+eHDFs/ZGdFJiiZP02Ls8fRK0eYWxS
HFVDgVn6QjX5zlJ3pS+D7H09kj/fwlGOlD5xVgHDdOdcXvwDjgvU174k0TEkx1JESUZWbo0BusOa
MfPdeFiMvFi3ozUG6IqxECu5Hy+U2JSSArnurCVCs4HvRXcK4uEPQbOzVnYHbfrioqZR0Knx39Nt
EuvK2bI2pNZQUohYtsuYH5fMP6FFCXSNdFI0VUS/5uIKgerubFPFJW+YA4523BaVwTC8pj486qaR
mng2pg4J6fyXkZ+aa/miQoJG5XS679tU8CP/Y2bBWdJUog8VogNDK1l4S1RKBVz1B8cN7RMGvwtC
rjGjSfiRa+MKmYc84OPs6n3pEBspWx1qrOa6lsHZn/WIEOIwEKn11U2iV1GvoK019PGxRPuCZTDD
h2ULR2wvMyR3I1TR6gM2dorR5mfSVpg1Y1fWy3Iqmp2M7TLGqjZpuzhXiXRmjwEqk/4jup456Gyj
3B4fx5N4qJIc8O4Na3AHyVVaxUahfExAB9bJ8MZHkNDs7YiJaDf93+89MD6gYijVd6WsQfeOXYCG
wkqFsR+n1l3TgJHCsuLD6yNwSSCcQn4lfLlTTVpjMjX5dCudFRKN+GDIypg/w4b9NOoevPNT12XD
NtvXHVm4hsQ2//aC5U8ll2lHUtOFsHJBF+ERccUhFOoefAJ8TGX7C2gBsHImBOfMl7qODlMsQuut
haL6HitYXjr6P7jJOpFS+GphPa+f51zMca7Ugdo7oDNMPbnvmQUpF1Tq6pWRz7rJortesS+uXyji
a5u1Xk8xz8cGFpzgg2IrhWu5fGtv9+cutr+xo0oDKQLszcYYjEYEEuaN90FKwl+SmLp6uGJgjYFM
ljNMOI7QMt57wthiM1zOVAmWeaYCf47hQBdtLsrUosk2ZlqXXADJirXbNA15jMitBHhVxkhvd0zg
Lsp3SQ+sqG2lhXpO+Sy8lBHA3Lzzuj5tWHgyDCksZqMUrh0NFhLVw7PZXTVU5KhPXAEf/MGc64Ts
wMsF/Nqimoum5ntcztHGaAztwhtmgeLzXFplxSIAchvyIz8Pjld5vtp55zrjrlUa3m0SrS75WhhE
yPJcEqxIszpll6kRAZ8GpYZwKw/8SkCPJiDxb91mtRh0mOTX0KWWJbG540kaApseh06DpOlgUl1P
kDe8oJlKwhkLxhO9EJdjEOatIlE0fsOC3KAQpoiidNKmgoKocr910cg2+/NpfB6nnMYTzjOKZWUV
JH5s/rr930zBbwqTlXGp98ShDntJPGoxzh0+lIx+t1zm7ziP8RdUKNjExwgdGsqh1lIxBIMWP5Ls
iNQ7aFmk/uv5azpOFDI9N3y8Anty1nA23rQZ8Js+LYZl/QAspSSZYNVkY5kTAY1FypYEaboLDTHN
344bZwfaiMV6WkDZwM4V8JO5tihPrHdYOFm8VWpQHuLXGAdfarOXYvXEqpAU6ADJv3yuEdhRNibI
/sDLaLeYslf8pha/tMmh69avsCGuq3UBoECzbvUq+0zpWG1LcfMm9VraxpuTsXn3I7AgufCIvaFv
H20EjDlHX661ix2uNvqJozzLVWh3W+rZ409WHuv7O5aXfbdX8uG1eIEyJDFWl7WQ8r4VhTQ4hDWd
dOPdx8n6/MMmSxvfT0F/DVfs2SUsuaeL9dJXnmaWA4shjeyvw3NnQDW5+2Nfd7RmCOtwWM2LRUkm
NwNSY2VXz8fuPbIlBMdJ2pddSUOvWmgRwsb7dkhPM+6A98/B0HuiVNgyIT+MDrt1+5qjdB5wY4ox
Gc5ZLJc1rFCK35SjYp8uG7pE1bvRXbnZkAfnkYfv9os6qG9h0rebUup4fxiN7+/PTMVHVi1pjJc0
RVBk8P1nfUiIaKH0CwgtdQr9EY2AJWmN0SOFpfAMWVTqhacnBBSGG7TdYZ4sd9SsFahVB3YwM1Yc
i94rCTI0DtOEEyyZxq8HAg3U7QbbT2T59BJ4hHq8KJnEZoBHrA2ubp9niWyaKAqSXcKELv33qBdE
/tUDMoQzTN7zD2Sv9wnlynWJ/1D5T5oce2/ZZ3D9nwrI+AYqm1LtlsF6e8qmP+4YdfWRizJ23TDs
quThS8cJEU7LJUFF0Rk9DXMsrevbSUXAOLZTn0wFQb32S4xIqc43djGv1ByJ6bmum0RsMxILwM1O
GRcNltYBOVC7OQeLtC4EUnnkHt/uIUyuan+nzGQiAXeAzBAaKp0wONHrZeVvOawCciST2eB0BMLA
RI77YrCsg454nXNV+EAgoV/76/UZ9YjAP4mXMVjahTqmYFoEfUPWcgRQFYcq1oPfuAgbCucseYjA
FsspqPkccWNVCMAtsF2Ohe0hXu9nouX5widA02IuURaW3cAQemy/C7rHiG0JTBsNFZ4aknyR+a96
uo2sVfNa8DnRXgjedHp8XGitiBUzwirli+OmurqG7neu7KFpXRxMCf5n6iRlZy48MKskuGE6r+jc
AoGAklzkvRzMTZo/uyjG2e94iD7nQ2BgSZyobA53F8y8dfVoDnMH1QondPj7bY4uP9XV3hZfr/yS
f+qtMGFzFxmNuaE8rzdpYM6pypOUBOM5LmTmjbGPfFC3uWK562zzresG2MYWwT+9kqCWCJVfZYQM
FayCwcum9n/uWcSUVjjpkejLAq4+3SwI0gvAK7SgfgYZIOC4aRSdq6RxfzWwSs612e1eav6HzTJB
o5fD0XFg0Uj78+ZL7U3JL91cIuo4RQSBLMRS3pITxhWu5+t12Re5ChZ92BxgybYO2JY+E4syYiv/
Dd0rqHSnaVKqzOV0rFKp6eFmC1jONtS9jsqr/pV+yuQiTvLOGM5yHV2iPkob2PRVJUrTX3m1Us0k
w6jnT3bnZgero3UQbsBb7WnP6yaaG2dP3N2tZPXVPmEaqzZv7vNQowJptwPlypRxMJvt9wNGfxB6
aEudbSWqPkF2gxZ2R5rEbJnbjXgq/a/jUEJsH/YHDG2KnTAuGfq7NZ/cLy29CwIeU8jcAV1XjUp2
+9M8WpDd1qTpDjeD7v+xmrhqoBvY72vY3c0yuckwN2HHvTf3EkPXEP0PRZCoSBq4Gqf57IdDkzoq
fXWvNTJ+iKy8IWbmQkFwQ5a44bxJUySJoJvQ2Uyc2IvlyNXsoUkkTxZPyZCUKMZ/Qy6ICETnzL3w
Slo2/rDQ3Boc+sY7aTYX8HvDPdQNUobhSkczAQzKPX75F4ZDuSyEmCufUhFu0AjmnGQl5/zLeh3C
NCiqIGEjgKGhzm9GBwizO4XD845b0T7pYNWp5SLkh8BiXWN6HIQmCi1p5oyvLLvotd+FBy1EpewO
S9QDkX+DUAUqhRC1adhNBs6Pt+Aqu87uaAiKHBB71oaOEVM6JYyJs1ii2SNdHcp4Pa6rIfqhShVS
54t582QdW90iPIHWAlkIz7WKp6VN4uj+jF1MvXxyQM6nc3Kpal6J2hZJQGkwErq1OePbWvFjalJr
THsaYg852EeJ2Fin3Lxz0wEs3buPJVZixHdwSpX7nKReUGsQHsr2neKd63kpS1NRqc9QSliiS9lA
6eRO5pT0TEJCY7nyXBmGEcdV+6dJRPKwVsw8QKvSeCt1BH61ipWuDoDntuPMMY3zD7YYkkkKBF3a
VmJjlXUuszdbGC+ONz3G/nGPsjYP84rJxQ2BI8DpjdoHYtY7NIvpqdWK2PxDYIZOPtu7JpBcT6A/
7IphQpUgq4tUmHXlUhCSjZ0bMMPGBdZWGj47KmfdL2iHBMyre2kYIjEwd6xuQbudFymnpUGKfXnh
HVmQkMDLe3D2iGuAzIF2GVHe5EYNtq3LTBWfk9py1LwKKCup+qbTBwnrIkGQsx2kpr7cqglinMrz
a33fQLx5yy85Pw8b6HlycxnHg1H/9GhQaspxZh6GHbWpqL6BnQAlkkBzXNveSaEjDKULc67vNEqO
AylVoA7tROLoplUkaCgRozi4Y8M66D1W+roVPGi5nwm2J0eLDuvMMk/GTpDW4k+Yt9YBm8JtMAtR
lbN7xgIFXUVIh09AjgomXriKPpQFgpxAzLMOm7JxiShkpXP/ZSd8V0Fbs8z7bd5KAEnqZwvXFRYE
UGk+b2zNdvMRB4zj5jhzN1Zd8I6LQvdjgH/9t8v8UFaSb/O3oR0H2tJShKBPjUZ6dBOxNGEuy+GN
J9aB3Sh3LgkLQkKro2HIfAocq2Vs3yVrh9BqC7OQsXsuub49v71hLOvaGeh4JqonqZGD/LTCOAIn
Qm/cJTGULYvV5ulNTo6f8yqqx2kK8l0Kk+N3wFn7ZypgwKm1+4oahqVKAIpIWQ9Qbb9jRYSRbRdE
sla+bEe+X9jCZwwLAu8VbjytTshab2NIcVMKiLgPrQ5I/kvCvWDYdmZ64abz/oy1FWpHoNbqPDuh
U3INPc35vevJfL847l84UUcJXEormTiEKdlx8P4q07KTXajjSyYqJcO4HEyt3Wet3Mfyhtx0fwDo
bthiHi4+bsF0dsev4zQmL7ZaKe1DoNqSMW1mad5Xtyieg4hUER+0k12pRWTRHyVaIb1Vx8TlTrqh
OV/ZVPVGtDmoQU6XQ365dzmVLjMo0k7Kq/1cWaef0SADbD8/LriK+MiGG65WWHrAN4mDP3ROBJgI
ot55uWGAR8/o0D4cDDPkhadcKpkGkT4nXkSDxF1pmWdi7qB25rEj3yDnqDWZoKpk6gFQb+Ssnarq
UxHDem1y2z8ckgY9TY7JihPHGZ5yhp6xuXb1yh/Hx+aBDJlorCi7CCOXSveTUqEx3OX7sAR02zMB
U4K9OCZvb0QkToIs2nEnso7zHSmVKwoOBcbMLEMmhd3O0q0vVpheoRedbUM0YBAHI24aBkPcLs1I
av3FUqAKBx1W/LFGtMce+SPCjeTVLQO5JvxfVSfIpnxl6N/YFF1jdbcTE8Pm8EWKjvola7unthCn
cGfbkY10TYZiiRDI+PApq0LESI3dyq1tQcjDWmomdaW4OUFdTz3fZmXn+U/4fo6eWv+t8DfL4lCt
bGblfXuk1rum5Ak58nJbw7AvKjkxMKZGb5UcREAtI9CpaZANIOb/OzxkKDL8rJZRWk0WPmGNI2K8
nYS8lwgi8O20ZzBOa6HhH56Gx0R9sEH2BcW/gXPDFf2TZLin1xclCooquk/myKC3ILNmcAk9/WOb
gIS2qTh32Oj3mbfx6gnr/XVl5u9RtUyAlj6N/isCxEvk/zcF47Ph8GeWY9PnWw/q6ncYeKI23Lyp
E8tv5yuYL5p++HKX1B1wpJqjH540bn3NpgK/Sbsry1X64D3fbFJ7DDiWaVOUYa2dm00QFRjbPQpm
v6sRf54rCzC99MozIcHYQm3FFhjcPxYxA8lwkSJ55/rzn/BHh1g138P+oDtvVDtXV+Ildnfc/UQK
t+Z4drUR9Ajz7V51bw1JLQnUi5uIjW97V7dtR0Lmtc5uil3ro9BUC821v+EpEjiCcYtVcI1UE+lO
emGCgbkAz6tdYELCd4p0d+kZdnrQO9Aie5J+uvT5oVLA3Vb7Wy9Hzzyr7yLIaiYoUgZZM1yfGdrn
62/S89gSRvXzMNVbncWm7KrRqpN/cyX0pKmCONgsjyEzgWfEegXCNnNB315gfXnlmMz9UZhKb55F
o0SvTp1R11aFifR+573l/pwIBnVIGKWf0B7qEHr+YMmdE2dgQ8Hw9ey5LwpFo6HLUHU2nFv5ef/7
a+5vJdJFub+TN0PoH5E6CGb8e1Q2bHhk+o96h3wLq4GdL6ZbvZHlwCseq6TasAKUUP9zgPDFKJg7
kLpajxW/v05W3kii91Df4OjmZvSyCFkOL9e6sO09ufVLbe8t+9RqtpfCMRV8soKxS3gF4wOVKkoL
tpH2oXEHxixKwD1joCyGW9QpBqOaE0o10xrqICWK9rwYXhG6y9IEPEwe1RgDdpXtD5IcnTXQDzaa
L76TqiylBzcIIzLdKRgblLZLxmn+CC+8LzK1TuMjUywFQafF/RY6b82Vltqcx72AYkNUx3IFrjB1
sVdTXBf9QUOnNSgdxKwjTxrdsbT1bali3RHUI5Van8OKAOf60vXk0NYfCy8iAMBF8Bmjt5K4qkbc
hZQkFhhxMt6T3nzk+dixkSjkgKYf/FumrTd/F20gvpsLzMiW9ACnmzb+yquyRTxtQrzvExEpsyNf
wMqu+a3fMzO0HOYdztJCpAIS8SjkGMxqpnYhbMMcEymZwED9Mo7tNkCujimx42Lc/P3m/DnG00bQ
A48hxvHO+pYoq4TNOqQicorD2m75jiQW9XRmFGEA3q7OKZb/9cMUIlkYJO/3z5Z0xFuSSj/bSZnX
Hy1q6/r9GUpT+2b3yHxQc4DVHOHUdsyfekI5KoI4RynTRM4s1xLKD8yUF8+iC50gHsuRR/OdHlOD
78ouTstcOFXtbFJ/lfKZVg5yWzxvPcYOq5frOeeK44t9NK1yACp7erzC+J2rCdgToJoBhTbg+S32
tjrGDovB5l/U4vb7EJ1CGN9ZPXQG9acSf/zEUrnJ6sXJONNChD9voAzMyR3l5gamWoFtVYZZ4Pa+
WJNpCkZg1mpfHqLGd7i2IDbITC2tjjO1TX8ntAGJTJDaaNtLV18v0iIAwb297l6wXK9dVi0IM290
WdKn3dC8bVjcNkjB/BNUXh5YgIC8bo/5KrLCqEwTpmlacWqHTFobeZF/Fp91UitmqljH3usO9+Zt
kguE3n8SbG8g/a/5wDPEyfN9sAq6/zvQLEMtEQ807I9EyYpD8GhLlPL1crhVaG9y876SJsTp9zm7
oPviv3NemsUIbZtyYGNC+WYKmYkIviiG/2Ru7kh1Oyk6mw/XmTstwYj3oMSz/HdjQ63GPgNmSnGG
d28NraNtC2hdkfUScp80MJDtFYVnkOuDI2ZGTxRH5TKDSJSpYQihKEQ1FZan+hZ6pV/cCJgnfYPo
2+8IJZCQItLx2WLU4xR3qmsHpBBr329LQkl/7OK8Nqg/TxaszPfRpAC3zJrUSdsJh60zi8UgCzgt
hMLKV6jUKDwm+16GwhN/69bCcCDvghLw/f+iVRITzNdh7Au3PaRt341gJEqCuq1bPfi7i6dyW7Y7
tnp+cv4UTOL8VI6iHHZtRr5N4X0sZ/ASEQWb2wa3wAMXxtMu8M7CQChLNa1jETah/O5OqZJBSIvL
MqqsEmHnrS12ZVmyQ7E0eLpKHUssUYUvrBhRJSi9229d8rnmwKfxr18JYTDOVynAeznQmTkNwGtc
PgtivKSzS1VHhKQBw6Sy96AEYjf7GWy/3wndW4xOf2y9roz+qBTpC+zmnzoix6zfgTb6VMYjR/DS
tZDLZp4J9M3mH5nnPVgEJDLNLLXzpeaCprrt5Al0OUfnNINwdbS0CTQNArX7gyJMDSoq54rIJuKK
2rt0OPS55xYLrz9jTFtuDJ+9DHHDhc7q7et5fw/yN2VSzC18yPC4/cG5JWkrN4wYXVQAo7GasoLa
EXuQqwtesidOGv+rU249KB6nljRwLSjtBHWa+1uO3XXa6BXzWzg/yRKDP0e9+fqe3EpJKyqi/SAK
yTlUbGP9gKInjPy7UKi1IHEUynsHQ1q3cexrEQtdhKyZ+8kSPGdDX+yxuEMRhM9Jbmd4yqfeuTbm
FReR/NYgChsINGd90exoIUmVmAuI/1XwKCw3cUTJjyEPKu59iFkhyw2k5YQF5oD5k7uJhWWGC70I
aqa3gHmp5UrwX/7XxuTZ5XxXoURGntX5KaOXorm28OXEhgOfc6PQe/ncvmxih91QIoM1sJoennus
sX1HjOuNaQNsELzmGfOZUcWy/rXVefPBeBKTozRaJ1GUrbQdExPk6KrLXmZo4Mr4XPbhx4WIzHXi
sq43JLp14OXihuFqcacydOf4Ozf3Edr1fzGtoGQJsbLlgcagrzTExFUVz+ga4ftEH/3vEgBgC4bG
Y0r9IBPXJPKbgqyogFxg2EgBXWbUHBL1YwTnjtz5SJCPOgowiGSgbPmJt2FYtbhdfzW2tBJ6jplw
KgbIB61eFE8/blDcu90K0Etksu6iIZyKVenimAFsUukGvYcm7mNBQWmVsw1sgwo3VPsAaPyeX1ss
g0njcPh6BDCHDhHJR2Bfgp3kTdBiU5zXtl6i5qp5lFjyxH/0VBtHuppWvXnhPsnWza9IFrJW3u7o
OS4QoUyIaF4SZgF2t2cot9a1AikGs7YpTQsInp9jO8rwXgwyc8TWFd7JftRPwRZYTOZrs0upywdT
S5nG5O9/5KDere6jZgZKgZMUMATqd+oc/5+AWlrYNYohizVK86JbkIULq6HxEkq4qwrFJXULK5+t
m05gJtT+TTG6rNDMZuwhGdux6QPTpK9M/+lZiy8IztGdbkHGOCTNMH5zzKHBv19fGjhB4IXSfbqG
KdxFc10W0FvuxXBc5I//nVKlSumwYEInZftVSaJ7Yw2SQ4/ebigHP5D5vEDZasF+DE23pAHlpDpN
2TdeXzSvO0Pa5MJQXP+ihYTKh4IXEtMiXckexzCtN/vL5B1dVTDjtYlk9l605badf6O5PUzi7wyZ
SyTxU6yWvbwFDGGu/d6dm46TO5m4LAuqv/1xurFJzVNpA+pJ06bOqr9Uo1JFU1BKhCK7iFjYehMF
RqJZtyYSPMU8+iIkrllBSwIm9p/9KmFpxpyMjo+V+czSxH/7xoCL3PhOOyaCp2NeN/8VH/aQXf9m
xKG4Z2UiTd/7F7rfGAObx9GAhtrZesafRcj25zMD14NXL+YA8nRT9KyQ1DuSrskuM6WRrdcqFHkP
dio0g3fDuQBB6fdHYrD/j98iz8oWs/8u+Ajz/WJysKWhWSRcYEnK+t1GZZk4wFgfGYJYn3Y/uPKw
QUryo+SlXoTFf/bBA5fZPBYHJYoAKWPeSSPftwRzYGWWi2ztfb2TRY6ohWhVJe7GGZSgDWwNmQ0I
t+dD6bULTLxU9Ozdb5nac5opP0NEC5Yn6Y0XbmfXkU4KCUMS54goSyjDrrkxvFG6l6OKpF3opEfU
Xab7JAA5bKm4rW79KP26/H2efwNtE3wTsza2ROYI2+of6lTfy5EwkhYdqlFFSXX7M0u5MAo5ls3F
3LCK8mHCu4xEt46MhDJAuBtbaceir3Ml6FmGp02ntdSQJb1Hm71X1bVyhY1XZ9j553PsmeRnytq3
tcf/Nm/FGuc5JrUOueM15Mdy9A1c3tiXwx2MlgL0YS6el+L+u+AYq/F/DDXTbswRqzM/LCm5nWZt
zhtnwb8brNmhDTTSUcsiRMpUQEoqA6oTQUZodvyLjxu3sANdVp/S0Nf3ThlS4cujGeq65lJp8JEB
UFn0TgRO0zQxWIBbxDlBB1giHgSjykL1WKG31h4VeyNeVK4AotRyYbIGbGJNMR5AwC4lsD+N+DWq
66lnE3aozdhDKYwhSroB1RLIHBRucr2ghBcTM1p2OsfQb3o4pO7FkIMoYX1uayxmmXieMhbiKVag
jmXq54UnQk1aNzsL6f91j4oDBaXilIvIaBqkcH7nSPBl3fu4MAAWklQQ5v2wZIUiftyiTcuUAqTV
I7KRCUwBTuK2jXLS9rw4fx654A4U8oIqA14esIwmsvJQ/uozy9EqUZ17y/SPtiaN85yDQ+Go4PJ/
f/3WJ1J7XdNbU5roUqqGCTrWohCMx3aF7gUosC0vJlodaUoM/Lw3w9YVuiP/dR57fw6a7WzQeELW
a3SKsU31DHRohWB9MOrwNnroZ3JvHrmWXBj7MA7TxbaRCVxcn8EnKY4rSuHFchsON7+YZgqxpyL0
izCoVhmYZ2wwZckrqvJ6Em4KsJYwoTjP9gPOtdAk08gj43WKKGJr9mdKTVp7FEXwPpxmSXuPW4P+
n4S+by41DI9yNCMOet3d1+0bKBGAuZnFfwX9pN4ZIj8Y1Y6Yr0gLGK8S/a2sh5e4d/ePo6ngqNLq
fGGqBg702AIgzbCrluQRfHi/T8VHJp2xbKOZR92LVXQAjBOgeq33Rs2HnhC/CtUQ6Sbt8heqAuVS
sx6XW0VPFvX/6NYL+7Emj+rleX6V1wu2/bbL9fRrdNbQxfnmNx5RaCakWcDWVV7Q6FjrLOJTe9OK
/uk07VKjDEDhjdNWCyG7xOtYAbx+iy/p6/GwBT0Q2m8lqF2fXmzP10SL5jNCds+Q56cAfvgcmNLE
ugRLoX665bUA5fLTSbfaU0t8fVzmbIVza8YodvHf0MwigxMCF2uv1hhO2eJ0w2eoV9VD2JVkVTif
tAicUWTyxvbf+4nM05sQsywl/l6OAd3uL7SARNFRPp06lsLEMDgVrbA5pIrOEd3x1QCEm+l7C+mC
/UlExxMW4P150lC0f9Duw5MVrr1Sp8f/jaj1x9drpwvAs3n15c+/rV+N8AsiaylEpZXTsjJvrFu4
DOjsuqFB+cQeqjGk86sKVkux3DSzyOql68N87XxFosBx+y3XRh17cIYeOCDlD22WwCliZlp6aT+Y
f9szSdgxhbqJRprJQ6qN9MCyHl/orsacMvLnhWZ3L39Rr9mNt/i8OUqt87bau2rCadHWJTgFs1+F
kS/ExRWBUXsTaKK7gWv8cS94mCo0MUYLYd3Ysb4jhCEChdJZBn8ni4Oas2kroyoHikZ8kiUFu166
lF4FqK7vPBkmD2toiAdPG79+J/8ezVmJjcbfdQlkK1duxJ6/9u2t24lIPODfygLeUsUDYaHQ1rE7
vRucOIB4Xoc6lf1WrxFIYtuCXCjHdm7/p3rq5oy2SMm2DxvzuEx+SgzUO0M2RGPXk/DjpsFyLnqT
xqU9rDJEoTC0WV7ZV2PSGQETtIj+c6O8zG2mWizES1h9qY37wMxtDFMA4yLL1iqQ/RbyqZq3F19+
BSCf2SwKe4NijI930TXjZH7WFVRU34vAdGBRVZQz4PKlUcCRSJeeJKdYCtmQELftKFIXeKadYVdh
E2Jqd4010ivbqRS7f5Oh1qQmDnH39s8dujsN6066K3h+mvMIaaqX1GmugYVC5yCIu1i7iACQlu53
BCbUkKyQ6AhyqvkSkgn/DvRm4GrTSW8s5iM0pUmB9wjxexr8iz+bGcrIdMxp1s+hqxvHfRvCmBpz
nVxQ32VZW9JYu0M7qAo9EkzEhVGwl+GkdFVYMLZVYwF3sFAKk790fnURw+DGiUUAysw8pTX1t9M6
T1mc04AEAEfYn0J0s9kP6qS+rO4X4RB61n8QkBfbL3Sc9/gO5R+76nxuDiIwaqiE8p9nUHgeC1EQ
Sh7daW6xILMzjXDT1dsrKEk8wId51bU/AmOn5nNpzp08exkTs+dHaZOKapbftSak5j2AkPmOxZ7+
yyLwFJbIiQ1N7NnRsNBVOKMUqEDGMUSDz72vf30P7c5YVQYJvUWkZmhFRx81nni22AoTziuIY/F+
AweK/NZNRGovCfssvdpMyN7uvmoUcnd7ug2vX6Rg9GWBkEqZYxBvr+h5mX1VO4FautBmXL8ljVLc
3K53zur3HB0REfzocVveIyRIFiQx19f03GyDXLaR1BXTe7z6mD2b03UR1MGoI1fEWUlNTUk6+wqA
KkFRGfSNSIEa/p5juszfDWko7kEvl7DK15CIpB/hDKMK5Jgmqvv9PviTB+KsaPLzTTo+veKWUDz/
exEBkTwGf53cXGHUpGb1AHj8NaeS2pJhOxP1mSA/ABcNhl9NpnQXe67pQbZwYGWgBJPEx5Rcpbse
+6voT+/moJpwAyU0PZNJXr1ACkQO2CFVWnEA0w1g1gzcO8LOKKTFgqu3B7PyCQC195Yxs08bTHcI
14IWwvKQx1NIFZpFyH2tUW1Og02QE0b7B6iZeR/PxQ/AQ4yhBmfsAvvIK7IOyzytqBgrzIzHUM8E
1wb5rIhjRMtRe0pL2n3Id5Iy3Kn72qb27rytuggY/R4k0Jo/4oIYUy26g8UfxPkA277ZzFaTTZwC
G4DDbN5SkSFrGV/viviLdecuBY66aOjU67OtBPy0EOEU0MRlJzLiLIjdTQ4b+wdhTNfx/SAYZqyZ
4xbdYgaTy5q8MQCvbW5vsR6dpNteWr+zJ7FLqtPCdUSs9swKI9X5d6mnopjWcJO1U08k0rZPodQm
f4dYD1vBC3J0+pc9K6NJBga6KG6YpkeodR5JtlH8gZ3UMHAy7mKhEOkwDKYio2dEP8MDshZ6PfKo
k5OxIrjcmjtdy6kmF9RCG2aDIBrJTpwzuTBfHlaSteWMJjmKxF8Ui9wXHmrq1OU6eYpl9+YMzt80
RG4Gmhz8rbSfA8oXp7YpZ4LGHblk2RN7ryQNEf8uSi9OQFJou+16ShFlanA6fxT/NGr887LfJZku
3U0a8P3ZRLvbi2wg++uklkF/TlpqYryKCi9uaadrLrZXGgSeVX0suuAf544OHg0l9N5vbIMF/pzy
eD6gdamjVN6g0Mud/vgO46O8ws8Ku2xlcFxd0pXxe9y+/13ZQ67SraVfIOgz02hM86uOdUMhoDCk
57z7oBuVy3Qvp6DhXbImb43Akw4IepewbwdmYVsQqeAuKoGJSddDJYNzbYzpDD1Vpl7hj0BWw6M8
dTO/rTtnl9HgWcx2ucppufHKGXl/VKp6qwn95F/CDgZUNp+tvETQgGo1W/9FM0dQn4x1fSJ5jZ1T
D5rVGZ46+P4O0LSipNx+GcIg7nO40X4io/NojIdFlEdVOwiVC1v49HYqVTr+IKkd5Yk7tK19o4ud
A1SuRhyxWr/aZn9Dt9hgVsoC4TIIn41GMe6+A7iuPlA03YA8nmINOcCyovj/2xAxl6UW5KLxij5w
6z+anyZNPa9hZpTEowbx/225B6H7MiSiFxFNIomP75i+/VXa0CI30EYWxK9yGa2LmprSvo8884mo
1axMCQ8Mew83M5G9P+FTFZEjPSYqpRPgihO7c9xg0/iwYifeLyhmFcZMKSREbXlKnYPnN8/xjq2H
ZA1yI1lch9keKpYlhqNCTj2m9e83l6pioYUfCuY6yESpKLnquc8QpawPUaP468fdCfsnstnTe3bD
QOtn72m4rAUIx+AWX3RFyPt6Th5jV7i5nuTgenr/dpItab+I+oE2lYV3Lvs1cBeC710kV1LOshCt
tyyKc9CMXJudaNMYvOi6m30ciWWvILiqYx5oZjQykBw72ojfcfJv+B+arWawXj8H2TWWodOUKSc/
ZnO9kboDtuZMUgYOkBRs4+0knmYL9vQEpdupSDeEdSiaIvGymEbtTg4w+8QFAKRDdGYLbykLKWwf
6UwkHjZwxou9GxbEYD7NvH6Pfh2wg5DXaOD6t9ph2u7wMRUR7HWq/klpt30aXOozCwTRm7vTaOyg
4nrQOqupYOGTqGeeSjavlISNYhdrapRDbUq8IpO411PFepg8Px9jrw9jrAqClY/UjgP7WfXZQScT
Tr5ChXml5h6MPXzwPjt7eQKibKPMU3HTNgOEpPRxJUadkn7wsa8wTxieqGFE2l+G+BL2iCZ0jS6o
Xwi7FCfFZ226WyKwvry3RTfs3wyIUZVuuvljYA7nPZTeTMmhEki+lFOE+WXh7SEsHGvl9mvSoKmE
appp52OlOIM7CO/RlaTQCf6XN681SRUyNa4ZYeoRlSdz2L+cEntZK4QehsHiBqDFqmzijM1gQwg6
1pF6kHR4nEu27Ddk8rrvfPrevealCVQKxgJXxl0T3vXqQWfgLme6c2gBToWvSiUONzFFQxRzAAWl
NZ5jqiu0uO3vjajFjuJ/67XbEs68FwLHrTWt27DIfpI5LzKsRIiTSrIf/t/PqnKAYqkhMjGfT+Uy
ZsaTXudm81PdYixoeQbbLI00Qo2Gb66udoWrhUyyhzgI/1Baq42InnKPmf8Btm6VgUgSllRhilc4
R9WzfWK+Ko0HaUxIrzwlohhISojQ1UmzLI4D0+KbLyHNXR+Gdskyir6J+FCYqjU8eYuIm3sOWNM0
dHvSh+LNjp11DaUOdfCFEmzbQX8DIxh19sM103Vj+8g9KQUnfnTQ2bZHCs5/1/EN/9HhHuthrZNc
sl7udvxVvjpeMd03Cpn+z0C1cG7pT/YpXZknd3valqH4EwPhPrcdZo8VgmpOtC/w4ISKCB+CeGOh
1hnbGRjkMKTdP1he07sSNvG5gIpjrq+rGURRIAU8RfU0i1IBxzR1bqR4/3P2rJUvebkFy7rUhJZm
jl8f1zIIwkBmab96E61Mmu49M5SYKD3lEa8AnWJ5qrqpZ6ETmUZb6YuUee/w3pZPyYLFekrXq1za
DyUXuVGVIy4DfIAV9O76aASh1SB+hjbEE6HLePU1V6g0w+Mblw435tlMJBKKdr8zWX+tc0ffxgz5
bUOaY/E7g0TLQckAY+Ia0/IiVHdum/Q6TlLZWoZJh2X5Z4MZsrY1u018DYd7y+7FqUkA6h1gTVsS
/5qzZ8vCBbClreGLkyvbqjAeRkhys7iA9yOt5PsSNG5i9BRLYXMY82GuahGKvtGHqvzPrFG5fPvF
70picrpX5QonUFU5mut8kt6DvDwUkkL2uankLEdnPuIJwbhcMq7o5UhyyyO8Wxxzb8W22fXK2sCn
78gVMqfpQloeKtK+7DmreZ9xXY+kQ45SDhkNvvGUl2XhH9Nqx4ogFYyWCtXWrkKaHnWvnoEdrSCB
sNDXuEV2Bn69W6V0NtrmEmtPtMRmK4DU2NnUwLmka/kU9ADDoVZnZqKHbOeUTNRfRVxF2X/ckvUb
8vHF0TxoOZ6mI3zDMbicFgokUSUKfYf1b64A9sIzeEggGUaaw7pDb1HV+tXEJFl17dYJsZEGLwB4
R2cS24HwtMB7hURO2u7KWK7rG6h1BLNqlu70W2DX6Ask6OeHTUkGlKHXGiNoKezayVp/cTmTc2AV
2+cmTCizEgnUJxA0JjnAQ5suMqp0QS7TD80MuXg87N8zxJbJjJv7cs8TBPWi9GeAuqqC57zMsAdX
niLvN0niGa8BsHkoH+tcbrQ8Jg36TgQpl+n39w1V3ndCsmAuyBcsPYW+7emoXdny+Ua6SCZq2cRE
UFwIWTYE2h17uwjlJ27I7Iys8dkRGemhIqaTt0EBXNnaxaQf6wXMkIYBH3CaQXlMSuVAP0UI1V62
EUanH8mwv0EGP09oJx/zic/Hkk3H0UbqLx2Z09ZD2gCXmvMCfpanQacWKCUV7pYndETcspWBbVTQ
zW8dL4iNI3+FS2KweqsjWipiUxJJxj0+IDHKlAo78yZ+KQ4m02SRoT5JNMMj9A2zHbZd8YT2Lt3x
By5xM1zjVS32tEjhYGuL9yO+yQxMc067ikPfbFfQCZURjY3Ymorr91QxziKd1opQreRlYTuRdbHr
RWNSDqMhWt7UV6pPhZUAp6emXNxWCtwIFPR8yiSYa0eS+XfuURb/ndmjqBTtg9X6mClX880HGLPv
0QjBBP+zU3NfskYv1X/NP70YTOO9g5f5o+Y9QrwRDSLwW8uhd3tBlIt3QoI97IHScZWYbcBE5/Ci
HIPUANFVirDV3rO6Pi1DTZolgan7vJznKvjWuoXCPNGmsZ9JuJLL9YccUiPqvG/MUN9aMcoPpw30
0Yow76K0vaLFOMMEGpFoECpgxSlBooRebciGUHbJ0poXZ6XugXsj73gK+sGvmquOKGjP5CmrwnDT
QhDxh0xKmCqEJpwaEs5+9Ab/i0B9Hz/y4HGB2TISqnbzgHWruOd97V4oRKloPPojHZGAeHur979j
TZTQ2BmAbb7Nt5rn1CVjnxt+9RXKCZi97Q7EJ8RvWXvWZB9b+vLeROX8+YAQQamIyMRUtmy7wPB4
Bh1z36XKOifoj/bfHA3tsZOFOnndzUOi3KCIX/4B/POgjR0AWe87w7k8sFKzLW+kxO3A9Mr+UxNn
j0SJVY4XU7eVCujYMaEp5ozLm1oeQrsvwZIjkAwtGK/Yrvj9HgnuvlzrlD11hm8HswxjN9TH/xw/
HWATL6TExtdqWRWy4s2M33yH/M30ftLiSquom3meQHk/8sBuFwi51kDSjHzy3vdM3KuHaZoYakKS
6FGJJyBWj4PRwj37tAq/hj6WLFijF1tob6hx7p8frLuKhQX/FCwaqC7JUKcImEjp0FZ9SFQhV63C
SPS3SCKkx03P4BUdJR+tMwK1qd3xJ+n+eu67GLP35OcpMSQeldbxhs6MPtRL1WZXQilcHcUaVtmR
Cm25TLvRh1OvNay5QR6ycnleLFc9+XBlMmenjMzR6rkpnKkfCrLaq5szKbS/XC9FUYIgc1Hu97/R
400N7GYxjYOgqjbx80b8KOoF1y6iG0/347tex1V2u3eh6PqHCnNzhj38sN6VeqfgV9S81oMRy+BH
B3coDLKyZMJg9ouuRzEk4lMT1sBJKXCsFe6gc92lnqqvZudjUIKSdZvyCooaWfWBOayGPYAf3ga7
3RySuE4rNvTIL6vkwRi9O01PAf+Tirc+Jl/iw+qE3NeC0hc8HuAXCHiDj4ymN2tat3XMeULenV4f
q+srytdEt+IX7iaPoa7saY9IYezm/40peOVzAT3PkFZc24waLZIKRnDkTmFtHnsDyMm+hXuldNgq
VUwK3jC/ezwBxBfy6NhebhYQNOHmVnpDX5q+STXo2/dnWbdwwb40aSNlL4yLunB5y8FS5cAndkoC
9uJdx3zF7WehMY8ZUfBDuozE7d/rdyZRv4EpyUMa6NP3q6FzxNPBJIAYZmdBB85s/P6m2xm7Xehb
3Nx1J/rmyMq2t8uU35JAq5xvLWlievqUciXFrJe/U8brJ4JubcMDg0tsb/1P81t5N8zM3rluiqrl
SmPQ7DdKOPbYiqaZuLE9AdGvO0T+OGSqFZsIDcKDmlhsoFZq6boe6YToWNyHV2V3xm4eQ0bqTJih
/vqf34XZrmtGHBpfrEHNww3ltGcpLrdSOiSU2Arjwy35i+hqrfTv4ObN+eHZhi7SpBadRhVeG6VO
uIdV1ytr5TgtoRzwPGv4tbuVKG40FdWGQM+G6k4kRi2Zpcy0tzZoyjr6LStFvGuIVs0mXkmmk3Yg
UNIoI2VvrzgPhtg6OS1qFvpxnUNP5S8+hVjzFWIYTe7WHpRa9c86cV97sFyXw86jDEsHQRHCv+sk
wMOMPEj5I1H6Kv3HLC80LpY128UvLcXzD3stbV/Fv1n3wGEsDKwb30TlOZfqb3H7wDO124fPl/0Y
6xZjXkoXMqrzQPapuad1fWjTJREd2KYNsSjECWSxHAgJnnzTCd/YOkmUOyjONH3EVY1jQTEy9PBY
E8mhSp5dTj7iNP9tWOx81K5lz99FToswGJgCfirQoRh0LIn1ZIsE7RS6aVZfQEEzjSUhGWZTSxXa
R7DMecDmHok3xXXIkTyA/499vrPDawAVh3KNfum6DCh6FeSDnqAFxoVkri3YC8d9JhLtKgnliHfL
m/iSqpP408maqQ9vyrzKmhaokbMb05uskpiNnRvXsVswjYkOtFEOrhZWLysFixw4VL7U8Q2+w4Vz
Fzmw21FwJD6EppfUcsp9y3XdW9WiHvhwW+JKz3vXn62+8CBp7R/NxeD7tDrjsgfY/io2RcGZpODh
GIVuRzoEc5ybbN9k8rcfvj68gSJeiln3sduxk+GhZ3ZvQGvdOT4U61p6JNTv0b4hE41y1SLLzZnD
sunoA/V+tqPSh0mK4sSpIVC55jJWmiYzArknrK6J/eKk3Pw8qcasV1EP8eJO0tvaOH+rU85rqW4l
uskIArJiZ1Lq+MqrsulB/tkgeQIAI+d3dwzHzkI+yu4CsOegC6N/xzaadQIJX6U/n7KdN79KBk7c
934oFLrMyFLvsVt0dDaV4yp6S5g6qLmLuL27Eey0DCaI6fTItJgmZdYl0cJXMgpSAeA25vkN74Ij
i6zt3zXM+py0vCp3n9UGpi1ojR7jHmoc/HIC9iZ12ESlOA6NKLS83XxZtWeGT/FwH6oYBi7MySzh
Rf8qXBqYLSqGowm+9PCB4Sf+8cd9XXNkesUKUvRNS+ATqSL+okaXLe+pukx8/mTSNETEw04VROBF
kotjStUkUtinbcsSCyZNSo5yvjnXvXCPPmgYdftRlcZz/mOggbePTWMFYQjX5mRjkabguM30mFab
6Gv/8BrITRMMiSvDkYyd216Alva0fL294nOfr4Eq7vHvBDuTWJlAVm0QtKThWc2RXRbCCh6Nv9c8
ijBV0i5QZU4moxCEhXAt8A/LQRwUKbu5841hde1S/dGexeL3yRvkd9PtxAnG7Ei5rIYQ3oCR/EH5
2Qj7GrE5w9HzXSJpdqKP/P26PRodP75ro0ENGEdypEs4u6gvyN/DRJtr8tLzMLGmI4HgozgzHpxp
XQfaWcTBUGnfjCbOuAchOeq89JgyM6FIN8+wXdu6DLz9uaoFoUHBufnNjc3VpM9lhWAXLV8tUy2J
IeszvBEXwINGAo+cAnOwKnZJZ6cK4EpTxAgbBh1Rkr7hk6U53Bh5ZDmth5cKr5zBTFwOjsJYBocK
dn8p0qBp+2UwijdM9ILSr2FA41SjZYF+La8N2lfkP8qLT2WKzJF86taEL5RXqqjZl9xDNSFVHZtp
I83mAJMyNFbwl1k7PSNhUdBNtiypFXqPwgUk9jEnk6U+2SKz8mcBV5L7FIm2KGl2o38BoBXWPvFX
d/TFatobTc3v5CbBZW5XmsxGsr0Bi2XO8rI4bQlYfFWix5SWjV87Xx2FRW+yLm5U3jwD0W24epCm
CSJqPmATjB1k57sU7v4aalUXbcWUcb8yHEBbuMq3GfaMY5ceQsiSXXMFFxQ+FD0u8NccuWJ24Lcw
9RXWt2Kan9GBpaGbq3FtHys7mPnCUtjMEq4HG0HK4aq0nDy7Tb97MDWqy+Ty1Xc5pymY872k6u0L
HWC4kU9Dxq7uzmiszkM8/yp3datA/RDjItzTLf7suyiX0hiAqw5/fzxWsezcmUsYsV86dVsbidTl
lOyYZa7tp9hg74AsbLrQTjHvjrl7EYmhWxyDu5aiR4TNX5bbO7FfHWmfe5U0JpgEyOfBtP+XtEFL
/zXy89oPkm/21WENbj2zfTv3BPJbJCKKeUttqnVIt6FHB5zsqCjVoIZTmqrYN6lypqS3zPg2dkbR
VR4R3/08fuV/0RD6/MdVyNci8dSHljgZL7c94m9fDIOiLwH3A1IuPdxiPb41aBGvvfi+/G7Hyyuj
2dPyznTk7by4sR14SZZYvodKndU/FDBoVVn7jTmLnKTQFkJbQjOBUXBfrufX8ZpGN1uxtOJQi5UZ
/3DllnnmjznAqc0bZoRFCLDevMP+Kd68KKQbJVu0oWXPSxC3Hsj3RyBTxUeS/lPYDzuIHmLHitwf
YW7V21VqtjJewI3R1+Ja9AlCBg1td1T8N2/Y5ZmsF3VMZC9p69PYu4eYnhOlxlq1FtLFN05rijbt
8xbBofFwc751lkQzJPSI1gIvHRRBhiRF0Bf2C0zoySUGzRaJ9nuGj4gma8qyox61eKT7vzHsnWdI
yElN4tYdtm2QMD6YArS3X7ROet1b7aHWlxZ6rmmpxsXCMhoN7L5UC5LIhqs/VQhWWEbyoWyjRnDk
O19M/lg+9J7m/6fg5HtXZ6FeRAuOm1derpf8aJDpfTDMf8A8Wpotn2JwZM3/IGIEZbQM5V7uJ+0P
ViS1jW56SfR3QpJFnwDG17/8XaoFUQZSATJmABwsEezV1jLiEHyPQvb0eyrOib7kf8J78cFLL7Xs
kZl8aBAFI2qV/pC1nTAT3IspHWVk72i/LBSyNzziOJ+q8roMqc+UHkBvRuprDbw2pHF9cAb/O+Ap
k/Kr77nx9c+P/DpGeYnxIjMCFU/WEBb1C42zmZ/3AuRbwXga77y9zC4iqKTTovGNdbQ+L06VOpLS
8KhpyifNeLMRU5P4aaYSXRld+AMylvZvIckHoHTSSfnrUmzYGQgq8nUrCg2NN1qC98I8PIx1TSgq
mRgYD4YNJPLfvtZIb7sM+Wh052XvgstM13AeTSOxRIoLmM2RKwNX2r7IdppYvlwr9+kuE+pQNeAE
DBK3AqN87a7AR03WRdbApvfzcgCLjWmNqphS3mxJF7EfqCU68T4eHLzSkX1jPXlIAIKaPQWbPjsI
S78Gv113/h9RHYrNUfEHE+pdrKcea7VdIyXDbLII2pWewLEg/dB/UoEzgWIB5XrUwpfUJIbyWXFW
/U/Yqzu8WUCUyeb8bVSTtgGL+T58KGwJ3F5GzJOl8uedZKfirvHZIhHgMTwz6wxIFf2MpYEYZ5uu
Jkwj2/jpsLEym9wAQ3OCeTa0xdBQzvnB7RRpYe0WXinq+mcAN8OqS56LZQvF59W/lyVQY+HrrebE
TFJFspJZ8FfG87ZhMOsz5Zz875R/DkXMeOsv2oDGaWzTLi+IfAZePhgqoO/vbKAYYOM8GWGKrpeP
kzhp0CPzznVCq05fNH81NQEJ4szuivr2HUvYW4ffG8mKHnbQVoyuQzpXTpIV39mCvfIoccchnQ9R
V4zjkClqgj50m6U1GnK9XfLn5zKnGU0lJPe3Z25OQioR0A3RKqafJo6aG8DxsthS3FG+gZVUwLGl
aluvrwV24e/rSivxG3yDgh4JC4X+ZeynlVQ1v71FV0MWIHQbdsRq7rWDGe29pA2MKKNLf8c1HB8v
aBvNy3uTZgStvfvlG31WwvN9TGlP3zjC+j60pgtNLg7uFH82mxgBOZgP2kH/uOs/NJlaKUmw1MyC
zAKgFZQ9dLGI0wLPQRN7cn3LIqcxeol6MAowZ5w5YXdii2PCCFWkskG+sZScWtU2CNXnhi5ghoyW
FfA8Tm7aOI/e8bPjHSwcGmSNfER7/i+jWghoQRvS7suzC5ny3U4pQrKpkc3Lxp2R8GShb9q52hKJ
aSp0RpQe3bbSMLJM40Y0itES0wcFhyt+91o/6ZHzqE8OL57iAtzqf1Xlx+isSTQxxMDQzI2iBdO0
AkCHCo5gVbX7hXuBpWvXT00ycS4eaczrnIkIMln41Uf8nUEF+E9BCrrL1nMCS11C6D4dOQe/+BQT
JymnCrV874HG3rAbovKeYSSqLrNUpDgjrvmvL2uxbVsHKOQjQD/iw04JxlirPGaAn3FVqp/Vazzh
LqprZfaTnZ0lNThyW17lDLGd6qbQuuyW6xjLKyFPke6QgcZ6cQRR2/bZBV+n3P+f2UDhTAZTFVPt
fc9UtUMQ4SpEbQXpf+hiliys+fqzxt2gkr6GH/zBVXzat9YZ3StboEPwBTpotgCovcdgOQNukXkd
Gj844dN+3tp6IqMxs/Ux63oFOutPJ7sSDwGgCfk9AvIaWEAYj8uOSv1uk5owE5Grelqo5G3PMDJR
l2jXOIAkUcFFiv9pESuEDb2v41VctvIvkxmF675WbV+HrbXsCK8wieSiBjb4h+wHSx8Vw4oIEtdN
US2wPzQ7a018a+AMgXNATjrbJxRl0wmWWtcJmIrzZ6YX5nqAVGZNxS2xCqkqEuUew4vXYJWDe2i8
1QDH9WeSoSz3V/GrrDfSsJaaDwIKKrK6duqlP1Ks3Ztw0sR5PFtd+Nzx9RqtnEO6HdMg1XC3oygY
FBxSIwW98YLJ6ESlU6hC9zvJqNSqCb9otYYPImEA5yGX9/wYS/UGDmD1+pj0MxqD0slh1vVTwfN5
NYoj/Z9DbJ4W1ZZdM4NxrwmsSIXdM1P+x+gn6rebpDPPU0FQW0/2PaGodUAgxHwvGrz/1s4WP5su
dcRemg1p6H30mlvt8uacmsrS0QLD07RRAvtTmDmUusulb8a29BE8oFDnaFDoUUSxR97xr3G53BaR
WTnfBAH8aFTfJOn+NxOkPljdnpdhtS7BdTQhG7PN0OOWcNp0TWMTwjQA/7N8xHss2YTzCVGr/xd9
JfiIcR1zMcSI5c7QOYMdfKBewlJ4GVxjIK+Mu3zYuqjl8AHOij8o6yu04hiKocywuAcsPkrCNvU6
VnyZefUNKjZRCj8zWBhNxNQzQrIDnMx0RfD7CwJen3lcpix8gadZ8PH7bXYL7ASAMaJgAm6KpfDA
pwoelY3bUu2Bq6cT75avuTwKgzdcNQ6j9pqnTBT2GK03KeQncnq3dz4G9ARds74zsOOIYMy+SJeT
wHg4KK1mi5dFERqn79XQBryQ08znasshHEqnQJR+JMP9YVMmiv58mMptQh+gXps1UFl+kIU52NTh
0NQ56O9IOsKomLe+7NSTePxdFZMmYZ5uATdf7XD8ePYqHdSlMqwEEwRLMeiC6ZpEbKtQ8oyXX50l
f/XXo8xtACVqUBZtN2RvKA4t/leL7bcpSL2YxknJlDp9dATLoccgsds1UC8/9H3wL9vSQu0iAko9
l+ZfxdOID0c5mT861ClV0OaAyTMTqahOBwyj/yV9u0P/1X6D1PhJ6KfzIMkfVdDtCIK3r3HzOBzc
Cy0u6pMYLk1vv/NcrDkEl/sJZvvUsLGhzJpH+ngx/v4Q2a4zxpprCT+LGPVWI6FIGCxMm/SgsZCs
nNDQhj8UE9wWxV9m2NrO+vb5nNYWdT755aAyAVECDF7vX3jXdm/JZH7dcVc8PZxiI7n/d/OsgLEF
XeAkqrOK0K45T5gWsnqsiugIsn2oKBmGR0WTe4I0Su2Fh/vgwomuPjztH30GcBykXgpvBzBOg6Go
0bNSYpFJBnpPlvMubYI2rpJqBM+59ksvLjh59OmeFyKkLBDGTG9tHO3uwuJRaVqbluGXAEvmRUHH
AySomlFNTlTEYZunrlV5knuK6czLkJOD0VM+hzlnIJt5P1BnapiQCVPkKnZAJK2GLKx5LDhCR7oC
WeZkiQ45k+UWqJCrhmM3JQb9P5MoM4ojPXsQAqO86sUsaaZIhl3+GH0o7n0C18dQxFdigUOFqY/1
V6FIlyMy4b+ARDb6u/DNPg4EYz+wq6MhRWiRtw8cMY+/Ygp1PsMSvMNUooJgLR1Iy4qeZARpKWMI
GIVKfdW+UWvGuVmOdDwJP8oibAkW+7LW+FfYUQbkYj0RPZbdiGGjTa0F4aPZATBAwTjjL+ziyctJ
wAUJIo1QycY1aECuCvQretybTlqbA2aLLBamoHezwsP3COmH3XEe9RXJ+j4Ku545piey+h1vb+sI
saqaWxj6Fa+4mEZLBQSSzmZRgvmgM7Pa8B9hby4mlPRSInEuAeQ3UFfK/N8yjfZ4Gn1RMpTIBQRt
3s6UfRr61Cv6n7um7mR2d/nNIy+gbBk1Wv6I4H7rFLCEFQw23QbZ3/6O+btVV+mx1PoI9koE29qi
2FJXNkZA6ZcVMpHKVyfR4tw43700CRxQMcFlzNDb4CQwYmEbnOMceZ/n+nBbMNSzNmrYunbLSHV/
fzpkeuFg6RHU4+cbdX7e1j1xQTQYPwF3JKeYr11sl3Bb+defVPjx+0uUPOSpEzf5e9keOoTGV1aw
ZXu8LhVUVQ++MTy9HQFvKXYk3D3h2OSOuVmIsVzOMcHK9r5e7WV7R+y9z4zWEkO1L9DDOTrbHB0c
1U8hPrgLCqO9sGd5f+rpS5CvuHX6mjeEk3PYzoJGoG0HaYN7nZdNgbmuefw7UvsE/9p7occjrozg
HgNqRBsjrs+KyfOrM4BX0yX+8oTPfH4ehBMitWdC0VcQhScabHUb2bdqTIYVHWgEBARdChSxt3xA
zCuSYrrXcoAXnDidJ33+Zi1Mh6sC2TtDS9R+dfZAa465k9VNIXui8OEPpO8mTaDYt67xihZUJyNn
9HvU9rjqVXMOpVuF0pQNIsSzkdk0cjEP0siYKz1hPX424Vjrnqlti4DDROWH4Mepu+s+mL2FjX47
pVPZBNuJef3aOb/sD/kn4AgRGFtwib2GcLCceW61188xPlkeNPG/mzcU44pWIjbyilhzed5QB53k
INadi1mBKc4LyV2+clbjH/SAVCHhX0XBCffoSpPWt0Ow8YBQPLSPeBPqFt2P4f1IhIaMJwD1kKwO
wDt27vn01P50RbS21SV/pPywWCUt0OImju8NzrazzUXvABvn/+hDLmvB6CHWj5QGMF0mYbKLTd7A
KXKGUgvHOHF9ERYJ+YdPG+ZBDoR/pd+FHE8cN1xj3zoOFsVTNavSuaTCYa5xL0Xpbs5Po6iKv1CJ
eyYqKSQ5E5vqFjXRL3PDbtwq/W0QfVNf3up8kcC2O40v5BY5ivh18No9YBBeXTd8a8inyGV+iu5i
+5oyxac+MIXpwjpZJieAZfP0B831T483KfvdGDFAq8B0/+/39EMXIHy4UCPI5URcODgO0RvOr37j
0o5bRJs6XUu2q55tz3Xn3PeS9ILkLlCF8iTNSwd4EgqAy4Um5vYVndto/x8j3OR3PRJAiMZoDjYe
OQDBKqterc6XvRVC7ZfReLcTBLXFuUb5IbyP2ZD7eIQrKgU0vOeF+tkRF3aTp6Zjb5CPF/VUCfvZ
lJkgLaQDkRsY+fQAV0YsZWTTzfxqIsuRef9UeQO72RmDuhDTHaFuMAglKMkikIunXLmNnO//2vCg
ltCbbX9NWMs0o2K+vfW2D5SnTEfiCe8/bD4v8ZiYZrdhc55EfRVc6HR3wKByFUvDlE4lxh91AWLF
5saraERxbiHx/zVJVRV8sIsS7G3QdgvpkZJe+/0tlTUFLm0G9jT3JgydxCCrxbbbkbRNi3mvkUWt
RJrJBeoD/2LT9orn7BeVIALmk3Os90h+er6WlJIxMN/a9Da4IfJNWFB8F0vc/7SvyON3ckNdCwE4
Z6SpkX/RH6C30kX3CgUxDCfOQ8NvI/4C3i+KIKovn3bvyqpz8ktVzAvOMAofiH+TKTqSwcM6Z0Wg
mLW/C3ZKR5huhm+EsjnJNn+OK2+cmczGo+SQNMdTJfBZR/qC+PvBj/xAKZb5Gh5q2RcoorXR00hh
sJz9IwSW9wBpwg+K1P9zSBwr1xdtmq+2aaC3x+KFF2tiF7CAY0T0ysmDC65oVaQ81Hx0/8G7uDzC
1x20/9Q8Q8TVcZEftZ9jlT+nBu57hfFkMUFsxZYeqsfbQ1NDnzlc2iA70igkB/0mBvP85YQ3rAUN
2WbSBTy7/Xq73igndGVsf2wPiQEZHeM88V+ehllZG7kJr7yQyH+7APskmsLO/J9tKAo1hIsD5/Sw
dqVh4JM9CFy2pfvfpMxgBOou6ZNwggMgGG6T4XoBOPM0ZU0ys2Hu/GY581FYMthVMOXKvlhIhIsr
O4WVTy5O8HMus49NssgnX2dhs+VZ9DZ2IPB0ClyvnbR9VOzY4AuyTk4aBfaHQ1iYfkFpVkLmuAJW
Gl0xwZ3WA2VkRFqn/P6FzEe6td3oA9oQqaAFGKSi3aDnKGXuoMmyGCcGqCdqdyl7KoVkaKQ9T0S1
A3BQPqtp6J/JB/NwwW9wF6d0eJNAZLdOpjH90QdGLexGCkDst2P9Yp8JB9D5OY+vp9nUl/BnvXJK
G75Erfj6SRJzWK5I6QVlCBcwKqDGguT1cok+x+Xe1HH2V++TCSQb6Xo6LK72fNgHCRIkZZxfy9oS
mkzUVWQPclt5Hxq9jCSOlbEBcK3gzftZXew9f16/YYGGrfmZi+J+UqlU4NeFQu1W7E+SJyvniXlk
ARgVihk2nPrWwVQeb8ut8RV4iuy8XEb0ySrnYthrHROUg+nJQ5QfZ3mQCWVJC6rbSAKH1H4wfwTV
ntMvTFwbdxZbbfaiTCDCCku3FsXV6n8eerLimwZ3B0NHuP+4MNX+vhlh6P17Tghxg6cJhJpwSF86
Q9zSi9XRx7P9X0R7enhgQtnJbcD/GNFHejJ2CezJ8zcAg48rRSy6RBi8c8AOIZBU6doGd8nLnBs+
2/hZFsKeaJDVGyLYjp9pgLAOIDoMTZGiT3Zc1crIZ9YrHmuBPRKArqGllyzSGje4q2zUpftFyhGG
R/0DYSXiINnIbgzcI5luvOB48zZvY+UbbtJQe6pYbYBTD6UoS6Mv5kKTL7Z7Zgis1zFfNIUyVXqP
YNh9/GdqVmd4/TtJRMPw7PmqVxywgUFV/8eitSW2Y5gcVNDhes7kRZelrYGempm7bap9x0WfHz/z
7v+vQUELSsoH4vW1ToVI2xfZ/KM2ozjzU3D50JvDanc6LvILdcFj2ieBOI/G8gEyrX6TRgGxp7Gv
uJK15bqaOffd/Iz8QEtwPbB4UwEfY/cQFhfWfXFEEG1kd82oUWiTNMrLtwVVu/27tsWyxgVZX8uX
x3X1UN7+D1/sJgT662/Xvt2xIKttGvYRpV6PFNqAWTZpdBdXYbFesaEkSn5udLaJi9XM0nAk0FV9
tCl85jBpt74gby/LEFdulM1E3L1iw3cMJUvnGhWVO8IUmmn5e2WZ/SY+tL2PETWXKRt6HL1dTMU9
gUvrB8WSkG6wyJg3RAZLJA5rGHgxVDwlUOQtImWb4/SzRo5gAZ3iwV6GwOiGO7d8xvUpd4v65HZ4
6Eg+lAZUb5DFLWS1jdndnH5RZs60xGdaC9ZZZXoavrK2lXaVwToLEDLQvGVpTe+9lq8WjfTe4kPt
oLietOMgTG4R3BVU5QFC3ySb6awt4MgCPn2yQttf/YrAKtGmvAArTxr/kRSMsRa5l+g7wAZwp6OO
zL2Yh8v9vqTuYIj21ZX/Ic2481a4ibFE5wVGz+GK5PVThs+hlOurAxdh+WjYXj+vFUwJ/2pKgkY8
SC9wR0y+M/QZWvtUPlJDBi+69lzKwo3Kyb21YEAXUhLteka7yAQFKHZ/cSnXZafod5oFRfnZy8IU
iYJtPeloh0qfXhdOdg2aExz4I6yZmCM/7v89In6bcDwA/lbP1sz4zHzFYq5e39GM6jvqIUGc0sAI
xdFFVrsHAfUNMlU7nodLFQuO6zu/1y6RQprG9exUNrxCSFmpFVXo9D3tzaQQEcrAZYcAfqxjqCEH
FbWPCc39cEUtnqJ8+fE30zEPBYGrmydfIRm50UvFDAqm04sqfDA3h9FOwXRfIjIc05ynIV1o8fPY
SlOAzQGm5RFoiy5TXk1/zWBhIrsfNM6emKZFxru4bZdzsp2d+iQKH2dcYYkF05mhjoFbSTnRE49I
kW3rx9UgQCCQC/CvY2GAj9E/1aHUM863N77DGQgWsKeSmvdHo2+j13+yNKBjIwkesgk5q7c3ZqAf
exqYKapPgxkqcPfbOc5+fcLTyNLb4sPihjsSsKVGS1KIh1mj8LBhavIN+KsOVMgk29NarbZsbszV
fL7zSZgCVZARLlal9A571ZAGLSHkLvhZhJBxhZwacF/b02EyccEomoEzDSsm20AF0J/ymmpqhzXE
HYCiWozwaJ1mk3fe5N22oNqKXSaDoX7qJogJXwGV5/XWWsR39CkJysjUxieTwu4lBZvDn72KEElp
uvXLyTE+Tu6YVoIYdipex8I6nrj12FMpVLfu2pDZEVFCP/cY7SoFZjkoWEZBbpDucmsmIb7NZQMx
HGUB5EqDCjOmjTUUEIgdF/XbVOBd6M4wJYp/ak0XPyOXX33mGshpZvQL3C9eKvgoXpIuv+OMa6k1
GfKPlcqLwVTRYvOvjfElobzD/vRPmj/VnfYS/WrFh+/Z9kWoQM9oFu30DdQskhTvLmiRvEvzMDxA
5vtTe9cY9jLWHrwxnbXBPWRZ/avj9H1/5sMp8ly5CNtgcBrAeUpoW8JZyeDeAh+BvuDosm7mjwPp
sWff8N6/ogRNGHzFzyw89Bv+yNowGS/LITQ61Pdmefe67beupKv8cB34OtCYhTbxiP1mW5xWHJye
cRSxVf568TTMYd3Eo2zCQTTwI3s5JVIzIC/6SJApgK+rxkKsxbbeCS26QBCyqhodAW54A/HzqfkM
ANXndJgvt96wPVNXESRx8EgJaV/fwvVj31mVWbgoTf3DvW3HjipWohTY3yqXX1hNj4wZVFDxJus+
9+dRwrlHXC/HBHXDKWsN8kppTS8588nd5CHIF7Y5o5Hn3L8Pfep5l0LD+du7BA2JyHyt6ATnh4I9
SKGt7YmNunn5haG4ohP2eAq0sXmqVPpuwsuBep6ymiGl9x4L0lvTJslTHi6fEfmIp/YBPNkcjov/
IUePHs0NN69kd9hNKh7t83T5tgjWUUyOiAfPE4lZNIHrvYBH2TTOQbv/1H2dR1K3QFAk7AQ/pHmu
vyLK5MRxaiGxB5EV/ZgeOctgvSulpxx1SmMYvra1BPpE9ZXJTrlXcqkjulOaQIOeGqIiPFXJAQzo
cTYFgglJNw+17i82LDXa8PqC9E4XZqEw9dblf1pdHYmmcKamVQSH7grZAY63PZbjZCK/JKZBz2ph
ccGhUTRcPs135EXSQIREVLi2Kshxeh5nchYzXCWeg16JWeWztNVChZIrxvcTjtW+9TjASU+AHMVj
IkqaP3y3O3CGVPfC4gfYt/9GEUkZitsHSiMFAszI/Aw4YoL5j7fqlu/N8HunNjY+lnc/2CxYkMrV
xW8jvbB4V8ijNBjs/aY6FOgsP65hX7xE3/O9LatHNlYiUb2ceDbUFgaTYUZFSSC/yV5fvm068iYC
prhfSCOJLbZtaF22t6Ty7xsmKB+/4QCF4MvqAQPKPHFZNYPUuLfP6jQNaejRRc+q64jNOrkjKZyJ
uec12nKIHjPYlwcJQVR/uGiEhMK0qBVWQO35zo/B1SeZoAahHdnZIjQmfSh/7oLE0A7LdnANkBI8
Ctunnk/lpDqBMPSPSyaCgq5A/zwmypjLIG/S0RD7LjfTVsEHSRtAmo0IHkhsayIBkwW21nMjD2+w
7Y8txCRHzALHpir8Sf8Q344OFsrjUzkEfy1ba5U6bhzmRqDEGQxhqKkS4svDUTE4uSqQSaLLrZON
RW2I0nOuWDCsTpcoNbag1MdHwblRBf1GPVSgYWMIhkMXkUEN4LwLSbpEh4KZE6Yk4Y+qfRRjBU89
T59SdaHih73EgU/jxHDOAyYTrrZfeFYKBr6MXRxRktElBIlo16mtPVLpUs9H9RHdPIMx78F9xsWM
9GXs/F7QYVvm0DWP0HpfJa6ZZ4xgJllI8KCIgP4HbqBBXaeB7kLyPEawxxtp+UzB6H50afX8qRSd
BvPUgSZAWDXonPOhIdU2nYIYTc/zYPllf1v3YKBShiRTk6bm+orCetxq2WWH/wP0BrXsZChl085G
v4DO6smNsF8duX+fVWk0ykZ59a03d4etJMTm804W91q9MEvpvOGO7oMJXTRjQRB7pHjsWBAbikUJ
uX6NBNdj8i0JO/PbY2vB9vxhKz0oJ8K4u7R3dmjIg/LISrXLFxKhBlT0XzUkoRuVaQ59Yl0plFy0
Y/94FjOUJqO4Xn4ju/ap5abpeMdxfc/uWHktqg0ke0vCRXJmQC2fn8o4aWaW+O94LXxV3yABvirE
KVIFAetLsbxQlxtBMIdYQ1n4d53AVvwJSEydjyT1mcfjMFaWr0c2T/WZTJUBTPqt6LlQy7xFWxpx
qmWzIv2e8X8CLSglWwGYHQZTqWMErzMf2ciCPt3BltxjaF0AD2Yy2RwSkvohfSL0VWKivdqcLaOT
hqyV77FXwCUGgY4mQ8gi0hI/O2SMES3+7pWnZ5bG9Min5bcakjjbthtIRrIYVSC9MzBk7D/0rsC+
UjnI3f/CWuQcGLwkQQ46doV3eMH9bxHBFmF5X/Q8NQ89cOagZ9ae8r2TVYzIKOiAmVybW9CWLjsi
v5NIHPscsD+rg82HLqJNoJ499ElglephC3nGMpKPeujU+jrIp+P3gBtW8mO6PUNxJb9JZnhRmtbh
fQ4/tTx3wluIV75HHCL+3uBitKGeTegdffUQgN/Ej5cfYxxE4oNuWqg2n1hIb6DF8Aowg3Re6zqI
9OXoWHIWoFoY/a+iFAH5zOIwVjPlCk+nnjW0p142Ix3XF3CyL63BgEiqYnmRT05h5vT4WNtl4wgy
axWzTAfKsE8naD0xumHcJPoj14JcO9LW9ihoM/9Bca6601xML/XexoWk+CML8h6jpxkMA501H5C2
4KZjLWWsfXejbav61PvxwilNBJvcfR4vMyFPDEj4IcQLPnb2aBioh5jduohu8OYcfUx3MjMFUFJL
RMUHa3C4EyoPIXQhEFgjqyolL5uYWO4nXbeNGxmQWu4tZl8/PzH7Kr4lbXYn9zgjj83e63EvKJyr
n550ani5LGFkI8IbL5q5YrxQU2GKMOiX+AwNuP4sPHLyEsoBLTBJt7QYMvR9TahktAFsRIrv26Bo
esh7kcFQ1cSrT7yiRgDx/lfJep1qPeypr18QnP1RVGVNjVUWOf9wHwATNl8MVXY9iOtBQVmDl/7n
dv9GtxgUwM2IZIDrNN1QqNgjviI64cJBSFqUr/oMOG9fX6GPOHJBmKMPcmz7HLBUmq5vlKO5aWms
PQ7BBoIFL+EKbVFsDf2OTCpsC8S7k/AvD/E33MPflQVU9Ai0HLAwFBUEQA1HnDDQtsFIdaH6zpCd
uiBW2yh0RdhctEaKLPW668ozpJeOp54Ii76PMT1U3GLl2u5gcEqUj4SOOJOhLdoeRmj4u8MCeHzu
/GjC8dZY7BqCcIyb/Y2szem24M9EK6p9HziuCWdwFoXSyqPNtMpiENWHXyZd/i1+cDKXyKsFWWhx
iQHn39F/oGUgIhwpq2ao7eFsHtqmGx2zOdc97wdNGX3h+0mKAyKJ5NP1DPn6DMLwLC2Fr4SKUwuT
c9KoKgraVZa7KlEwkGUBCBxW0ElYpOOetyIYri4NTlQshbdByodiLU2C3P0dvhWyCGJMTNhIIc39
D4WWNNkrjRuXXdncFDgqPE36o8CSFxC+fxS2uoa0H+BlPeIDFmSvwTP+/sqihNhL2g5Kw1BVP7HK
8r497Bn8DkAUYeRNcZIsM41fCqvt9Yq+K4czmt48dFA1sWFRTXmZM30sUbye7oF4+C5hd30jyF6A
W2EgGPEcybHxAw2WMUbGVVxNX40mIRj2zxG8GV0Ojo2XlbAgCS/GoIktP1fpPipYKNk3X3I4Wgfe
kTV1wTFkV47J12GDLESpE1H8okkNbYZId+TDJE7eYsxebeyi9y1LK94AIfa6XhJ8AIRTb5IKaDns
n1PckBfBv6XYjYL7jzs11ApGBfcGTQr9vgLLW8fodIxwFIT6SVGulx8Iy+JiVUGOdzpSkwpQ+me2
KXTkNO1+wKNF+vfJpLoQgaqmZTKYSEpHMDINwJI+cnhiXKlMdqy9PwWM0lorhzKAGB6nViXoOYQm
bDSWLkcUnzvgbbNrxtb3rX+cUkZR/T08gXqFho7N/h8KCqGI15GJ4Got6sY7fXhovGJAMqWUhrZS
fLu87J2eahmo0ojP5H/Q+A0gGjKWKGHNr5iA8YCRLYGRgCNKR5+HjqmyDAo085Od+kC1QxS3LM7O
H3V1S+9amW1pL1PSKX3HVpzjsMCJG3hcSaj6GD8TPc7A9iW3N8zy4xVino2appqhofGal+XYCKav
ZxUIzRFXqaf5KaA2OmjWdqRUUHBdclnhkuO3dUHj/u/qbX/VsiF61gQA1Q2O96R8fDcXAQVin3f/
mKtbGK0N5vWWgTUmhRyY3kC+eL8SxD2VGwq/ud0SL1GCQ3fpX9QiyyZenlPesO4gHn6FWVE+kDMS
I69SHC7sWwaGYvwuiUtQ6sstsOqp1PYlYaf+fwnvTI3ZOw6DJcbszrHDCidmUCVFBi7QXHQs081G
qOZtgLn5Lek/8iU6FeXfpuefIYmzFYPW3xZuY5v79MFioZfOZpkDUxxJgh9Tg3KIu8pPoD9HkA+j
QNRvNLg6LWYEmsebnd6bB7sbd72PC74vF2Gm5V15cAbsrqb2CBEPoEEg0ZgHvj0ekt7//NdxL+SJ
X6thP1iFgCcH2Cw5EtkqxgwjfymH+mEPFOydBlP6x8cxMfcGxH7vpWkCaRahmtMGPpJrsH55grJ9
h16mgwrYW72tK4ZBffC2ZACPEZZMak0Ei7MLMaK3q/6rDzqLQc8eDvWq7kqraWcwjE71Z4eymhyN
NT4MjIkVnsZnJsB/ofTvyktYF2Ps1rieUI7ZBcIGogUrEQ1kcKqdrimsXnCcNMLR1USyecip1mKm
3A2brSuWKrmQsCfC4o5mlexwbrPPLIxW42+reikilCC5NPwohnl3lH/Mhj32H5ZbWm4iebFrOTKX
Mx4yfrZfWr5BBs3DpAwshytWyHBdXq30H3pgQ0H1OgDD2qGLYuDiNiYLV0KyB7zs4BJJ+kv5TMzp
EDFA6bdZKtr1UkZVfglVuZ0PFtwYMhp7jfzl0b8sVnMJySWSNnhd5ZUwdKPs4SedmXytKQU+8O02
b8LndJFlHQd5xDcLuc2DQMcT27qHm9HKoigD3I7WbX63T+AJG+oOk1Few8BFC8ldZhy9sC/wGMmr
m1SjyXb24mSbhW2ScZbgUgfKayhHpcPCv191cUUZvUh1guCKQI7oCNXL02KSzODAhLByph3GPF+B
RmhaXczJEeRYaFSVPHb7FjZVDG6aEdb5nFPuD/qtzV77Jwtoi/7+QMJyOEMD0azg5m2q3Ww0yF6T
AsUdjSsSK3iTQZ44eA/RqipWkhM3usAg9q9ZIE9FX5Bw1z8zxeB4MbBGlLhVRtJRAIIDGyyp5gE+
H+cNWwSb+PuxAf+SPPLF3JCuieHKOqeOAq2H06ccrit22EpIp86sNoxyteEtXqf5H9E/kDdfkaMD
+FCsee9PHkCLRdcV4P/GXz+z3/xnmBHkhZuu5V0CU/V7nKQ5JJPNVpnHjQSQI+KjbGQCF4Mtk7Rr
R9Q2CP0lWwNOuUtT+//kcesJ84psk2ZqORqdwS+GXZIX2q8JTrUkh23xI3jIA92GZMbKhvSajVcr
71XWr78ubZKU4/oGpHyh3JQ4DrqB7okPwkKRWpcqk/zPKj6A5oMO9E+fCIiiyRfhnHAK4p5eHYrC
9YCnuWT0zPVcCsO9O7B2NhF/11h0iMhLA8RclAorny9XaK5TuV3TE9BXQJWGTc2PBlFFRQAuYR4u
z9lCUpfGQddaN2WzC86wbYRzItjSNb6wQck1ctT4xPUp1Y3bwuz/SM46itTM4R9V2b+gv9egCvoy
wJAIvi/KluScPqqD8YVTHrAMdFDIKO38JXTEGFH8Aom21F3GX9/enPQhuw4czpgJNeNPFxnNHkKH
En6eT/96oxvI3t39naYhoM1lTAcwkxGGcaOvX893Bf8pn5PVIf+7HTmLhCe0nQvMPAWNtDAUaXNM
bLr5tLGO8IwK9r65EU5StglQijGch+xlEn44yRnAj9CwPJVbreH42bkb6M9d4LmpnVZj7UkmOtd5
XwJQ2elRaighALQDzvWlN2YTiyiiNv5IzA5ReE/b/+kr/icH6GJX5OovCiseU+R/zMszDz9ups+g
ey98UIkiOLW310LKW+KWnHykpg6NtMDqh2e4unnAqDF3mAVtl+UL0mZdXgOgGsrK+sr7nhjMQ/gh
EL2w+cZIY+ppQSSADxxKxyj2QRUdtw285+wI/uK1a6IuAdkNK+4ZIXEktF//PToSgX/ok2gVmtYo
hoR104uFKtsdkpaW8yh9bNHiYyKLQVB5we7aqnycl+XqtkNZ4rq63Orr/XIC4Bx484h5ggWNQuwo
TdhtiUgBzLjtLSrsPi5etOVUu3TP0MpwHvtT/xeYp8/+CiDp5LuPNkSqh3zDnr+mW3pBTH/w2B8t
0uvaUi0ufFBekIuF76Z/gxxt9+43QW0b21PS56hXvGJKi4Hhuc8IQX4x21iwuGvjQsan+dY+7QeN
797goZfDbKeGx8Y1j3UiAl5WqRSmJPvcBeaFWmGIiMv4V0ygiIV96cLGARbfs03tAq0Ur/K3Mtgb
WqLcZpnuIAxEy9Jh1tHjvaos06pkWRN8tFltBmTBT7PujKdWvyjm84mi0P00yyJBrc0JEw3SPpSx
aCkmLPcfO+Jg/zgAVe01j9H/iEucx3tkucPZj7DollqtwtAeHGH3OrtaLUIVVK71mIb1L4DPvLri
nbwMRfiBoF6ehNXDNnHolwpdM2LdT4SDSjZz0GgAvkV2dDerpTMr10ib5EnQQTDKe5iVXjIr0n16
uQ0GbEm42XzoTLBfD5uFOmRRayfmVbkKPlyCprMgjAMorWLrUcGVN8JDoqtNWVRSuuiHqFVVY8mj
bl1wxxtYt1/IdHNxAALPovNWLhvZ2EwwNn2GOAiqs14sQk3PF0mOHZQbH6BC4ehFdj18HB39whKK
KGa5zLDOG9o5DglK+3VYWwYDJ5Zlq9SLV50qjn2+wdF1B/dOqW2cssMnGz0wS+Y4DxniQo69Z+s2
AOVrbfFox4n+ztW7gI87l3uPHeVwxPuZr8Nj1ltR0JOyjZMwtbbYMHPHCgBd5WI90w6oe0rl6qOd
rmNL0bjA8BhTVXtrUK0xJdCsg58xcXywFa/U8NgVwq2wnCz15ady7LZZnEmaX3JrPxUW8fK17a1w
K/r0PUPLkVrCVSgnkNSnB4EgpsMcgK6MAKtUpr3RUB/OMy+aWvBhOExrKaYQ02e3W43qg7dT8P5T
XAn9X5DAOTFmkPZW6y9OtmTjqAFT/aYfDNf5PeSkb/6FcSO6+YJRmfw0kBDwcidd3QRcOrWq4a2p
zWKU1DVdu9MZaO1a/D9VYGhZ7IsNM8WeiNYGEgEspsG+Tu3H07VNxqHhHr4zzqTmOMD4JtRFN1kI
CVC8Z15dvviX9O7Q66vLawV1n93dayUOpwCHH8371dCyfCl+byAqrKMnL6VqTKpZ0eSZG0mL1PGu
8upVUqlQ4POr5dBKOnlAXFdhAOfYiKkHbLiWaPzejkZ6ZY/p2UAzEGDsSEbEQ4OZVuO6Ee4yxkO1
CNAU73wpQdcjffA80542Ke6S8m/G8j0qfbqhbWCbM9kUi3bbh7q5r0GRpPmqYb6tjwXnb/qmS7N0
NV3VizqcGQadiGOge0MYFk5IW5APkLSsJTHpH1129bSQZiavQDUEd0P16py37h0geKtspobFPeZn
nYOnyN5rY6EOnuVe5fhU8ny0WDWS8ydWprQW/2zX9CSsFEPQpXBqUTjYPld2iJEphFhWGEvBlwtY
Ddd8KOQlIFymMTeg+iuPXGUrH05Bmi6pATW4lr2qFSukLJJwKKBaHlt6RaPCt1wyp9Fs56idPUn/
54spbLtx7GnkOjw/LuIjUsu0mYkMtICIRCtlR2VGGUnl8ErXBpfuzO/RZlFmh89Ie2W9T7fnU6w9
yQwcV4aGtZ5zITEVrDYWAhZVY8R2jllGxRkGKf1nOs/p/97KZZmwbYc5RmKHWQspjy/4u2ZGJE7P
ZlEWFqJOCIcc76nourhO3msXWL7z93p2Xi59vQTT5sjoknTgmuJxN9h5FWZsb5Rrovrs6FPmhNSY
voFWsVkNN5L1dNmQbPN0mRgQPIfxYpSZtXOY5HK9HpQlwJYG07xWdfz9UQ3GUVtqXBtVrtpCQHya
vczauZdVAXl+MqrAoKeST3fvjKbYUVdN00BSkOeefGkbQTE53FE/E1tKGzy17honL7a6EuS+lsK8
svBOUNKqXzN1YbgRGl3Me7CGWdype7n+Yp2xKbb4aQSFqkrOo4o0XTiWEPBPy5nnj10PobO+UT3g
dv/LTw8zeQQkNS3jXNEc3QLXBdUAB4oaDz2LZKYJ2zAdc8dBgBvpnKlmogimtZ38AYEWThKK+ZPX
JUBsz1MDwJKjjVkf4xS4INR2wymcNuvgP7N0u+kGTmarytur2xm4oj6GM6aIiFTUJuOIV6e1O3EO
Ds+6b/mgYqWRi6E7Ve0iNgiIssBsVyh48EYxVBjXlRW6hmYFCOQk3WjvdYfPjc06xu0s8l35/Bm4
VYwf1p4pfih/dnf4mbAh7J2TpAFJBk9MH9ggcNUSv0LPD1AOkOyE/yTgrO5mGZSmM0dc3y+cak4A
aBKQGCkjl0vsuKRjgqh20ZSF5HicNap6QILiuaWAqyelpbSVF1IsZweKIUACgZKGNoe6eaLaW4y5
vqyBdlSdI2B0pOAU7RdhXLosPRTcdZPyo8Ro6otWabVY1BfEmA2ZPuHl7BcgAqT3uP8gupbee+kz
0K06SikeqSgFDKIIdOTCFLoxcNv5o+GmZ8MVQr7RaZ6rRzRgsunZKP+uij6pMo38hmAgo0ZBsMy+
U1f2b2daep00w1LksdBQxGRIHFonez11t1Fub5GS1qKmZzqS2eD1J54HtktLFSafOD+sym0Loku4
X101xCOaCokRpvD6v44ZTaDyK5koMQ8LdF2wXTUhx1TrXTlrtc6rr4n0A9GnxBzGVeThDlxTMqMY
OvKAF8gDZ5Kni5hucDJkQ+NKTPwFGktYgVPQ+PRCB3Dg/g48q9fQwvI6Sg1MOpHnXS14Lqny2V1/
uidb5sX21JD97vWydXDFJt39GSWOyJ1sF8SfVwAzCf8465USJrashxWYJm8PdXmFfqqyTayfapjk
JNP26HAXKldwhBUduocXEDseQdaRM6zgapwMGA5NCEdl0evUfGPYLY5ZGy2pzM6dTH9BKgAXNPoS
qLzE7YHWjGEjU0wkfY0rXlPQccOtMoe/WDP+X6HdBZmBbUVVI+zZNgr2NRfTINrMUhKlKCTojFKr
/AjRSma/gkoD0N2pP81QZEgMwzvgC22wPri33o4AQh7HHjYNebuIcgarh8MuVd9HAcJ9e3K2aN7n
hYje6DTKsP5+TR/5MhH3pmZ5ck5UrSgrsOSLJ+rGiMSr9WO1NZm168tkY/nIXUfaEAUkVa3ll8F0
12ctSeP9OmdQx/U5VK53ZPf1P28ZB7QIykX98iYawz0EZ5CUqZg9ECIFXzzEy7nfoRKP84zi7nPk
v325JSoicC4TWmZm3sWhpc822UHo5YwO0vrE1vrACbQ2qrBHODt2/6j7WT980bWnLGcM7/Z2Kdc5
S/agDrxOYSf4rAYWtVuOpbyXI5tVZMlnHE/tjtZWJnFZEy3/Dwu8E1q8J4cgTLcoizPEMbt9bhCz
gx+Mhy3k5gvEtcstFC7KOuLcZIkHHS+DkiKzwryMhh50wRjaktnllwhoSPdU2B0XpjCWczTr13+H
3W7VKqFp1ZwIf/hgNuzwZhG5lyxnkV2Q6XP5G2qeT+ZHjm1u58KLgOHdoarQu2c4PEOxo/w/odbg
4Na1Izwhu6o4FAhoMiQSy7oUCbEm2oW0cfmENcL+pyg4+iCSDhkSiN3s9BdRvZ1Rb4qOdb7H+7r+
9nGRYjCOY/NDmgJ7jrQSboC70IsylKfTLVljtBTzHqbMCu0hMBxbEHn2xZLMtJgtTOWj4DOWXdWp
iiDQn9PzDnhBJr370x24LEK31x3BCWnseCfSnmKFpMYgfXpKpXDNs6W7/giaRGOk03pKdurYomkj
Fh4TqUb3ZNTIGtkpJzsuAvyX0bWiW/knHsW1A3M2x7IZs/3bXSTOIAX/pZKuT+wbm3OIySrR6hEt
xdwZMrs4HyQgqde1w52UqEgrGZlnoVJu7efoy9zuu+zTIMgUcnbW52cM/VIyLFmjvvnZzSxs1y6i
6pOd+dPmE6jQWOltfk01tUAUZc2MIiDMPwQvd4frI9Vecw7WZOCZeDC2bmYpVQz2vAK6+06Fgvfg
kNgVa6QS/elMjRbjyyztKRg7tWFZeu4RwcHJKJNmIr4bBFWWJci4c9MQggvp9VXc8KJMGTv/I6p+
tGvfh5QB2lof8XKjdDUGwE6L86w7OXzsJKafmv7rUdzTFV23wYC3dcO2JzFYMcl0RDeaHRgmfm61
YjQW9MjqGs5A23KA3/xOZxN01MzprGqYRfnZakX12LqyOonS1pBQaoq/SIfxOeAhfYArERVKhTe7
1oUt7Bg02NEyRiqigjrBVJIR29BSxwePIkBMRWrJsmNUQBO+oXMJw63nQfdPFf167PHz3Sc0CtAx
bxLYYZlTqFCE6n2CVpFwzAn3YPzrc+RWnb+5e9ExLsYT1/x43WSnlDGuF70AakZm7BiPG6CWKOOs
iQRy4TchtpPs1jYxu3LnMm+4KrRpcSOHTqU0trGcm0SwBsuCa8e2e0bqA7XM+GqNReNSkE2gvgXm
ZNcz/CbJGCHVAp4CTnv1eeu5KioKfsoyMZPwhXw56TFSxGGqnOMYFGb7Uo6DKu1oW/P80u/EWyrQ
QKxlcJEtNX4kwXJmo4IS8ugrs9Gh/CyXmZAg5HYpqwhGKTszr1Q2u1OFF/oFB24++Bizj2lUy2T/
YNJOUaAapdryRX06y95ltUkVAAYDdeIMzf9GscWpNtXb8VbvoTnmaYPFT9ke3OUeNLfa1rSrRpp9
YGSqnNiUBdUXQl0xfYu6l4fymjSHekMErnYmdaqSToIpK9DFNm78jmyjPFvZDpA1pB00j/GMaeFb
qc0FJsmAoyybxNDHErKX2ecLCjuQtj6dHv/VZYAe4EW334tfqbDFAhSFKrwco28TGlUJ0RMRx5rv
bzrWUVSP9ghOy3/0LXrgsFimTiVxn7Zs+ExG/9LBAWGREiOAKo/1Y0WwsfA+qGSQd06x66iGytr8
qQwWhm1AoKW2Zipjsibh9tKyWb1j+0wXWOH4raMYFDAbQWUMGLIvmNvLHyrwBqqCwJgFl2oaPy+e
SHF8Wg5eW2lrQ0zQ+6ix3PY+3NmRXB67vi+IkpSAmgGLfAp7mx4jhMSd5qG0JDfhgcEdKosZpXVT
lizOJm8au0tfJMFemUrDliktSERcogSbk/eJtOC9426B9X8NEi5bkinBqoVFioNFFi0b85Y1ODMe
3xUyqrhRAVtgn/VSMVoj4doUEatAsbu0ByFwQfJXQU67XjW7s6Fg5X6Q/AfpZfJ/6vecpLsIya8H
NFVC5QLxOr/oDrnEQRAZq27IXNrctX8Ko42UMnZA93ybt+y4y7JTrir6PWc8qvgISBPrusgH3Z0F
kX7K4cSQ8Cdv8hInXI6OlH6BfTgAXyZVOfN9xx6E3Q/UtqWKqyqjcHC0w6ftc6bjwKabByOOVbLe
e54JhTIowRu9xEi0T2WeJ9hN5+cooBOLuWtvJ2sZJnxanA+bke6RbdcdpOKRtAmHofD8FNakjhb6
JlUt95V4QJbxAoV1hvuX1s2ejHyd6BTlf6ZK1ZfEyujnw1VkFwUHCd3rdzEANyMnwCPmaUwej96T
gCSBFSixWZG9aZe2hmnXzrNX5XXBRMUVHd0rRG21h5geN9XSJcfVjSRNNrFqCqld27NJyqYHpVYP
ggkmCHXIwlvdWVYhyLsn85HyP/tPjMAcgEwbqzFuOQu2Cclu9C8Sc1hDMUMM6GRCi5mWdSnJpxit
Onn5UiXDY56l0U/dey67JfSZRz1gMWFpAHRNT47kWIiDx3WD3btCg7iNm69yCaFXKtNU7hjF1Qtq
KW6o4PGu7HDjYUEpk/6rxutuAj9vy53kxg6aZsnll9nEw7moNJ8r0KBdj4efILIfWofwSFgZza4r
1gMTUDimOPxl1YJzcszrTrtK5A36O3Smei2qMxdOSVUq3iJd9FFiZYshHDla5k+sIWFkJqTS3AaA
8AN34fdScFLYQXhg0WVvH6cVMR9FIPYqeoxZ9zRt+aqtc5RN0OUzuGFfq8cSyU6RBx7jL3vzTnsg
cGWNdI86SlKwUNSWOIUMcCw9vI3QKcm/Byiet4GWOjkLxDL2LAiB0/RzDqHKAbkv5Vm6St1T9wXb
vsYY2e6X2Ibw6KckPRYaHkH3oYjdgbTi2oAtKaT/33y98ovQUqLQlLbrqN30+/W44sM9U0UsMuSt
ZzV2OsD51nfCR9ed13wjoJdgb3X7PqTQ4mmMDNRA9Stk8E9HMzUcsgWl+1Cb3XTFaV4XH0QAWeTY
YMW97i161LVhaKE1hH54NACHUaYr74EvHkJrky4LKmee5kaax0xNhCeafsHyqnQFQRhqFIIS90bV
6D74GW4AGdtyo6R6C+KNynHFoqliO1drkRoL0UgKcJfyBLg2PtGsnRU+p9Bxi1xXpAtRBg9/z8EF
g0FE7sK3UpztDV9QoxlY0Bu+m5IvqLeDuN+kiS7UZHFnyA8bbzPv+gnuo9+qfeRJAxapFltkLslz
mg/UkWsIPs61oO1tQzYXaLGp5CdzGTWABI2VMznohgxYCDJpwgMWcFn6s8btauY7dkXL2wI0PBR0
aClS751YORUsg3ek9EkRiahQuEORymiWKe3acsweWEbxmSbXCDN+NgqFOb/NANsb0BT3AA3UjVRN
1FW5sXslYJw+SMxbUHX70XFNtqdSxFBQpPMMJlkVEYq6phoxqTfUja/BIUvKXlcFGza9r3yeQUvw
wSqDkZKNPo2rQtpqVx424dNZ5Lfo42Gu+LOXYRDc+b9yF2BdlsMaLqt71hI8tN3C+riRHLnSaYJW
Zcye3ynPS7lgbcTxb8v1CFoPSsGctbxpTaX1yyEJhCkH/syFAljSa9f4UDWVSfbo1YlOGGY6xtzl
GUjsmk5CY8sr6FgMBHXH+frhC+I9dRhL21DD7qAQ7oQyanDP6Eg0YAoA2zsx4H2ebY9kvqOulYK6
9RtItJEZ3o4sqL5DIfFQJf3l3hD4x/OO5hR1yztGJiNvfDJEJOy9sVdGK31UKzG2VHjJDwaN4db2
HLAT4ohhyEeLNPet5ncBDXbb0XbBQDa35Fa5Q9OHQnDI6nGZySGa70wtDm8MOtZvXyPP+QWkhjNZ
SL0MbJeuxp2MYvS6VcR3tFIpqmEKcml/DWk06f7DNaATiC8hS6PUd/C03cTjSNoywpehRIyD/790
1D2Q/TuXtDSiiYLjZ32o8BSRbvn5kYSA4YAZWLCJDr2BNQBMUBL1JLanY/upaxRHBUvJhnbiO4aV
jJ/Rhqa486syXLF4AVST88i78WWYRgYASjNfpGochKzvtHa/LVo9LKNx00bqL1lIDaqBoAm8bx2v
yZ5hGkIFTPMTQG6vRcFAGSRIhTRwRpKONAwkgMyqdzZMdzd0Fpkgd2BGKHD1ScUg42WI2VS0sNqT
CuVBlYRRnrQwxN4b1O75iAtWW/pBKmFAem4vl83m5QKGYI1b2w5ffA3XAsjrVftL1/y028RJNUNi
ilmN5IawgNkPBNHKtKrPiNaYZlDoip+CUudgMARzk1XnYWQEnAXhMqcdfsznWlLwr4OkT2byFQ/H
fUW7NHXA6l3Oj3iMsSKBFilds6Br+SBD/4bXRE4Yx9xTpKS3BEcw53owQnquPjwZm5M4PhnOmlHF
J36kZM3sgHUOagy+cdvLLRJj/+NavCBLl3IVuzahKMkemXPOUA4SYvuGDKdI9Bp1iUDEFMW5qiQY
oVFEd2fAWe9YgdDUbkIh4vHUo+eVdtYCgqG/oFr2qyPTly5PSm1a7WEDbsbO9iMeIH01SRZi2TXI
9Z62JnEUEBr+Ekk2k6bbtMUlfXZrQ64/0jTrsW95ztho8ueryHc9GwG8gq5vI+SQ5/hMgmSLccou
Q61iuXU2XGX/8pyGLjWWLzK/k2O+HKHz73xJaM9rBYH0XVMGGkYV4Tz1gq/hdOf7QHTTKpk5nF11
CMbQqXOCUFasXYH9yggghvESV/6NGmjx30YLmE/OqovPdGtzuELWNaXtHliY/jRM/+MAZmgS0eCA
JEcBW+OXyVCl6Bl2R8QW4p3eW+zbTSICwdjOicHfnD1CDzqQ6RzbsvZbwG3mmHTQ95ltQCc/jPEF
WQ+6LuKv/DGRX6YKoISr2S29cY7bPFN/zcEMWzBE551LVpJLeSx13Px+LD5/4qhtRcCknP2pwrMA
jdt5HDMFea/nuZaIRSUYY9Tore9wqX0RTpoFzljHTjKVOsY3RBPWex6YoMYMQES4X22fu+m7rgvn
3NZs8bJc+O0pfLPWtN2Kj4ufBUU9Rd54Rckn2Eo/KU+6LKlmXeUFWgLEpRQABTUSO6zriRN2cqxB
y6f94kFfSwNBh4g5fSqfZ2RLB9WQLtxcXOtcJs9rC1CdwWJd6AJztNYYS4s+DXryfWVJzJAy8kYy
mZkIrjAFo3N5203f6yyu3G5UBgaYswDSPatO/9yqGNTxhMEGpcyAyO8Em/BaEEx1RHh7Zs1AY47u
uO5XUqktHwi/hW9XyCVEivAemz2J/8fkJCFVBdz1fee2bqQXVta9RIq/+xtxVzhZbF9bsygfkW5d
/x/uxRDH5+cBH8ESdUCJHdXIttog8Y/BH8lcSqUvs6LdWS0+pBoupP9VYk/CgiKHvLAs08Ced5+e
IUVjZNk7MayFiQwAfNh3PKsH8aYUvLXcB2It4oSBUAG++whTcoobAOJ2PrMePYEXoDj3JZrPX1E8
ldNjcxM8OKKcRIFyTrcMEH0G+2wsbbmQLFDia+8/bslpaREi4K2Ua3TMTSVeAHq+KkHN0JwomMWy
IH1vEWjZX/JUKH3FQm6i0d0hwbnFROY0Qa6T5EVJ1PW8D8pVmZ6eqb+EhQq0OharDPSAmQqDX0gK
WR997iy+iVgI8Ui9CEBu0ag+XlMURqH1gEVqJKaSBvtxVnGNtzTcdmW4aya15sa1vK+a6nguqxEP
+PTxMos74pflbruTbvsW1s0RQhbpMAbXLuiF5bFG8wUYOHC3cptTgDj0IQD3PIO54cpThjEyw8Ml
koUo8/NFsuuYY9TOn/i6uMSqJjy2U7MNHHLN6Ec65NNNUUCChGcwuF2igyamfqWOZRYv2QGfU3CL
TsyX/M+M6Z/V0pKUGTpOKrlAVNfTzj7o8hTaTBMTPhlJirO7xTcZ3qey0T/Z3kZ1a9HE55AaeXRz
ttzM8mXjl/Vo84zBSgtdPezow2xAjl7hZv9d2LHZcHiHC2W83HHiyQxoMonmCG1eWCsLji3/jiMS
Edj35BugP8q4RWrAUC1/LVKMGlN+2V2+Fp45nbeeOOxPCQoo3GDyH/dUC01msfNosh0UEu8zqWKt
xzMaJehQWZ6wD31KvGwr6KubftW1c5mScwYB4i7YKDI8xzOxn+J32ya9zx32aLN/Bsg2VhmDzqx6
nHSKoVTZvOFE/27nPnFnPji5jhTzxU7MehYFHsyPUnBfA/f4JmL6xtASGX+JOoBbx/634qYkf6D8
2a+QKhdqxFO0um12AxYoB5jVSvLNGS6e2Zi1lRTDpUZdfCw1fkt2zqD2mUy6EFf1mscqVkE47xD5
TSa5LChKbOs6fCNZ4sgB4vSxzF7327P496wpYkvXI6I4/SQLandPbvkVCTXlJiXqoER8YwV8yjuh
xsgWIeMjOTOCgqugh+ajXYlpVysGPtvaPDKTnrUKnZDMqMfOqITHouPV7a4HficdHxq9Zq9CDYAv
UVt8J80OIlRXRk0BjMe6XLEu3Y7tdbnfQlY/mpN4/KfR6pzGWsi0KXuIEA0avNVg3ZoW9ByGiwAj
hrQd+5Wl5q3LUA6mmhvrbjXhuN0MjqoK+5UuWDrkBYgNmEN8o2ki822jjsgOVb1bpP+zMGV0AmL1
Atgdo0Y0XSl5IjsA6dICimLLP/w1GgAgmk7RGveXoPNZPav/5UH72th6dH1r0BVEF9FPob2Y+d/z
xskwY+aPHGgMChtIxehQ07Eap+QcpNhUc9npD3sjp4tBcUBHFjmwSR02F3+R1RPR7zQHDDq750vd
YbGhAdnPbyVPZgpT07GDn4WTkegSZzFcfKFR8HsUHlThrdKvGzgrKvJz0rzsNWOLQJb7tI7aH/vF
hTwLDQ4LrTMVQD/6eCm8xp6KdxmBd9r8deMalWXCZnndi12PuyTfCCBrXuAJsP7GmjDOPq1Ppaoq
3u7dlyfSQv0g0CunlhwfDoSSNGNDv1vxkTrfJYiUfre/ctGDJ3mYAqyvFTGS1xydhHnQt0GmxLZH
RftU/0oWRMqST6UanivpJCJCcGrfpH+Qd2MnOP51bSmt3Tb07pO8thlG2hqF8R/aaiPQcFykBEYZ
E18YzWcolt6GuzVVo+P7Vb2RaNch5QGjJ+XhQaAC1s3zDkfL118oHEbBbmCkVi6BJIAdVvu0SGbm
Rqhoc/2RTxqvDByayft4Q2BnTS/j94RTUd2W0t/EtxQnYtRZrpZhPZD5X+UCW1AW9K5w9/IYvKX8
QLneKo8fssXUAuzHwC2Fbg/YX3jir9bT8LUel7eZ7kv2SpMO3HRFY269l2A1S32ahKxa58CrpKA+
9FufrGXGkm60BENEtvc7VsWG/0465fp1GJP9Qd3ZZN974w4C4sYmMgdpRtRw3E9btE//6AB+KAiJ
bvzkGf+Unwz4BCXkJ53CoFtMz4X5mEkDHU2JHtnoZcZHMeHPAwagnG8awkUqZeBwOhfroibzjxtg
kSjYgzPR1ULJQS9PSAzYkJp8BwS1n7HcWdOCHbQ1gNtpXEAwPfdD9sVPHVc3BPa1vhkYqoewKeId
HWJeP6HB/1Mx8abF2imTO7VFYNMbLYNiC0eWfUX8INRngbCmwa3Q+s+LeivhXZDrVgwpgF/fCkaz
rySk3GA9JxmZgedV+6MK3GE0unU6VOAAAnuBIT8XA29ZvTtUt5Cp39tr4Qg3Rm9SH8ra6/Kg/T76
iJIlt+OFO3q3hWV32xWg8e+29sD+OsoWP5M3xJoi7BrVLXd43RYLtu9fNhlHQp8bq/vS5BSLOF1F
HqhNRCJSoE6or4h5DmnmyUmBiwzTopSMesurRCfBzkQ1DWtu+3XRuBZ4BOuGYd8F1oRgNYdSYn6P
6ZCbcA9TqCeRrMW81m5o/JNZOoK99QOM0BkV992Qq5deE936QZ6XOtG/vKxpoaIm9I1Dz+RRxX1b
u4EdUhXefs7yeH1offCpQ5f9IVuhVo1JRSOLsF4SnBEDTFiCqNhuNGPDafKTvgfOTj7nAMXj0+CG
HkZsPoQ6Rd7WOLwS507JD7QgnGcBiotatUmKan2Ukkiq8stCAXXaRUZ3en/+v1gBeNj1prCvx/Hp
GlW82mLMn8TN0qCQ93DLl6WyAMXzfZY+5VHMpY8MNp7Bot/bLAgXqQ45pajo0gNXgc2ABPdFPL03
wN/Z1jpP4ZQaI5duPGw/tM6cYnfboShOCNNrm3Hl+S4mpzC6emmv0nYes89jmkx3khxbgv1yOhB9
eTl1RHJE7CKez0Yzuw2GLV+AFrF4l8HqjMBOJxkyCUXG+c3/FmD9PaWhK6z4T+vy5+aGvYzno5Fm
LM1NkPEXgEfRSYPgq23EurtzxPzJuFUWKDPv1HyY/+rQdUlMxy3XCNa+jEe5YKGjIkBE6X2e68fe
MiS2O6mWCXo6JDW3Ty5titGQsgqm/FJYzoyQUURet804+YfgQOkfscLO6L9mVHKzljMmfQ7BcvxF
LgEbnL0KdmNhsMR/3rgsbjL8INruNx36T3g753cD+lwzHHhEsLz4a6T1UrtaZwmmuBWzTrDw9PFf
s8vo7lo+z6KPVwZPaKxAMcFeDtQTUiMEbp5BXaCrrq7W7Ww6cHfbYhnv4xkAj/axzPDo3OHf71q+
RwGKc5LAWRiXdpFaFbCqbxAVmYMfCRZlvWUaGgZGaicu7ehFu8dxw+Y1epNxof+D75XkDQ3swET4
KWfml0KlLhs24dV+nk/UBKwpPMKR4+T+91nP9OQtGgU2GYkUFps5sOBHMBOtOwGonv2YD18MQ5sJ
+53Q+Af1dUf/gT7kZ4pkhPbV+5NFE43pM1ud1UiTVBcv3ETOe5nxlndVRv/4xB6oU1OPIxk/SUby
kpVSB6x3DuaEaeRQfGmLPxtBxB+1RfAMbVf5Jti96DMPgkuOwgXGpaeJ4b4hEnrBgNQUGferfLAm
wNnW+fYiNuTOazFFTzUEfBUHpgGiuFPOXJV4YPo0UtG9eh96n0LptXxRO3mwXBbgIt9q7iMG+rRo
aeS97z6M0RHwjlXXnrTBEpQBrBgzxCADMgOThlIohRa6e6zSl+8MsGQZAeYPlIVUZA89QdxGNOxY
UAm14Eux3YoDVgxEWhajvyFT7UEiqLU8hSvR6eckD8UCR77/F1LGwp07v1ZysIb9WCV09Dk33SOE
EEjwf1TevArcER6B+z88dCxJ/p+0rhBqE3CL0Rg1S2Nlx6LV4UcfB8OR8eG7BPvGq9wtCmKV8/xr
Li1V2MsOuI1//X6lr0gvcTbpI3Op1iyvI/wC7XbtOfP+/ClPApZoKljVBfS0pBbaanUabIkWi6Hz
OlTJelrVXLhLR4cNLzipgq2Wjpb62Li/Q/kL7+HiTYrEvIPJ6bzwxnIGhhXlf0nu6U1I//VWL6pk
LEg2IKpQCcgOGlp3a37OTH62AP/qqzkMo8RHmDJDuj4BKY7NIW0jFQU7AaA/ywM489Ftek0hHIMx
KnHUQfpl5U3KtYOlzAjaQhrYAxmFThC73ezUaddOSaZxk9EZ3AI7lc64MjFz51xiucbko9ILcmkV
tj+V9M4UAgPccBZWsuNJQp3LkYn24Vu1sCdrfw+DZc/C0kWX0f5vNuAFsS50htMzEtCAstGbJzUD
iwiPGuUtCg5SWGpGgqXgQMvLTlT//8+z4c1PNfLOqY371Qw+RfyOO6VZlx+oTfBV2CI+ddZ7m77A
xwQ+XVzebljPFbR2Uq1NkA3/IcIkSsQtWYKp8Nf2gsqK/4mUxdWZu9O+hNFPJMZ2i+SscUmzsr19
+xrV9VCx7JQ5+3So9J4Os8Mz+PG20zEmQc162HjyBBf4mQHG2+hF/iX2XdwD/nGt1odp80iIXxgw
FilxtcF04WErgu9IaJ5BH5pRoFwhgYvOd3A2U+rQV7kJscYviG9NmXXqsAGcYE1wj1kCjPwjEprK
shVH9B8NiNovBPvs/1IF+f+SBzcLUqMw/ghb2D0BxwdCia/GBlLpZe22KNDyNwdkc/WpcI/5wpvE
VrJ5TR+fDVf6k7DI/7N6YCT1ResEvyB9SYYUQQinKLjjhZPpqQi7YAbUWZGlmOZfnFwUZH9WUukX
KWqSgfFhQ9198Edb0I0je9T4oqzBpUkmc74lbjjl7Mj/MBNUS8kdgkPUz/BS85AwMSO/YXnMP+w8
Y/zYQGamrbDmYzeMDzZd/2dnIiM7hUqrQLvs9Cp2jb/4jtM4esY30reUOvGxYFTFRd7LKjotJsHj
gBnY1gFgx3bGCV4nJNjFok30StFFb+LCrpFD3tzUk/1fBAcUAcw4dsu9B5zblWhPw85sVoVlMgXR
iwkq0v/g907meC7V9xwRhvTnPCKmVyOSZaM8qErjN0U0+Uu35aaiMkMOTalQx1BbZk23zCDaWu56
VsHCwwB82oqNK3RHsN2P2pHYHkKVm8T3DSHn02g5mgcbx9aGjSQ4y0n4dKiI/a49C31MlDvNp0pa
W/P58RiXLVQjbXQAzWqiXARTVQrirE67EUvtsrYN0PFsiih1d2xHaEc53xe/YXG3ns/RgN+OA1Es
Ckzsg3D3oX9ribQ2uDiNKZtaeTasEy8NpzzTIAEB8bNA9bI59jJbRhrjr3o+Hw1lOcvsyTHU5dMb
WIDY1yttVTiHrnKAk6yOCk0oLyWiQ3NUca4r0YbLR0TMoV7XAnH1/vskgV1d9EjHMAfAyd39Cnwm
aocVCBZk6imanjXuI29+esbYQk/sUcR2ocOj6TPuqX8cboyJWrHw634L3NR5SCN2SmGHQXtDU9WK
YhOf4Ock4IDrHFOzM/P/4hhkY+qB9uytf/fdKC+/SSrM3zgThowE7Xwns70f/HRNH1nihVWVbtUs
0zfwgCYSkIukwdpeKuk2fH29uZKSmYNCoGRwIzQEOYN89gN3UCiGIvBNfRVAOkRWaM7jM7G167Ix
3DZTwalSlK8uzlxhttzxLH3YL+Hbr0ndZWUh4STXKoYNg6bm8aJgrdVJY+3q/bBNoS4W4RUn3qXI
jWLSd++mz7007p3HUavVPgmerEG8l5cEA2PvALm04DCGTI1nGjjZfwmODTUoG6etL4qxTaL7AZI9
0elviY8NcVMZTb1qgR+SYd/P2B06+lxeLNKpd2UoQId0e9jTnEug16S+m+HC2Vo7vZGyBzVaaudL
gKgudeRDaZUTH+FKlA/fJTIHzt9BGTtuy54lzkGwBN6b0FacMMIcv/FBUEIsAyozfSBDyVVuMiVG
cS+LPyR13ypZaCwwnD/rTjctSk7WzV9pOxobnedfzlNxALV6IRt2ek2xw12hK3KLLN065AYjBIvA
u8JNgbVBr6+xW9TMQ1EzkUGJXgzVLdvV3+T+g7agu1PqUri2pfy/MzsLyKcb17MPJK1fx+u/NMHO
0bTYoC0sJorSVfUGmhv+uc5y1UDygTdnnFQQlYL99K0YJ7eDNtK3SMVNkgQkzYn3/Eh419TCHOpV
CQd7nWSslz9QaClmzK+D2HwQI89JwqSGvfQn+dIy0NIwt+AkvRoz4UqhLA1m/yaBbhFAc+pqYTlD
1AzF9mu/2P/lwfgXIfGqa4qzumaxPcUDvIvepqQxHN1cWjzgjb+YbmgokPtf3RMt98LQ1DF/qczo
MqHnx6LBNZLpJGJl01vc7wGO4X3KbKxQyCilTZcVpSSqWgoMUu7Kn6vrhzKQv61ZONy9U6dsDTVP
UzlFAQzYlbgyVoc+ed7uPAobiYYHOKrNNj44gx7/P2O4fM590wM3y55jZEYbmy9VQtzGwE7U3swo
n3kTxzodjaTxDVsacVFbraYzYYNyvF+TFdrA4YWQzp+galO/DatIeoQVe8o10nP14bVgO+Yzfn1n
stQbsA8dtA3LIKV6ZI7f2p2lUGf3U5DMGpFmEzpcQt2XRyov1WiRK7IltkWy/ElZ/MiypN8bkuuH
Xz1L72/KUPbtX3oMDjJKRJCHGpZC6awM7uL/5MQIT5J6VdB4c63aNS9wnw1rD6ZjtVqm8tBVZG4l
X+yfPDFkmyVqnyndUaU3RK9yl7ZHGWJ8FkUGXFzBOJL7xlLHDJkiwTWpOghrUlB9zJkl3uvHUUGi
uUfx48tFxCYmPMLko6J1RdCneUHKjgD/C4RQtZbTi2xy8FZaJpkqgXA74S756DRM2YA6uWnif6UJ
EE079RarjpDq1F9a71j3B0rzwrZA2w/niidX3Ks1KueUS/sTNUfUQPQcv/twUKCo2/hphpM/56Om
8URF2kVavVTevHTSxZ1XyPs6w9/3Qh+YxyisYOR+X7PojD/+CH0WeCfYjfhZJKsc/3ZOHEL+QeDF
dEniA4hApHCtBlRz64s+yxmg27wU6oyM0iCANgjcCpcGfhdzwOBqgUZiUTTI5KflYDIjSrqhgZOj
vk1Nr7AchtKfOoX7snt9euAMk6zMWm61HvOo2gBdo6Ywv7/8U6HS9eQYCGmH4TKiPWEMFPeFvr2u
GrqVT9u3WgG4XZhrPp69w8MPxCgz6qrGVDYq5R+CZcoW6twATC7RsuKXJED5hY+4Yk/pj3WeeX8D
gFIVuUJ/dEDtHpNYn78fxdnm5Y2rUH1LLRWpCVzWiSF8+o+4nMxd3FC77nHrQQt9qnfwTVGwQ/WS
RXRPNCgZI+626WM8njGGqBCcgAhKdupvXvh1SJb6NU9+FQtMSEzpEX0ddV0Eld7ZenSRwYbCAFSt
vdPXm8G5LertzvEavgSRprkL+4XhEbIEmfHiH7Krho8iYIk2kwAi3cwU/KQNKlbXWH4oNSVvlqTM
5wSwD73nyt3B3H2A5dEbWGD4nE1Ia/u1XbywkHdv7vHlGgEVceNu1rL0kdgha1xl6hc9B18efQYF
JPvz2iAdoAr/gD9Y/1Eglr5bKWlaitwyeBB6HufaJel0l8YYWzvCkXuNOo06pzBJ5LBzGXx177Ml
lG5NQtOQiR52ZzoQROQE0NFxbpGPlKJwhJLXdng+Mt5THl3j5IAlyuT77JphmJ8q3DZPfXxacxjQ
1HTE4183ifbCvl8Bx+ILtCw7W3fKChLa5AMLiuFdUF05zqaUpjjNVZoaFNEx/jdyX+AG1GvZJeqt
eNDwvZoFOrcS+gPef4mLUT8jWc/ffAk5s37TCiy82TGu6S/dap07uE2cMvgs8XWj9rVwffdj6Xot
HjxdmAVmFHmZdJ8RlREg4mc22P1Q64vkBSoYeTNrMYEtMm+VxBBux2sxmxwloD0qXt0A8osdtVkJ
i7Ht1aMAo/e0F9pew3mwDGL7AOt3GDLLZCpLxbSWqQQ4/GJ7asNpMQnHZYyC0WNowdfBxhV5VZiW
EkFIqCNZGltQiU77D44jWcpgQbvDpR3nYi4h5x+FA0Y2v4FZdodxE9LXMehENisHAQVvzExWR3ju
ajwe/+k1iSESkvGKHk9dvsGLYvpt4CrF/tLr6N9dQgS2EsvQh2Ga289BHi4sB+NoHOJ4V0zuvfx6
bkdMFjFwQSHeZo2t6u7VGgbq+s+psbCX9BnmmYpiYEidY7y2dtmin5FSHB+xSfDIw8roOgx20Xaz
aeNlUEJNXdZ7Px9kJP0hlClDPOa99uJwLfWtEJsjXi7LBPixmSLA59/DpNnslNfehVJOxqfV4tys
6lWF85/S7dlCaMezopb46MHhPOiqO3KlosaHXrt4EI3YPoWYcgjPkr8MHX9s/79Uf36syhEqLsjo
q0+iHmeMgbFmTn6Ac7or5bRLluvCVJJfUcRtxjwpEjRkIjl362ESLfIElyDLTCZEaI/iC+XVKUtL
6PH1Qff2apWf0eSGfdNUX2Mpc9JW3rx7IQb+45T5rHbtmDpBkeFPraXB7wkWqLHiOXb8OQgOn3iI
03ybZvqIML9PidRlt7m5Z+W8pM+v9WISWEwyvnGmmEeYRnBm6Ecz33BugfAXy2L1KYxI50C5LAPb
Fgh/YWQf7AibZXJksenQ7JFqfz/78WPZWii4X3gYcIuY0V40TT+j0EvoMSQiTk5Rx+chbVVMyz+w
xJjPaDzor2Hc9gnjbM+4HhyDnlLtPrBRX4HOnI47YDNym6tTtkM+wwcixhbsGuqd5AUKb7FxvywJ
M0lc9jia1GA1QCSUaYSNP3EuchEE9d2VndDOWeYVrG95q72MFNAPofOZ70L2quMBlvrZo5FjsBAH
FLZgM8OdlsXKxA9vkFJiyrpTDWH9RyYcfxGqZdXZjWnF7GMkIlWsdr+ZrFDQOG/ocNZaj4N4Ilgv
RuTId/E+ljxeAqgOw7B+mBj3M+S7TU4bzFr80VbFk9SLQz0jGO1kYhuM1wv/VohDMvQAE7fgcBK0
oy1EZwh9D2JTArWwl5Ux/DKNmgjh+KuUiUogUBKbj0n71ds5HKz11m0h5sWbh/Zt9bCHed2xsZuY
Tys1xpIKwgg+71W7Toa1BqsWrr1+daQHGHxVChog/G9d6H+hYpIA3fdah6A8UVjJ74enecovfKis
21OtGyliuY75CImNGQR/mpUrYYhui/thSCBwKuU1SPvWQHEEisntWtfrJQql9q3VI/TqvM+7/S6S
Nec3bI/J1VjPdU3IWWGxuhffcsz5iCG+2dFWLzt4bAseDMLhbMcvEhqgXw3gLOCsFNkStF1/qtjg
7TZg1ELJaoT6XlxpqU6MLwY4o83mOlhB5pX0c8n+mj1h7DrZ1GyhVMdEkFWsvh+JyYI3UluzE/d8
Y0vJs0EHs6fRdfTrCTj9/2lWjHAN2raoFx5oXLgVnSkAWWb1dDi0xFyN+yY27WWbUBZ/9pJqoF/Z
LhuDquc4TNlGIfZxd8EASGP+WU3uImD9va6lC9OlLp/3DyUdB9C02mNZ2sAlQFAJaEipqw/Udbvt
y/27pLu1MUkXfIMF2do8AUTFpqsTzQBCg9lYRnfma+06Xk2CYMxmKnEUUPBAQI59HT4I7YXaN0Wi
zg9fsBMw2bbSNguI1Hnr3vCMHv63mWgELWwgU5wj7MKwGVXin1lkrKTvoUBbLqROka42wX9QKKXu
u/hfQn6jaalCNfX0manZqmM7iF+R8ioiTiI+7PsIIXmtHbf4snAhPvaW9mOue0Tl2BoHMSven2dG
j5UMoYncJPGzrRxdXLp7r4hVIDLwyCI32jy7QPV2zcsVw26EeN/sDGCVakQfTx9MxNXM27CRZWAv
3oPQWoMwe2NohARNdFeYhgZv/bWdVgKJHHjq9uQrkTjLJWN9wx25NgMPwGCFJ8G+oGidtKPwPEG5
9Z/w4tASzqBjxM074ue5FHLFTZ7iBQzkqqKrmbZap7BTaWTWUz/LVz1Ey74B65KHT2hGNwjjVq3T
cF34EAfaVhvbs+PTio4JKvNP4UiASXf3pWSOWDrqAMgovn0rRkaxWgLZZ/5GAsNxBKB2VEMj1wpy
yZsukoCwFb6bkG8ksgwiUR9cmbJaHsdnKTAVvNp6LnvMOY+tuwJsprqb2eaGPa1iuHkdKUMo6cxG
uZLCpUxiUJzo8OdTStTFH2Pm6z1Qu5Z3PeLSIq84HBOU8vdkKQsXqa6PIBKw0turaku51LJ4OAIA
KZRBDeMx3Oo4MYFplM9mmtP/evAMQXQn30QGITzWlOU9BTbNm+YXppFdO/8B38rABaWZ6ePL/ppA
bn3xlEQrImYSiSCS7ZzdiavkZqoibFO+87iTKt/ZxiuvVr1sDzLkozVvQoddeNpmXS/4oZi3d3lM
tVSx9QmxLbEd/CgpE/uOo5/gVB+1+BfagWVlE2LVs25V0IEmVDtbrOVJWPE1mFYd5age9dRa8Kcw
wt1A3GM2iXn/nBNniqIKAxoVoww6MRi35XS3gwugMHDAI4fMZ6J5sj8aRBM4WeV17NRjEHelhfyc
bLSZsF3VnZSwlSJpWtnf4Vv60FjQwU3eC8TPLVxJEhZaNPjs5E23uTHh3SzgV84hq6CYDfEEL6Mu
nFLys2m99ZTxCWOGU5aPvgJbQzvphHbTIjs8spHJl601cLWvC448AbZ8H+8ar4bZUFsRxOfRLnlk
4Eqz+YgvMr7V1Vx9/aPhuK7KrmFFPUTDSHfbVL2QwpYIaze/8YFbwUIJBP3XeGJsS0wGWSOaUxKY
SmY9uDnhKg12WvG6JJhAuh6HFDiO0czcWWAY9ey3BqIcUI27UsmRsYCrpOxZe1kIJefProV/44j3
i/dYT4I0R3dC7rTz6jQMgFqujGw+XN9NM0dYddTAIQpjZXQZo1KAGU5F5TZNzP5S/dsTzDH6jze3
j7k5O/BkLVJs8TNODezrXSO5onyFevUvJQ4xwfEdOeKgmsX+y+InrZ5jHePjjDQ52HI+byHQMRCp
aPmWBhtlfjxintJqGJHtdSiE9Fgx7fEyaIVK+I4kmhc5XUv+VEEVsdzUsuDJWmc6hFJAp9pa3i60
hcivKSYIuqlqFi50Nw6BzMPXUm30L3V7S4nKHYBkTkVnQSFo4cab6lsC1NO1m5pRJ1Bv1GNGPn1D
bHigivuyBYu2R1r0j1Rcna/i5oADZvIGhAAv6/AnA9Tfdv1iDW4em/67CXAl8fdr5t/uUkWyichh
MeBs6VpFUrRHeVseYE9flOIPfUbPq8o3fn7ylFDG+oSCbuC7lH5uJajrfPkr6zxJZn7Q+CfLylKh
JnWMFMXCpG1pDthUEyf3du584hJOQ9HhGR9YA4xUzqTZFj+4CRqPTSTNJq2uaTDIcEkLNpvFjRuh
H6GgCaKdvSxdCusYauRV+f6ejyC0+nfFLdh3pxtXguXOgU/FMJw2qa3mc2ee3gVzEJWtT2s2YICE
Tnpl1+QvwzVpqB3DM7EViSwh5PTTsprU6X3WShTtuTj6CTULj4Ki42Vkoqa3SpaemZvvxTUmHJKe
yLVvdb0rkLbsfeYx1r0X/IMfcMb2ii1eWyo2pJrBLxoSHbGaO5Yclk68nuxoZBym+p/Ti85pzTfG
PSR7v9zNSr/D7ESnh4rLZKLx4T1JHdsADEJJ3V3plJeAfLuu8fCfLHBzL5JpQGuF7zYN3MVj6oO3
feECFQrlGdX/t4NdznHGXzMGj/a8m9R/M9f4jXGUy6PYAxCGp/iRagdsr1BuJU3tCV9Wzqf2IRps
ig7Im1Z5KR8ZyCYzysadVbqsmst90+tyJsSWlYwVGYajnII+OHk3MciSD0ENZ0JOGdPcrMzIfgIp
+ybA2tu6v/mmzKp9nLM1YwpGiLBGwW1Frx0QfyakBUZYn3kkXRmUnwLt6ey5UhxcNPYdvxA7TlTz
Ke/nybylliKoJoSzVA6fqVNBnj3R2a/ZxxwOQdk5GT2kLrdr6l2ndTdWKCYRTYRIL3rKoY0lpkDY
Nlnhmu0n9+5dtSPHA1ch8gGsjKy8M5seKmGqqBOI41wjofY/iQKrQ82EgztMwptdDhfNJ6Xfyc3M
aeD8hyhfL3rs/nzGvdZOYK5NVEbAm4a+i4edGnc+FzZCnYv3eJu+y/CikNOm0QUDsHddZOI36gOJ
GpmZJ0XPMr5vO305cZoJqJYSE4lLZQ8A6QA24wBFdXXqe4KdNr4BDPUFCYyo0aM6LAGUSjGZIzsr
RtlTMKStoZ1l8sryUnamQYfWofxhSOxiq/8mo+4dHEb25vd3vLz/6gh3Zdc07mcLYrDlwfSAIbUd
iJr4KA4AULVtUcqotx30rqkCSDAp37D4S1mm9dK4+iPS36sE2OoxRy/RFA7y5mukuJPpPuLhvNij
UQEbsxYiiobnuuIOKnDPC7udrSvUJt4cT4/D3IBkcSwy6jLNvjUiQp8+IJY3+0h9GhKWDY5aaaO5
eR7K79bcVbbBaV32avX3LMRFPy//p4sCnj3txJ3O/KtBfxntg79PcqZIfWejs+jRP89U+AZAc4Vn
rPO15Os+6khue4x3Kzv5gYmhR9SLsj+6+eWUEMN0jearoIuIjQpOayJ7hboatHcmXyE+4O+GHywh
yiWiizt1b9/KhWonONnIqsQ1cHRJbdyDcNP0DH4001EqU/Ri47AKCD0ZOSZE/o7LMKmHrtt4QFYi
s4JwJhrLOF97+70gPS0mPCZhjzQ3Y6WNTlapO+Rdyi1eibVUtknNZh12Lp64FiGRBVOPsUrZrF+J
gKC4ZMuVB4q76z7JRVoERj2LxYV49CgnJ/+CohOazsBv3uWNm1E8/gXiN+g6Ydkf6+GqsL9pAwda
VIWAMsm9+HeIZYcsSzvoOpCTERlR+ta/jjdZNznbBfw1os5O86CT4mQm+2jyRE42Uqv5j1ejWVEH
QA+jp7IWeFZySaCPSgWYIEU9qOlqathKgMPFuaa6GwzbWgtFaQx3UPmVyexEnNJP2yf4XGgXe/Bb
No4hPW2cBdw1djsTmftYMFDR8hch0ikfHbD7Kqt54ipqEci3kVBqokIvWUtlXfWnQY4ztbkCIYCy
UyAG4H1WW2gDeVvaDwp2LOFGOJCEXP7p6/cMtllpTkrURDwxU9lrXNL142nt6gN42dRIeujU1yaK
zbFJuyJ1hUuY9hQ17qhRev8wKdYjuGubkq6zxa7B6eTkcpGO0ppBqMyZOHSOu0/Q3m28C1q5LzfE
QRI42yxv8zk1zuOxuiNGV3ymLcwcQL7SMT0htpx58zN2hqDDzi9Nm0h6wVDMp4T1ir88z4mcP+i4
y4JIRGWlo5Se+/JBHh7xkurJgXMsxqK5jUe5kAKj+kDijBptfCZOtNVzo8jYftcpBO4dMThRvwkU
jByqjqTLaLU4CHOqa2vgLGOeHm7Gmi5IP66DyHvPaD60gH+/7VButnNWYvKwz5QEb2o/09yE5uWS
LtMlIk9eA8UY+lzuPHx8fqvl1Y+4P/3foKKh5S1WZ9IIUE1tAyO6wShtX7+AFYQTTHjDGkPwfX2C
QOxnwcoCXt4rbmZ89H6P0NuOuJ1K7NX9TemPUl8hFwgn1kOtKB60pyL4FEefnBtd3oRC08Gt8gsZ
Yw2Z6ZfkRDn2ubffZk6FSUt6n12MSRVthJIfUdlanELTYcHj7VaIcVEJiZMOBJ35AdQx2wo3JLl/
cg3J+v7mYK+OmJQ0GLLL3tDri5k/eShlLaBkKZjsaufmt+fUrSQ5xYff7ag+omuM3by9k3pSZidi
WQJutEFHOQ+pHM4AQKtMIybp5IuyKg+zmoVnu+569Ao7H+VUKxA8XnztthctWpS3KBdhLq0aub7W
pJU7A+Qngl9+xVbJMdhPscdfkrJbXAPc6k9VuJSrUXJGY0+W36NU3Yjuv4shEapEr/wTruFemkGf
62KK8RsQEFoZls5emlOJJjQzJT14b/pm8BPnHvrSxuas8SY8YRL7XZWO2tuKth1MjT0tUBMerCMZ
VVEWqOUUS5GG3V7+io7Wiw/LMzIkmEwPKWComc2aAA+vWANHeVWkuQMJw03ssAksX2uZ4gm9Bw99
IUGQgFLJ1r8W3bRRMLf1Lmfl1RH2sFGhVpEzGLfPb+na7Foj6LuoPMJ6fzPwQJWHlAN+8jvktFoZ
/OPhUq5oJAl0yai3j+mGuLfptiX2h8qqwK1xjwMghKZGaSIhWD3fBLYQXC5EaOm0codGoXC95czP
fuymBN8qA9Rmma7+CrSwBzcrQ12+1qu6qYfyX/yVfVZbvo5gW3ev/byVqFXg10pDity0jQdnPba7
Buaa2kMYUFGtOZAOmMde0ab696z6+ENbko9dXgpcnJGcxBLahl3IpfP60GsG97izVBuB0XT3A6Fe
asqmJbDzKvrRy1Xj65/4cv3n8h6BU3MI6P8isiohR5mxKjErJm8CAQdaZ2xMsPJcPSh43tZRsdxQ
u/wuePdVKrBfxzadrVkyTzQTTjCxFXYnFWl1GjlYDSxKQOSD+iBzmpE0FwB5LjMe42mbj75cdObR
q6YGJWqWwnI1Wi8gr3CyuCPKyUn997msMSTAgLhnajr2yb4PR/sAg3Ea3FCwvtxgRPyYYZLfXukl
6XBhy1oZ+ofI3sbknH5grsbh3xfHde+DvL9EBr9NAN32Sexd/F1zuQC+zrQsLm1PlAatd5GZ1N5z
omFZPOEN50WEiShmdNb4PfSUhNtc0x4G+VVn0xXr5UJhVuSqjceX/BC8oGGh3ssPtzBWz9J9y3cJ
3i7CtaD/wiMO5MCV0SvihEjYl1DWD68sOKFVGLyjX+qPkOK1m+YZ9NvhbCJL6Y2p6VjZkH/MSBfF
1LXJPpNBS+fsrVx0xHihPr1WSAvR37AyIeO/LFhcarSARpahX+/3/m9y0QxwgDkOt0DLeSZemuUm
1UdfDgvakOwKA9M2QegnHaHWlpFA4rjoEb0GRZHoZ6K/FPixSzSBZwG3qpjGdOBcEeYamSuP9QnN
GUPh0GdudI62l1ea+hUOblJWrSzDQ7qiUlmeoL+KCrQE3iw6TMnhmN0rDLufdcBxd1baV2noY19n
TNFaWSyO8CxGFNgfEzEIKnmZS9vAd3T/ZY/1061bu98zU/KwlkfJLgcpij8UYAXlsxJbuGXqWJn0
wM2HnMeZ8lNiQwvoTg8ycQKsy/ZVUHDBCnPSpksQEGtAai2uFsdXj6XlXnOS3D7Ut3Wu5bU6B+T1
Svm1A2P7xVPVB3wA0n+e6vb3pI0uRzuW9YQNFRgZZJ58aUPqKThz1aiKQI/5Wi6/5XxVqS9/y5Pg
EtP80e765ejKpziJxOvVkEv4voBK5TtaXuuxvttmG6jVC0LnWQZM+93DoXJ+kJHzvpad/OwvcAT8
7QwnVJtJYSe3whbuolFf3JZmU6b0lHL/t1KjIzEBt8wwVUBmNuC9qRv/EBrp8SAL4r21P3q2NlPv
XE/XYjG9qC1MqUJ3pJ9Xc7gk/HMMGMEO358qrKCfI41+PqVJsaCCu28crz4EegD0RI+yiXm35oK7
mT2qefsD4zRb4llvvIvzBOeI76pWwUTNizcURHU6E+piCH4vRJFQA4yo3+YEHPrdP5mGc5gcmz17
kHW4yWqtgRzPx8vbOPY/A1YKI33xEpkg8oBqAs8y5ucaL3r7JEtYqV1YVgtGQOyvEB4A8QnxlKRz
YXxPn4R1wWuA+v/ep4xgL+RZjMR4In23VUOdqX/nRqdxk8fLn9a17JZHyZ3+NE0YtgOQQgeg3+CD
e9DxlMR+WGQK2DwZ1GnkgyyrEq8BWVSAnY0Qf1HJ+d9b5wW4a1z2bhLe2dVMMqLkGeWhh24/K7o1
ue8LuSHz+bv3lBf9hP06zCWdbljzMx357ZUG+B0rv9SBFfWkOLA8ljn5l7nN08mEtQ/4+qhy034d
POGWayoV/Sh0hyrWB4QOyih19UTcxxR3Y2bCbfwA6db0hurCoEVucUYACOSCyaOGtILPkDUIVqgN
ucG8WqbdsfYQsu8q1QZPr2tMoD9FfJyaUcf0zOaB2VeE8mXJoMm7XL1VQM+7C5GqvG69XBm9gVop
xrDmSDlV7mVaOjEqQ9VRXq71X8KB6AKCngEVLSuKuCRTcWUVmue/4jlRbSABHZb/SaTTvJ/VIZFn
+6TAUiubC4+uLEYV/vDJU5HUfWXkpda9dnsg9Xmyvms9+TYxvoQ185Q+gp+PpSy6R9jcMgEss9zn
8FkA+u50MI5/eShwcwBck1yWegq8TE+X3NlcnwxDRna5RgbL6v4anhcr31rcpRUSpPadCCyHXmtP
zYjyPNNZX8Yj1bOuuYS5c1cP6a4I9GkQcuSG4CP6pgqD48ZylNP3piKFXRbciWjYbRYaGHERDSdP
sUTsMuUhi4lKQKmumDEH0uT00OXV6/FauMGovSo613g5OfjN7wpvl7tdLx2Xm+B/A3k7EzYEkEoS
w9LQPLBvMhY0Is/1E6XcmP3Fywna8OCwjzeNSHCbA6WXsog0/BiAr8P8BlniS4hT0vBC7gLJcVMd
y2D7mx7M/XM4bznhqK7bdfNZYnepFSp2Y49RrPGCVOIaj2fQBINZdSAe785/c8Rw3nzEwCEN0XXO
ZJM0IyYWre7/SKS9vbKiB4VvEHLm15YZbeIhNvegjpcvbZCrzJWAS282GVgwJWkp9yxTnlSLLidW
7PmLieOBIbNquQtqz9wmsmVrQuaKDsOobrXQgIHfL8Ku3QBJpKMiAF4SqFzCUiMh7nXqhK8PlOXw
eblPegEZL3HevA4Qjl6w91WwAkeMyz404HBzNrH6hz6RwjyVhsQjw877yxvXDeCglUoyI9g8zVnI
WoYe009C6qgyBc4/llajaRr5XpaG1PVc6goUiG0SGxKUVgVJ1KbM8oFEBWTOwO9UCmV8rzGOKeRL
GKWkrizNZgVJrcMWIE8dUz+E00zkTkEijC5sHl9TfXtuTATV+F+pA4Nkh2cRW2KZGVIvOF6eoDO3
+hATcR49yskthtdcRFTWCxBw4CMebKbXSBgUXjHukcc1A8w2Q/C+swTQjLZh/U15UjBzH/O1NrpM
nuSbb713NvlsumT6jmypv7AcqtHQ7BQ9Q8EgZO1JeqRcRgIIGVjjxJwUikEJFk0NQkT3bwU5rk9b
N/z3N9tRp7uH0dXBHQbP11yH1szNZlF8P+K81rbkgMlOXv43tpJ4z5zGBRSLnVQTPe9FF9F3s10d
CwTN0+a2J1dWbpwUscLvhtFp/J/N6EL+PSs61oLsjEh1R3NHtKwigf35Ba4REwf35Lex0Fj0fDHs
LK5PGWde7AkKdVu4x3DpblZDlWheHKWp7jKCq3Ff7rT3nHBPVZX2QcUwQBx/dvmqOxwn5eXnJtXz
4kXlmDs1poFxGtXPnClaUyoz7r3AE2ogBrry5gDZXF4WWWmsRFIQwT0PSCLMVZjvUuqb60EreASz
Eu0r3mEdn4oGZaiR2ke/ketZlCpWIG+gI8S5oNKQ+qJ0rle2hWd2qYbk224kolD/IHztukbaL0rv
nmebadL0kzKMadmCGrs1mqyOcQqWuq3FGbAbHoCxg9Erxqp9R08d5z4qS76Tu5b2/dXpWwcYVd2u
zEIU8nT+GLLLFHoesl8EGvGFU/730FOXu3/ALxEHUOEOUmEm1LcLVzXTjxWlRewpa5I4djg9qSkp
LZIUch98aph1xJ5qktZAizaUQzSmO6ztETXoygowigZJDDBl0+6tDiFMalfuaju28O/lOdey91oy
VHPrxXpnsEGUZjz3zD8Qh22LFzyj5U9WhW2jJbW4MUsCU0Bzy8/1qxLvo3A6RL3kq3EBo+QLhdom
zvdZjLW/c9OlM8nSQj5+VaGmLIWL73eTFvnNG7oAjk3Eoyt8PnWdf3mZoNqyWyb7hPoR+EqWCpiJ
ruhWRomX+/kbagpBjFN+qbMlZqmNU2qkjFGQgaOhN+jPzTPtFKNI24qFTYOUqtCVHy1/Ijun/DUU
811U9N3PLaG0xPqLx05LVMBqJZKqYqfYfktZnMEx3ibqOzX/LOPR5p/g292Jjq8+P0HAEtfpcVmo
0h59CT1fFMnFkF9ZRLe6akLmgGN9FQhWklLXNR+MAIg8ePEr6fnnyZ5fG8qS6wMYAjFKZbrBEZnO
V5gvlxjZ8iU62KUeDVcGuBfe/9+jM05stbeDQ1PyziHaKsHV166PKqK1E6kPKGjrFI9gRbRdVgPD
XdOJYLSHXJHH6+DrvSboqK3utiy9Jcgy/rSiEfKxnr3o1EDR+8/Y71UGtLJHz1hjQa/lkGxLsBeM
G/mG44YrVKifCdlEjrF26ZeIFoTxK7SEJDGcV1OTC2vY/29B9V3JsONC314e76MLT/e66lcPYJA6
IwBUWzIVHZFjzMZuBZSQMTlQ2NdNa7q1yMfgIcEPy/emckSvpU+VW52KKk7ou4VB5Kt15jHbYU7n
90aozDrjo04mm1g2pZJR95LRk54XdgVS1Jl/ecylJ9ll0BO2VBRlz9LxbrVifeWB4AueXlbF+hM/
nfluHCXTlwMN/MSdiuZIqumG3rB6X2jCKR7iX6CN9nxaY9o58VfVy1xN5f64FX1SCI/pq7ldsr+e
QDG1IhE6rI1DxaTuGrmPo/Vn/X3Ew7AvAfaK1Do7Lf1jP0uXs5C7aREQi1txmiP6gc+fF5hr05AO
Q/6jJyfcgX07uEwlnuKQN4fwQj14iJTLBnwE1pvCqBYo7B4dyVITtgRNZ1YzoV3h9FAKUtQOqOen
jyFLpNnvddDOD0x9PiqCSfnZdAEFFxyQvJ8HT77mAl3NjUoxF9rmjTxIbPoK4Ol8lwfy7SS+2Mco
IXunflmyngbZ7d5D5OQDbbMa8zQ0qt+0s4IZNQRlGuaoqUVjLJFxKhYtBfFBtOwmcjnT8sXbkaMA
ExHAWuCcQMryeuFv+IbVKdhk9gT8nh66EZX3IimpBLxXam99HoPcREtJxLDN/M+dTdjDD0vq4kWz
Wet/9LE/CnOh21e8pn/RXY7pW5ivrEdE3k7x6Pvlh6iTym0wRP/ZKXn13xgi9BKlAfnA1xdX4GQ5
MNRh7ez/JldDz2qcgxwZtuC/wwFFB1qfSNvUjGRd+3Fu1cMYPbO/rXxEkSUqsT6aDBt3a8KS/no2
02jX07JgIyHLjuE2dua7HKWAK/RBKhPsin01Ih5OxuSbzFijZaS55keYlgUHx/H+jCMdz6B/h8na
rPu0oHMSLOeHNKhptgQ9oFqBk0or61DAc/yEH4sWsLJ9rI8haQO6LnCjJ0skJoYiSDx7rY3qiLlZ
BT8X0mOwRZ8ozQfpCxNCvSrPmhQQqWzXEOZry+qf1oTKKQdN3cwGuvtXyMUTMSo6lSqPGsARRhIU
QnogyGz+6WS3DydyAydUrJyHckSMKML+t3qiCP8/MG9CA+momtZqxyHZhBK0OSIG/pjEk1bHXVCS
t07P0iKMFH0RtK5JJAbAko3LNKWyklDf0w6I6Cj4DTEZRb6fWeNgr7RB8QU1eyajwPdzwjmGd+Zi
JexnwbOPdozQEjmREV0yx0V+LD4p4zB3OKFv5ZzZxhvU0Thso5p+k/yBuoUxcPE34xXzgs5RcXD8
bY4qw127Gj/kM6Hd+aDaYIZHWRXcy8RW9EHFfM6rdaYx9WAfCri+zjan4ICd10LWM7pNHmnnui/m
noFq9JivOhtB+ZVCgmYGQ9gLn/YwPVf4zaIgy900CnPjeVLtAdW5ZmAgxbIsIv10+ypPzHIlK9Iy
7k5VL2y+fz8wLicFtHluDPimKFIQ/Qk/CDb1t9mnZ2FHw+OxX9n1GhQFjT+J9tRtIBjcrxEEK1cy
vF14CApwq63Ekg3d7snGNSFpV/GUraUtpbs/5nj+fKgX/X0JL/TJTU9RiFHPulBBeYG4OEUY/bV4
+eFm2ut63tL1yOX7exrpDRrQdbQXvL22uhuRwK9zPBcu8vXirOeZ02wVh0lMDyf7YFCEDlId7i9i
kGsv9AAmCgsqrbl73aG0mxbknMidmZ1cFBpIKJe8p7LlmlQROt1LGymDwroH+C+JKMnMSURfRHSj
FjQ3YQxS7Yyf1zdmtAKEHrQW7kg1P6vz021BkVJSSyMDyt7sOsxf9cUNFWuubfBP2eeQTWwyVR/h
FtVx87DDQnQZXsTwVWqqGshfMl4vSxtEwYfitC/rWQvKbk59oafih/3Y1ASlBnjNKnIToSWDMYay
Yn7emQ8sh6ww5tYMLs1yV0dwL6fxojP0BTt0Q/FxP7Gsbp7fqtx9lPBC1UT5aLegDA/xG5RM1WV7
Cl28N2RH0u0WsMXEOvAmgU4Mvi1VwXx35Y/WeW6K60Uf8PHSCazmAFikPJgfN0Wy8VylGqKbXV0u
kXvQJl5W4MCN6r7nv2ZmMZnVTccgKody/zrH7cN4IGpZGenUXFpjkfG3HGClUEcD1mxmkJWHWoZb
j27wVxlYdF97+aGRCB/xkBRRfL6AVDkYI7vhzqbYXYSo5V09tUldxFuVRtIEIJvo/kvdlBaCM2gk
I52Uj7ztLzidkinT5R462tnjSu2mHFTNLTtAqmam+PxGV2G/aUmXiqCclk9MX1eyd4t7REaNlNPV
/FZz7Q4JRZABhFroSAl4KHymPTcHbpiTJA7scI/eep2j4QH92sHUsKkdJCDFTHnZT5JbAwwPM4F5
7dAsjGPRWJqA5TZyxo1t+/TkdoRXjvPcdaxD7gDBL9vF4h3Rl+AcXQI+TJ1Fqx77cQCBgB4XXyA/
0K4GcRzUuMbcfU+g5H9OH960g5Q69E//vLVnsjSsUUARLBxgEFmHXKJwOBKFGxJXuF8mSyF9EitK
v4yG+AdTQjVkvhWErkO4VmKsceMd5nSqtp1vhA6jYp4Kev94X48W73k0iNfauyKfd7KeWa/bGY/n
FDiyW/Zu9QJLYoHKRwYHZtjloOeZS8rkHx5Cg23Ql8DANsXM4p4mROZ8GvRQHIdyVPOK5tbwoBrl
vQW4A0VZsElqMrTQVYJOLu94BQ7U9JFO5xx5M/VA7HjUNX6HSYQvgEf8UYECHve6bwXZWEKdlZ2v
M/8W4D1M0X0XWAiKM2DEWra6HdCEV1HNWXIkXMEjfRS3qtlaT48VJ7rY6ehx9KeC22Qj6Dzzq4mO
5G0t3o2CPQvY5vCLMLqJOUd+Sdpld1Vj44lGA4ZBGJch7SEZhjC2vwRkEmiyfHHtXDuNbB57mr+K
gkGg4RSksr45xjyxEKIzdCP3ZnNHLDyGbUdd6+qVwGMDTtCvv56gKGUwDBV+rycwgRokscIsUNoa
Ym7ojAYk7wu7r1B04NWd3K6J76wSOUTaVBpZz2qiUtE3LMFUPKrZVyAYCumjHdKKjk1o0nMiNwtR
LksJTeCp3ln6ot7GaDQ0gDCLWQ5cr0TzohxkWSET1KIZFenDsRGTK3+qwIH2Wjw0ZhzZJxfUfL4t
doj5sMPyC9NiztJwgNojW62FCkUfjbrjNidhVAXk1nF0czGMFiqoJQ4jSvqvMOkcpLYqfLivWHzY
98d8P+ynsjP603Wt0YmylbpEnO0mVbscy4zWL7IPeA9Qeo/f8Q5R+Wl+004pFho6Psz1wvtDrAlp
dpCfQJ/yJ0iaOcL2jAP0wtdE+SIYQy+xhVidl8U8YfGThzeTJ7PpoR1Pj1INWr/QEcX5BOuwjXIR
JeW6qRkP1TWtOA9V4/qTrojuq+OaXvCdLZigmgo+OjfBRcXuFPbSoyi148mBH8Wr7P7d96r0RbgE
3opE3e0U5o9pg7BMMrkioQLO8hvGOMs8nEZgQ6V7OgC7mtAVJmO3WYOla1v6dsTDYNLq5rciLuXv
QnQX6Bl+L6gWQXQZAooTAj6Sznlc6vmUBu4JLkuRLBG26mgYhIxx9JoNRgURTkhMMF2IKYRohlxh
rYRVPMJSAPXf32P1k/YQ7mXd3E0RItmlKgosMov/ljKB2/TKuYqI5uW5HZgU0gBqAepmLSx6qicR
1apZuKMU3Ve+bXBC1Yrk+acK7bN59JxWGb/hhzOB+n9CLbDh0q3Uohysfb4v5h+tNPZ1jqOacGUB
kRwsArbzD5LVAxdguwUrFjPRDFR+pJUrSTvZTUz9oSNj8MZ9bEBXheCS2sqthw7Xa9sVAxrCs7nn
kQXdclm33SyE/m3mruPHHtioObHZPlL5b5cAKhGdYTH2rm39EuGmdrf8Hw9YPRnqITIgaZ7Ogsnc
edFH9RXuiLfWJ8/6DAW6E23MahDoDqujvNaT676/GAAaoo0y+PZiw+Rm1aCrvKrOF1wsui9+EVh2
v3zh8X7Y8h21S2kUAgdjQywRTaC8imy5DirQgwEMHC40i/913AkZC200BWl/sUuP2MHA5bXjOtpi
AVuDmHvxc3b26r1M/wMKcATonIZSCJHm5NVlCCzWwN266/7fia4ObfC7kNADZ+GgFBnrHDzJTcog
E8LPY0pdGind2eFoK3UNu7qx6mgN3VLV4W9/FXS1emTp2KGm+A1+vts+lEOGWBnXD3ZwnnUATwMx
cC/xd77+MgsQ3gudLy2RtELQWUtI5mdi/QcQA0Ce0oz2tdrR3sPkKBhsWIsUs3+aPsljj7JxI2cm
BKMSC45MLozPgF42FKcNo2ZAx9ML+2167ZAAy9nOiytgtdyy+XD743PcQlsafv0+oFVI1A32ODl0
DOYGFHtCz5ApOcObrGtBXzXJZ6Y6vRIMKJ9G8MiCtAbKdRadmFAOCa2fCDpWfId8b89GAwHtlOVN
p0Gi5hjkf0kV4yI+KQ+dYf6q0gpja0ZEEF6MSmQBKBMZpGvZAyYP+OS2KQeDYnuYT8LEfDV99ssH
Y3xjJ00Jv7e20j3lGqm0v6UIHvuPsrzeomt2rLrxt0Hmcfh0k3+Nl6a8UQLGzGhww7ps4q9fbvWN
Lcr0DF/nsJfkTzjvy3jivGezJUqK2sGwbpA/L7H+gYt28oYppfJs4gqWyu5hbiwLI5uQSFXfdMLq
9eda2F23PvPuhPkzzPLj1vUODdpIg3a0Jn58FTHqOzPa4/xLBChlfZYVTolzZsc8zZMi8WT7QKzh
uxyyl0yeQi48i8oej60cStqK2DLwJFl/tNnFlyAUEUEPV57Lwh4Mm9FLnYfKA6RpkwC1LrYsH0I5
SHwY/PuMjEPYX+ZhU+daP5iQ7SxeQRugdRqstvniVfCnfeXhfjzAXw8U27kcxLocJkRj4cGUHtQ6
G/bjo6lJLk3Xtvu00scTHse9oyWkfiUoAEIzmIATkFLieJyRoWOKH5WUF1OPv6a3Pr1DsVbdoAki
UbdLXxBsO1uBb1LDNG2C7yoTg+RRuSQjhOz6s+imT9AaW4M+ACkPZTHjY5bH7Qkb61TdS0W80x+q
G1b77Jb2AZsGmpQFH6m3ehR7zV79icxMY2qx4MC/3ukMCHGsJRn1MowEdqWoyrrd1d9rXACG3L8n
ptkEEcruXzYxtZ1lEVzQr4AiOshV4/rue4tdV9elMDKegOGPQnkY7Ew0wA+Gix4lNhS4VpL2jXNV
e1KbNoOFkEMoov1SBp82PXiuVJBSqeKo5rP1+6jeck7NTA3sx+r79EWOpppKhLnFkrEODq+HGvqp
wqMwxZKX7uugNArqgmuwap+KgQt1UI8yBFp7rTxpT6iBLKVCoBF4vb4hp+ysaXtGB5syOUarMUib
8xGViqNHZj52iqHv6cqufAXJtACJQ4yCr67sJlPB9i6J2oGpqhhX0asiVRU7VZvLleN8MBtKIC5N
cnHCSlRJ11iNj6WKvMXNiWadQHuJ4woKLPZH5uC0DQPh2xLIf+Aaqv2wyK8VyS8PbAu1m55JJuLg
umbUBAl6OxFGFxIZa3W4omDV4REZ7VnydcF5rmJZZzCd8xhofwR9ZSxdTnqpXxVJCyW/CUR5eGj4
JMmW41Df8aiHhg0P8OnUIu0uQ99mbXGgvVBrcJ7D8eEyUDJYPj9cUnK5yB/DKg3TguO1YO272oRd
psDu4VpbVBDsZ0djDt5pk3BSf846vqEzfxayaiWrjQdWOvwLG8Imm9NADaYAjnQ/zvFvytj+wFMb
VKuk+z5Ev0wTH3CqAZRa4qLXxP8c7IibM5h9GkzedvX5pjjIm/EIlygsDzDoKiopGl2bZURj/rrx
tqkn6PZAXHn1KbYJilehJDJ4BWGAUyAyf2w75IiMIBQRB0apTVc1m5Y4kW6VRShOcVAcCCD3y9vX
n6zeGZv11EeCQMzTkcIgwt9zguUNf8Jy36Hb8UkJ43PmJP4BLFRgKeiX5eVO0jhiTnyJdgZZ6wv3
K/e39bZGdlEaiZO2L29YdzeFsVVyjOFASxH6lEeJKNX7dAFZSceMU5JHRbyJxEH3oxIWIKMEwjzA
QeZeEq0y9Cncdx1G3OmUelDhpx28oJC71c584GiBpvDnlDs0j3nfZGLdcQr5M7Ne/T2jbyUbmlzv
mlXwqGvxS2VQDomWvIZdtsbHqLYCWed7GlYPo5US3wTawKu1qAo7xo6DNF/KNRe4Z2m3EdtuomZ+
+OXuyX9frB80xmFp+DgbtUa7e6/qluubx26YzwFZKG9PrXKDMyslIvHo6TO/I6GeImH36k+CE3YI
G477UQWro3Y5N76hUDuuHeJdoeyE2uPMrabRlQNm0s76l4CRtt21/apPMdZELgqKXL37F0bDeth8
XSqVOTBN6+WIHg4di9P4MpYM7Vp5bddq+igmuuP+rSp9orBTdU2bHE+AcXOJOS7PmSBNZzIf1rw1
lcaKafR35I8psA6RDa17s/+6xllAKIwIRJDKOF5UuULZMCGzIJDb28Rvp/NXr1Ppa8sgroqhfgYH
P3JewMYjexSRM1zzMZmo9xK/jsW3wguojaBoX6gfrYvxNK+wuyVOjxtyg76RiaVDbimjSj7GQqa9
t104LURaZtIWTWVaCY4Xg0DWdWLdnWaKLudBxgE21qjhgAiEmhmE8zDFoWHnWKO7k9aJm/QttI4d
g5amZmcsxIi0h5esDx41yYl1K24PyE7TI3x6tKZVdMz3/VivoiRmFs5zKHL4FmG17Kv084/7Qb7c
6vMqKcxTBJyjGTAhP97kQB3NfwHvxxb3H7lOfiG7LQp1XOP0Be1D7IwbD9wJr8e2aVIg4vixVQ+N
eDYg4yqZnt6XzqdED0IKNfNUwmfMxbKABt3RgwJw9f9fgv7yII/Ef3EfB/Nh6UFeRn+Z5cFDtBXB
O++6Dh2h+rjD2oBKKjBR9HtdyJdE2gS/eTrsk3w2N57igRwy7EtMYgnv1NFE9jGX934THY0CoFc0
gi2VqRHGIOYr2V89JakI58rgYXI1etSm8aHajKMlSihNsvYdigrGEPdXmdAMY4QR/kz9cNimzjvg
pZtZA83x8BbKdpdGQTggv1s0WnA6nh4FXOUdVrXD1AuR+mWTjCbsrCBRCP79FcmdGr0ekm7f7WAb
DyPz3DwUfIRvytE3iW9voH53/efLnICjGY+h8cv8+Aw9CTL8yMQGoU8s9x8r57c1eUZGckWfHnVl
+U/gzRG9doI705FwzaOqrqhyKbpH9xqiVS4j7FZJlNAfZcoYyZAmaU1sQgT5DLw73fyKlHNO1opI
FoppkLToooA2zTL7ZKmaGOHxXFEY8ysFrO+JT3caCOm27NnGUl/HIqN8uPtKhTq1YxS2pGTrjIF+
/TmshXB6Oi9NOQkC5QyfiCeOlUf0A+W7tKrGEpZWNptpFJQ6ZNvIrKNFc3bPLVavAREB76ONt4PY
TH8ENVvq3f8FAp6jRNMCrCqeI5w1GZEmI62F/zjUV0Vx8TZGc5ohXJUkxlKoeCQ+bH3psPLPO6r9
ni07NU9GPveuUdR78szz80jGka2qVO3/bcLfNR/kLsMfoISfR29Uxuhq5twZ/LFBSTZAxl4P7ewq
21o+TnFUokd1uKjlF0YV+8I1270NHHwTBF6Zez0h/+e1kfnqDjI6sR5kirmPrLKYXy2PMeq6pq6O
/nVwlCZPGWC48yTTpr+fOfsfbMhZJH851uh8pw5jRBpiIFQ1Ib7aafPW5mQknTqxfs+a8Q9l5EsE
CZ8X5o9hJWSaWC1QRqCTKelsj/MaDJxYf8rGVttrPSvenP3C86spfNPZEJt09rP0NN3QbfFDfjnF
8M1hH9SN7F9BXKXVUXoXg/oUEGQScWRv9/FIs3/scKAfW3Nt+eQasaXBPlJowtuqOfXhk/jXJFVk
fuXT9myQD7oAsiefwxbATo48FdySvfPrXqnUtoMV+Blp5mWOq29KS78q3UbrqEImaXhKdpCwSoGn
Z8amQRZGNOMX/UOs8cF/MrpIyzVtN+cyPEhXN1BZ4GYgRVZOkoRHTp2mDSDCJiZUyGZ9priKW0tw
HpQ/urfOtqQXrnEF6SuXaaZRKa3ypdgMmg6Bb6MDhoGTAwwpjoz9c1CR/PC34tdyQ/P9NzCqJCbf
WczwQtJwcrqmx5CqQ88FGOhIBFrokyu9lsolRlMldIOLhmBw8rItZwVleuS5wtC53cfbgXFxYuMK
E5cI2XBcGohOwszTBpzLk4o0jIRpX/vzS2ItTvp/3J2fyR36nneDkS+bBTUYzhuMDE4lnZlR6aTE
l78NG8B+I9dginRJE/2L83HDB3GPPAzcsD6aLQ3JNQNXdADzmnxudv6f9Mahl55p9mRzhVjiVozT
/qRnokOlJ+afS4icCytwp8pSf8eYVeqGtAcw5awulu4veNlvNzCYT1gahJw6u/NLkuEiinyc579n
TcK22lk+/d8cCwPhmb56CzX3447AjqXN9MdK7MJu5+y0/cKbxGO5C23cw6UzDkxEe71V7ZU8G9Ej
xpt6VXnAgIHEBW3QxCR+KKUZKYBFmCJEO9W8EqyvxzCOolvxh3IX/kgRiyYXbUUZvB6/ofbWmn9y
2CUpAapBvZaXu2e6TLGeCHihzB+COIIMJDkydlBACO3nzBNGyIjgUtvWDN98iFArXd1JWJ+ORIfM
mxGcX//Lql02Of7lHX4zJBVUp2ceJqInYCpuxovm7sAQc6jS6rNl1+ldMbr6A9Xz/+/Russ4BOZW
B0y+fmvsjHalciaC4O8oOWi5Lqw3U6encuPv86GBf6WE4kV2kf1+BjegZhkTgr6JixVhRejdfT7h
+If+wnRFfB8peO4pddIkKuGWfIodSEQ7Wct57PgXz4hXhNUR9Gm+hUfkkUD4eThfB15LN6lSLq3U
9zG9ILQ7o8dvFbcfXDrYiS1VrBth08GiJuq8TZDwU4/dQrQDoTvLjKo/QtBZO9rtOkXJTDJdEMGT
n1u1jtHojgfc11KUrEMlE+9YaV4Hvpw4WuGZpM2Kq7EG/zKZMiligGRop5lG2k2QTyWfyv3fBBGk
doVlQC1cLQAmhcuvOCvO3V4Vz9ePPHKjD+A1jcu5nWsG4DWgen9GnCpB3x5nj2rFa2l8t47UgaDD
ssuYt9q832WTi38giDI0ccylDRRfBPGksZaboHNtx5yfIMaNF5KJq5YFmRR/UY4cObyXKvp6pdUR
ceRyy5nvqXwXG/dWIbFdj4jaumBYlOkKn19l2Voknc86Ye3lAOEXx+aVcEtnArJJsRfswKZDc3lq
ldTyWmTZFFiU6FNzlYes3TshRNuY0jmO2bjPXlbi3ZK/AacpqsxEaHHKHOoBtGf29j947FJBQSq7
fLiMJZd81sKa5833U+jh9FuPcge/wJwyOl1yJMI5k6opqYsRw1wtksq+uTBUYNPfPgeuwRjSZWzc
Y0tD5Wh9+NYfOUtqLpuxVQZq5khBbQDjAlp83riXmb3arHRfbJtnv+irwRRLZJ/z0dD2J1ol+Qdx
t1WoYIxrn43ReFY8sfBIFhVJC33zc+kEI4RA5X5b8XzZiivPX7t+gnKu7U0yqpO0GchVocqtPxlK
JR5FFBTSQquVQyI0dwl4BVgHnRKd6DS9GV5dnuxUwRv832MBHjoC3kr4V8QPzokVVkLdd36H/9SV
I8DwqyYrbEXstIUUGeixjK1OOckqOQwf6ciBsFBSHpsc8Nu1zxlPvAYxoxDTAk5M/h77ZPO8jxM/
uho7j4p77hVvGjNwNueP0Lif8TPjFgx738d/KRWbmnkBCGtWoyQf0ijQQsCEb88HuZyYuHlwbZz4
h0+cDRGU9ey+0evVIqPwQtBICZVDMH1Pm7dQQ+0U3kSQLZcXx0NgUHN1h1lcuD91nnwpAVKHdYY5
lAnNPZRQkGdV9tC3ZHmOEXMpjip5Yn8hZzDRiJKSaM4qJg+IAeS3ogRsubuXHSIcUElYZdVOo1JI
damHWtAcKPfqXKCbJu4gHJiLbdsLgRyF69EayHa0lxkndzynbp2hn4YtnC/cnFPsknYWOXWgqPQG
+zRkFVR3ffFXmswCcIoixgwMK5a3yfzZhwtEJIgrzKwcW00s8XWKVHXynfVCTKxleOive8G/hVav
oFQdPBcJp1xcus5NAcXZo8xPiRp4JPFfgtNlFCN+8SoSZfU2fi3GaWbG59vuvjSepv/yQRym/RCC
NRGl1wO9zL2BzltJnGJ3ZwCn1uJnfGPU/xR9RXrx9smnjn0r8l1/H9tPHt7fr9Uub6gkyY4AQ0+e
egb4GKYJj+ZAuJ/iORf9N8rmsHqnxcB+Ke/ockAVR+Gx6m1hJKlh0GPhichUB6q+HGGCc5sIwoUR
1IcPJrcLcwHxy/Xu6CFZ1lkIg6vpRcJUNuHV4iVh6XKQMrmfgwmLbQhEQn7jT/9TTT8EhcI67/s0
1XI/750iVKLYfQkMNomXcUsJgvkQ5EL12Gn9tvCIbMqrEOuvAYocJ+HueHXd18aYfxgW2/CvhZ4D
lym5BwUsk/2Q19gZPkg7nXJ8bhR9+hZ7SYGc1vf599dCNB0ehbVrLW4b80TyACS8w86YHhI4JJRi
jnkzmLi92L69DK6o+hdaUmnhvrvh24IZvUa7J5X72fhdzpgQCKdhddakT/bgnfW1yF7qZ5KqBsD9
XER8RQjdTkgt6O6VwQDkSHWXtw9M5dc9WQVw6EB5V9RAbbyPmU3p0EpVLQLjsmwSs66/W2IBAtHp
GXRTSd88iPju+XEXc04U84Yj4ZrjahhetqvD3UynjbTFPz3ebMO2UDOcMNvmp9symSroGzZTIPVm
ihIxs6J6oqySAb+R8nvGJHafCcJpyIniaKvkziK0QmeA2Ztt+2Sxo+UfXVc094JHbboLpHt5F61M
pc60XSG2CRxqqQ2Nz+zDjSDsM3cqrznUBRb+9HiiRozp1wGMu9iSIQ4BO+DvkQgh11VC8VXGJqAb
7YiZgggLnUCF/XUfZq58p3noChlzVdnyPBG3SzsbxY6G03H0JXNUdFHktNe9vXjw7H3RYtyVYqMT
QhHwdu6GLKOLA6FZ6RJpfhM1o6gj7gE3u2SjNvnf+VQh8foqbJjEwGtGxsu32gbp1d+qWtmmtSUE
r9RWidwOYBHWmWvCEcSNCwc++Fzgbn4kA/J7feJekcxPjwQyshrmUVYxhxT2mJ1ECR2tUXSLoMQw
c6Ty34hfCtUUV8wv6x/ON+NzrHyKfasZ1i3bv07YUK8c32oKjd65ZwLV3muVufK5cehR2w4OqgPB
tUDZCJwnWmkbDH/ssLIKr3k0J9hiptwhzVLrlrsAwPEqt5HGr01nQ+J1tayf1m4s3IpMuRlaplMy
roP/aTJ3EeptsXmgk5Kt9tZ2QXe0cYqwWTFp89yw3yFqWh6k+Vngxfmn6xum+3r3cMRJ/cQDr/6u
M86HAugParW8pF9C6WGnbq5UrRFnFS/TDMb9+WcJJ4UfUVRJTrQA+sK9luKP/yF0t9AW0JVDzOKL
kxSQhZxMfmNTk+3Kk4iOovQd9UI5vOng6J8Gq3+JgYtc+TlpDgDIMSy0lAhPhFuoI7F3eVFGmux5
HRnAU1CkNji/ZeGi0PnvHrXGvuA+GK3r+0J6jTkqAxrZ+UJgaiSGDL7Mfo3m2mnrMapZ0of0xFq/
DBESOFI63jZmIdVAKu7LJi4+xCsulSE2lUAamgs5kYVHUCwEqr5yb3g2qphWka4x9sWDKNkatXqF
u773jxE/gcau9wvah0i15xDZWHkPBV2UW1b6lWbVW8P7Mlp3tR8kp8sEIlbczYhECt2tRP9+yDhh
s27oGnRjzAQ7qDwxwsovk45DwuS9ReHS1fJWoZr1HHoM4v0FXU69hiJWeTJtHfZUJvDXJiwuUssH
MWMvca5GVm5lKXXPQfbGkGhWh2DN/xz7VqtyB9qx6kgEFTIFcT5ktrvDwEYkMasYgr2LwjF8yrNC
tSP452P4dL2FzU8sNIK4qMFy2bhP2nDB0NbS7z/dwe4wY44qVrMwdI2Ccb/tq1YhB0VhdgEmWBJf
98iCtUSHv53vOGVlGTmbt+rKBDwnnVkXpcb6TsIHRy28IaXAjuwb9JY5keeAcLwtg2zRaKw7x7uW
YCjYne1FsrvN8F6Ope7+Lxqd7QpMjyXXiCzHbw7jeKTNtMF8GLqZXbxpE2fpPCusmHs3PNuO+P9s
+zbfVuSH+mhL0TVBvUoq0xF4Co62s3db9saAhn8/FRHnA7D+12VTZZP0stH7qLYh3cmWOxJlU9tK
LEkeCU9LKvFvg0FEZELuyGEeLz5i5AL1eBu9VdOK6Bhu5fCfwMjP68p0FUSWGhiB6uXXry494fva
4zpT++DkEfyH3AGTrgAbwBHJZ2prqLPS5TWUiV3iNs188me2MlrfglEPICg2t0Z3ib4/gnY+JG1A
E9exJSLpX/3jzRJRIIDsYDw6M0BXl/mrn/1DZC4B8GyU6eYNe/7nGsOvxiCfocZNMbUyhOixEn/v
hHrs/YunRkDDeDrHy1BYSiTZOuDhIuq0jLvhEXmBxYLGdZW/sjpQZXQVvWGNtKef3xag6kXlBQNg
m6o2ys++DdmJUNOjGVPdxIdhIYf52b6Q8iJNoQs0dQAOPasnksFsZqiNGx68fSHWDNAhp5O0S3um
ptbDOg+81rV2Bj4hKLhvJDoPJzPFEmjfgaLOJ7X2R30UMFjTxW5V9xVva6f/YqrePW9fUw+lJi2s
jG+9x4c4lJ+mlLOahWXRLPWgQAbTJRCFLc0sep+UXUIIKfVXg/C/9g2S9roPcDViWkP7KveXcb9e
gOjk8KusfBE0fbi428KA9OM6Dxop75icOGkh/+QEwSTp9xIJzQd2FpdGWpPyAFzVWAN70kH/E7rf
gten7vPwGvnbeFUOSc6pG8kj/nb4ZVejGSLYGRmsYulXQceFhukfNgGY0zmh0vNi8uDHWQpGNTMW
RsjMGxbGS7M+WM0sWOEj2CAtqSKUk4ZZbuDkYRX+hgJ/J6VQEyxmAUxSriZbDm4+8vSPhzydU73K
B7hY+pW5EBHMoBaoXzR178+E3R2DvPY/+j3Sb0mi09MEqWF5zkcyaAIYHALOEC4H6BbXiH807+U9
zStYqvjHTrX/NNor24Hx1F4YBSjUD2d0ZEb/zOZqVbbEB48VbxAuYB//v9erfPdgpJRCf1cODeIA
iy7SAwLXcOva9awJn8ivFYlWLgsD4F5hR66xG1jcjvD/8Sr27irYQGEQ8wuo7fe6Q4c/ZipwhlJs
hmvqIQzIsOaWjE+VpPwNscmCb57D2yyCs92C0VimpO9zRIG0eFQH/JMyUYaHtrGNQIVejw8e5ieF
qYVPKsIKHkEhNxEw6QPJijuq1hXss9v+Ukt+5/Y3/+BxiI40EjUmpR+Wdca/7HJg5ehNmOwaSBiV
apbY7t6phTfgee2xahqQvwSnkv6Y7LKfRjikdymaGVPM/OjOrKVn+fXP1N/KHLdl3s8hXlSHzSEU
XCZd6Ca+9stYaXv1bpnUqqr29FBc/9f/Jv3pYfjdOMQ4obQzjXERq/hvDQ6bBqy+DrojWwD7UQ+y
yIFCKZk+sMqCxD4UiSwSuG3uiOos7CLdn1nTUO8aItpfrP4mGT+aFo6aM4FVgl1f2ZazRbYCpVQm
pZeR3Z/UTUcTt3DvQIATjsQ9EjHPD35j9rANvPvGoUow20bKsklrqIP4NHT1v8Ptb9y/alImbiS8
DF/X0YzUeK/RYHnj7k0gUFFe2EG3FQvxwYNk1Lxpx0/W4tmhFxOfhWL0lZExmHX3z57Tpxs/sV4i
qhQ6KgdG1+rdHPPaMZYxZR8MPVR+xuo9vIxVhP5zvmCNh7Orv4a3W9Lwab29I++xd/XCPWqgVoxv
PnbSH7xfqy1Hx5XdfjDtRGCzRmGFfVdjHwdoq2zKeKoYysyvPjYvJjbLbK+OK5nxua0VmdbkfWbN
+YyZLtdhL7AUvOw9Ozg60japks9r0nmLpUl0WjtwP2OwoaJ57TkWN5NRpuWFeYUk5ZHUu63otwiJ
+PXV7cI152d+WqJEi47UubbzUvrHlMjaITCIc4sXft5QjFvY0qKUkb4d/fXZIubDnTkufR4TfnYq
fdNZzt9FrLIPwcNTj3B9SUHIg9CalBOTxrhEsXfs/K0lvGMzEF44EADhn1xIPfrmEldeCLKFv2nW
A1izBLWijDZ0XQmCvAbxpvHAJgjv6ClXBYmFxhR256YS6IcfNar5iDohtkkTGP/VbruqJfOOuuw0
SbGKLSsnA45el7djmNXsaN9Fmabob9PZ3eDrYsuvIB8AST8XNcP4NckYIT/kn4dC/hCHOUpqdh9m
kezz73y4oE3UUTjOG433m7cPgmaSHwdNgiud0eykzI0IVcK1Ku8tG1ueAB6hMo1BEjq1qxPrZbGr
lwfZAYg/oHFkqW1BHa7awansiSx+GkA2LEUUcdWeNnMpPBsi72tjLpFP0U2/bXKTy3cw4NVPoCmR
LORXF7W3OV8RBvKPRl//EAaHy2jg/T7WeiZV+04dMGYWviyimRMQXSd2OPs63bX03JYupChrtpxw
T09I0kp0qhSOfAo2nRX2qcI/m0s4pz9LECTd536lcrItoVLXLVHUbGtFqlVPPziaPyTAKLPitD7o
SBRuWjl3ekLhgonsf/FJwqJx/SbMONj54Jw/aarQGiWmwkNU+vxPvknGjCYg9qYHOpSpmkCee4UC
dwtIDqUBIQSDj5zmguUS4536GVtR7RzyaM76JlCV9yRW+m1yz+uzE6TG0yNL9mqllxjUG5xrv5Zz
dSO7beoK2MyLZSTrKcnvZfm2CT+nSja64ApYsDZUP7nMmO3D2MSt8NyVIJXgw3Jgc4wDj6AVzpXZ
wwoUP9hRD100kTKRDlvG44mSthBkLOl+ZsID76rxJopBbq9X/9DymljlePxLTCVy9KPEUW8Cy2kj
FtodCD3vrSOUTyelmPZlh49uB5jhH0IyTNkHsbDuTJU5vTjbOGMEWxGK5AKXQkPduHSOuXLmiI+k
zzRJbLUWb8QJVwCMG63Xei9qblP3e8KewPxoW6+SachH7FDT7hYKNHKxRG8Ta17IpQ2eg0f4NhAq
NFni7OvA7bz9WTVc73DC6bNKUxb7j/r4NqF1lYznjjCEUId+hrBfovKOfKvi7M2db9SpFAGZAiwf
pVE5/tDGKXj95a1G80vWhOaDKwLap/0Jjr8s1+kaeXnACPqZZpUTufy7HYQ2x3NsD6UMP5TzFYxj
5MHgQMx/04E36ylwv5lvPgZw/E6uFvWe/iVxhC+NoEg9QZmRx92oaFa1y2yj9TYMpjXqpW/4YgKi
vyHIh9pztXoVlXD3lCAL5mOOhaeCjnBJdP1Cs0b+2Z15vq2we1qfFTUU4K0pA1+b01w2CHUEZi5V
0wA14Qxc6eRKRlddZGeard7IJ6hwKZLVkfYiIJ/XMR8YqL/POGwlhmMr7b0df8N+FSSCx9j3plRR
b7nP6vxFR5Z5D9518dSGjKxMJnP2dZFqRiS8qXrNrvQOoCIvKq/0KwqwQxAoq5mFslYA4Tl5n3hQ
Qh6dxwitoouFuCmfCVG6FEelSCBxVTox7WHL3ugyjoqMtlNL6MOx+Py3Bnmxqiyme6y0PDkwtw5H
kgnby3jdOtRVleeY6Sln42CPlcMlyihfYtJBs+69QZiZ2yImnlJaVPbLgbApvmkSB+eeVHr74Mjn
eLaXVFc39PjfXAu9i01QH4DF0OTDBB79YLuA/lUB7JbtmyOYbvHNx5Ouv1XaV1W1RO3rqJg5qaEZ
HjeYjIIvq0yB1sFkRmPB/0emxIrnIMuq1loAG+TKQl+YyUEKTm6HJCiLd6qPVKeXv75k6O3gMbPh
VOEpu1YeK1F53MD57n2z3ELKl/amMf4xY/dFktnjbnquhlevQ5x1c0Ja9J3BkZ6jg8+M76YDNG3m
jwk19QoHshqfOpq3V6Oqo+GR3/OlrlO6KYNVbsdkR0OsBYO/owME+BomqAscJcQslwrF1aWDYp+k
SM31sVPxMzKN1AMNjsHQZG75DfIWe68ZHuiHWoBCZkhPBIP2T4OHFxNXGBaRLZMNguKmMlvbff7C
88I12dWhxNIKOQFvDOnP8teOAJNbyt5kFQNXeeZOWtOImK742A95klmx2pTUbwxHPGHVKGsNEUis
TO+/F5WTwZkhPqSInTtgocf/rO0mST9duEB5otTFkvXbVsPbr4WEFQZzm5kvTcferTXuTWHFFBE+
BOI4pG0pggutChPy7xhsrQVEM5l8pxbxuYmxTYPWeNfQwWF5nxvUX9ujjXeTL0eGoxaFVsU9nXay
su64QTURe0LkZ1POYPV9Dd7ge2s+8yzccKo4XDAk5q8Fl5tlCjHT4xlGBhAnzkbp+ohm1KPaB43C
hXGydptg8xzs90UNeP7FYJYM+GPoAIbtNdh6DMWXiSHbyEDYLa00cq/J6Q0ApZxM0fLg8q62Ubgq
gH0ox8Jqoj28Y7+RDjwIYs7KdyrpOnscShHbZI0lqPrYpEet2hjU28T29SU65d/K6NmmClW5NgBu
4EKt01ccJsy90NptIJOjDuhyuOtNrZclV5em+PeBV8z7TEt1FzFnjELKu48LFfrvk8ybKaU30pRD
JVmcJ0dKRa9wobGbkgXx7Ae6LsBP+pNEVikatyvnhclBfWzbeG898EuhmigEDUVTN+GcXYmAPihh
WLVcdkKj7MkgAWJ6xXsztbxPwmlcnxGorNkPWpYKO9NBdpFagWcbYf/zN77QO0aNDkcfN4e6BQsh
NklxLtqpYxFKRnG4mAlxyRTqRoJmIOkMqZRcYOaKkL9l8JvlcJAQ8ll8kiIycSaqGvUmoFWaEGj6
Xp0eaODlzdGq0SvjWHJzIwXCps3F/EI4/aT2Rq5AED752tPDqDgiepnbbTubiDauPOr5/QEhgIz8
C/g2cIHDqDZnt5WOszxumeQjjlt+tF8Xk7BC2u0kmOy7hZDe8H/sZ6kAZogsee9LCc15iJWS9SmD
eX7um4d/jxuvKsRwovSDmMLsBCLKmZfHf5vSI/H7FODqjsy5paIGIHMIqPZRasdLvH4Vv82MyuM2
tnK5Ea24N19am24165ehAQUq2YRAtcDiNsnYCY4vmf52UQwGM3vaNSnX/ItsEpU2zvJ6g1Ki7TVq
W7PcITH/TCSfwLc4zMPBnQeR7Ly5ud9WUdZi2QHjEBkXs6Yqz3p7zIjoP3nLz1B4acbe2gpAd32V
+xXhl7RWbnkTenCDkyREHFirbdzY4jht8igIvLm+jw80WHmPVMP3LDTFUg74eQMKlY7vlO4YktE7
d7iiPeyT3YscANBGylCrBB8r9AcrwhlXB1M9OAQzK724eyRfll5JcQN36Gt8MAMXHjkQ+O+KcBF0
+SqQYjWgS6Tjc+mwp3OC85VUSdEOWPVFD0FUOmsbLXGuis4aNeG11FNeZXX0hymMeGijlw+J1Eek
Y932Z17zd+yCTNoMzF69sX8xwVOCX0rhHFirdduU8W9f1ppZ3D3Ba2oIpBSUwhirstIfY3nLb03q
HmzJhgusEzGgdhKTuzi7MIdcenb2cLVmJr1nl30K2yngsZY4ToNkA30F2kSsZCZm6x5jw4YYdtkI
hz5h9G0XiPd+zP/mpcYPcDn5/SRxLqojItE4ogu99SgXnuAwKdtVTJ0AOou7IYVDA0Vt/QOablal
SwIGZsT7hUmUWJL6psQ0yRaeizpyIMlwlce9HuPh857QEOE+TtciLPSdL0gHzw5+3xll7OOSrnpR
tj5nJagg8Sefj7n7g/V/opPHTodq5J0zATULG1MfqxCpcJYVJ+ZosjmL8iIXigQD5mZWlmLK3zvS
BRPEFGCauahfVUnO8c5iK7bPNyo7oRITiaT35ELoo0CnCEwTklI8PMWfrg5dj2IsBA6uV8EmH8E3
zkDuAwtJC9PTJXpx6pZxvxaCMLF8ftVzbMa4U1iFbbDqf5GxE9+s42ltQDgm7QVrSh7aL6QNUMfQ
OI+QdITw4GoTyCiEMWd6WheLeDVEiuJE6jMSBW8MXfjlHvAbo2R36cUYOrICnVFLCtPWtVLP9SMF
NzNnE9muFT1ZIp5tStPr2ioLS32NP5VgIISPc9zWmwgymOoPq8DiEQDV0mSG7uALBobR7Y5mSN19
01Mo9reV1By5XpNPMf2I08jLVkXclmXu3i/6n9050Tqm8HUJNd4jlTpUXqF2NjH7p+AlB6iOsFyB
W6OpTPZVa64+BTYwFUR7lgGA902PLb/Z9iFvTVeczqtZ7Loawy4QxipBjR97wsm8hSZR+C1CMVEC
E1fc06CeYaWAWtHwA5FALPUsY+JDzuQ+/zsNSZvzLiON6g+tDibIqwVvrcRoKA91CIhw1zkpl4O6
AeURCTEvNTvpmCJgWD2e4nlpYEZbc/O4mayudVlO2Gkte62QcBsPHLRT7zqzyGV4y6GlOm0uSz+W
9Zb6OeRCU2kFTTjL/TqAODmsURL2IOhkj21UFA9Zh08CPLGL39+OCwLJqWqd0EFEDr90WTnsTRvQ
HGQ/b5UrCy5DSdE1JzlhL3NQRyCabQxwPpDi2HVVkCPfYemspDoxVZIxz09+cBPHIfbhs+op0xk+
tuCOx3DF4J+PsHPEChtqhdbvliNFfj1HRsuv9PReI1dPxUcHbkJ+tT86/gDGQ4G2sveiSMQ4xSaH
Ynrx2EKDaJiAPn3Qzybh9NSTdVP8XTC+EgXTmhQiTs7YRlfBj5AOVd9I/OyV2+bRy91V0wApdC/b
DtAKZbNW6D4UXrDzy36A718K7b8i7g+u/LxpAaiLvF+IXGHq7whLF4sqkIQrfh6Ihb7lZYVohrGV
Kv91zqtzcYQZg1IKqLLBdT7pOBUcbKdUl4CigI2Kg2Fc5ofeD2yatd/7phNVGOPsP39kSjWv1ORT
xAvDT4LWovbd8G1VNjHeWkPCl6wr1YB9S/5cbif/AkL3qtH+z90ETMbayoIbYPbV9bYkesrOnk3V
wkzDO+2kKfjCNQmV48el2HvZLe/ilx9g9jI1fK+tk7eJOb7FkECwfDpr2FU7ffIMBIAUOp62IOnz
9G3lWTaabjB4zIqk19DgvYvueA2wQ14D1C93h/ER8ZPUOVC/Xe7scUZi+7DYvJnJKhpU45707Kst
BLh7aEzTjHUlIezi/TCi6e6hE+1KtJ0juZwf0bl8pojCScyOncrEhbkgol9RFsjtuoFmeGZQ5Cro
EdDWOQSK9N6oP78dAGb0zaIUeA0e+bc10bqIiJL0Uumzj1hXGN5hFCX8CfdgVXuF1iJdb5ltSVb2
AGS70rQQpGWd9dnsywAOdDODhWDjKt9b2dyL/gWFiOkEM3yp2eTZfUFwuzxRMcSpkT1SkllnkP2v
ToGWVhtl1L5a57L8KWdZqXpHazrn2FJtmkQD+4C3s6NXusbYnOcUgFtOeuLx7fE291Fzj77YWkSo
dnWgL+Qkugrvpg98B14R7HN3guHs0mGXy+cwntmi3jWAafev0KU4Wh2tNYqECvnd/VTEsr3Ah9cz
fmF46TiO8/MCZLY3SOu3qSueAJ6Fj2795LaOYi9XSsZ87effinPge905lGo0ldttFz+gxQgHVW9e
W+J3TXs+uYNL3E9/gk+GsSUWMGwMZqzjG07dh+Zw+ZFZUQ0LU8+k4CgOIu5T54U7iP4LwNkMoGv4
VQcV42w/D0xa9ZX3Oj2R8BE/73vQbvAM4Eo+kh0b1/LjVvJUaGqT4yD/62Xf5sMJu/tjXbc5dQxP
ynExCJsT5TmdYuv5x4J5VEnyXHijZlPnvJTg1+upVRZzzR90vVaCeI87ishZ1EhsEuVqUV8h/rqp
5hFoAkL2r8HgcckkomG7laGK4A8ADsO6E48tRLffA2wXWcrLL8hdwGrga0XiwLr/JhCc9Pjd0YNb
UDo1QrEXOkLtMRdcKMP+yGa7VfOLiN7y27HFlNuE4pMWwrQ4yQRZ95XBOTs0M0QWGUkydwFOakZ2
/CphetTITiVqeeL4Lc1iH5DZu1KjR2OnjRqn4LHWEci8Y4mfXGzUNcAMEcyfblWVXglw7iTfUr6t
QbDSozIqy90yKk0aKeDwdWCxsYDPtdoS3XWHv/yWa2681IFM46jd0Jr/d3OOp4bsMoM5WcdgRIKx
IrsLA7jtrw9Sv63wLGTq31FRhjLtGk9V9zFxiTMkoIPF3NmOuF9a02YIleopaJf93NseKYUbaBM0
kBMnBORfrDUcoXQVcRlob933nYlkpZycFG9fgnUC/qqvT8pdRWLAuVP24kKxdhd4ZciXW/f/wafX
TJnX8gogp9cZjKKa3uu2+147crKdqPtpY4A44QLGgiAkR+c4C4u3VNJxoBulh2kCG1cjaAHz4oBp
yiI8LQ0HmFM6sc/h24mslM0MNJGcPHFOxDZEb/Fr4VL8bVLedaGNEKiLaWFzkNs7+qiduel/1N9k
oz2uoebwuCjUDtCSuIQHgleUIuHDUoLV/sN0+yLWFzcP5UBAyXzWehff3faAypmyD0gTUO3waHZB
Dd6V6FZjqMZJFx/AFWByQKxp5rtO0cVHAFL7eyTMnHXBGVjqTVexB4/3YUIuyUy9Bv9Rd/kACQz8
pcxzXt9NTyk5w5rGCXWAj1nd/5idNJUCm4e4YVnTagY7gNY6b+MHMkjXVIOu33ApI45VyotrbI7Y
lGcifIQpNeudR+58Ahac+y+A5krglT4fTegIO0Cqv4DHCyMitg3P8ylh1tRw8/aVS2Qlfwu1ifRu
ZYZjO1un7arRZsoqvV3iVJR3hY+Dy4VOYTQuvFwnX2+SZAv+Bml4NUSMCsFzKCJuP5dZFT+QQbze
UMiVoTMq0QNSVivN41g08TeCsUQ/l/Qn0l3WqOYDbB5ALy78OS/vcr/s6V42JzqdBwd+1En8g+Sz
+WtP9RL7eP1YCYIH97JoO9ve4qdtrRRBByXXtlMJFwithp65iXdwoB4Kwl77O34Lba6dXuBcN616
4TvHEc73sKIZh8fNy3DLLnIQToZLgNcFfcXyKh/X+0huwPqNuB8EgRTxGUM8gUV+7xirlAa/O+0j
26soQ9Z7eecf6lofsNy/QveXf2T/+Sf9Kea1TvKKzG2fCXc/GvjXteQ6pqQ+AeDFe3TU1KnzEheW
X7kSEGeN/WBxMRuzMy8h02E1ifUjBhIHqAYWCfSJKXHmKRSQJPkNlKiV6YIfIl4JlqBEFdndKTmk
yeGTpUbIKWTn0nWFjyOAr5xAr9o47hYfSoOqwikLaOx8iGPDKU1JPNoXrsn84hvB5Hpoom2zvNOk
n61oe7AmoLYrl6NTNqqO/6flmtWJ2Rp999cLszp3krBRiM9hRcwGnSo3UsYLew79KcOAvlJzbb9v
jcwryQV8Birby5loHDoyawho8xXdq2DKbtxBvGHrx+6L3FEu+eYvvUoaVPHPKCeUDtXrY08DsV7A
WzG0sRKUXXYFfyPaVVNXud+veudB+3ywovRZgwaZUEc66vakJGBS3iHruZybTopW2X2kaj4/9bUL
bKDSNrhzQRhgqb87SKOap5v6EQgeNH/mhujDg8CyuMegj9LZAbuRkkyhW7kzzU03RFjIaJfYBYct
ImhQ7vPMKHMsBea4JqXx8BHspcHeXK8BkRrNW6LiUkHObSGVHHtF6PRiUqWTy25lkglDV7mIb+VH
suP+YMggncuqW6ZZjAWOhj8YfsGGFX/e6h3te8lZtaxnm/fqKl1TOfoAI74qQIZhFzaq7qRlJMH9
zIwcy5LtJidND4vM6ie3vV0nAPp1eZxGE61e1EKrFTjJMHyN9pQGyJVStJhUMCGF8Uk3CSOPamtb
Qs2Upq5FGZEYsfAmRbGG6K7MvmmFR9jIgiHr5J3VMpXO5FDYeIPGx5GVLEAvpCglmKuiPxJ3giC7
0myp9EdFNmU7Hcgz3USuzhXmJhp50t62YsRLz5ev98J+qbNoYn3A0l0ZVq2JOZqU+nYmVx+LVRlV
Xt0WEB5EOJnX4L14EEO5Ruagw/XmGu5tqha40SN5uYsVbWqz+zpjc7skvzrSnwmjxs+RlNXyLe71
b6bjhr6m8CSG1pc5UQhA6ZBAHkR+gW5eHsRd2rkJd9+j/S9/NiDHtQaeSqjbi9vWDdvXJGCnMnvJ
9ZXxwhKJtK/FZtM8+nzhoQdgar+QTGujhOYCiAMQiKXw77T9t7PeOUHQNQ7mMZDn1EHJylv517rb
PNkpnf0tOidlw6MBoLBJ+tZcn7KZMb8+2BxPZsm7baAx/BICy7qhyRUC2CeWbSALl/01GreSFcMC
pTP+1OYD5AMRQb6/TLERRr8XOCjQyQJbxTCJzFOS9/5/6BtcDWOqjDumqYt9IubZbLd5g0L+kih8
k8fdiiG48RAsM5mMyhDPZBSiKPjdEt5drV3BD7qlhn36cGNQnYed4TjGJ2I8dem/kW1gHHU4Pp7S
SAJmAbaqV+/JG4DdZIyIHK22Yg8AyAhUGrt2YlJU1PjGo5g8D0X4cj73RI4BS4BSvSwU/A7Rqsbm
YnTVbO5voqVfO3gpnYahlwkTKK/LU9mFbxNys4X02UVuOQ4/h7ATEBGYizrvvZxtxLvxWXGk0pt4
iDclJHh6F/A2SMNr3ua6CnmNJ7bQzjjPJvInisGa8aODEzsx8ddZCkJe53WkBoXgS1vuGMMAoVSL
eKNvE9OXLMGIJH7H3T0dMPfi6zjz2NXfy/nmv+YFkE4q960aLkbxSI3hDKsWwdbRV80P2DEMgk3F
yRg9NpO2qK4x2nXtsBThxRr/0+nMLv8mAhPAJIUR0OCBz9ZjM9JmU5hl//CqTOcfWKV1mZuvZLZU
YhbZ/vautwSVDq+Ga8o7GvsdzbPZPl/JWAs5e9UOBOyBYyXBgh0/t1Ja9gPVx7rUgYz2UAM0az7d
YvRYF21Icw/eTsGqwOr5Clbw8COnK3R4QdSAfyYqlRtADnuhZe6hx7qBruEIxwxV439YgXV1d+IA
mT/UoqYJ6L3FTusP4ayjWIA6YMpX8Ix5di/yQ4A4cAmjqkSv7UXmeN2dAN5BBLtSEmCVa8osRTuk
xOFtwmXhCxtUV88M61/jAvFsMSPHskqeqLojJWPowXaWiGvxNiptcdXTKZBAU27vYBZHL3cS3OTF
PmzEKlo62v3L9GVKUgTTnRIiuNtx+3ikHL2oyBAsQd90c0z62wrjhgEGe/xHa13jXQdt03OF8PDd
Rey02Nighf44juuFCsC879hpcy1OlXZsw3dD3YfMKb7a+6Bk0srh7GNabp+tY722nks8U7S+ZCKK
V8rWoA3xAoNzqYrrWVoxC0HeyHqX0CQm3rOCLgPTJmo6ga8l+Ct0i+zIVx6linK5lIpAzpiyehVu
ZesgoLCsBklzT8N0PN8YdN8YghqrDrjhwVTxUlHpPdpyJE+B4i8Wvr6f21YzA8ifOLWpOnJm6zyh
ISmi97eL8tBLPSihVDwVFQQ4O8cZPCZvnEdJOjsDZgDBKesLqKByVrA3pQFpB4LA1l9y+FQM4yvc
XF42M0ev5sj1Tw4rWuJvwpA0nC9lfkm4pIUQt3t1WEZzNI0gcl18oDWsH6xG9BsKOAuVrmYTdQZj
7DFfrenOaqBK8L8QiapIDSEwMc1MmOpG8/TwX2170Jrc2ZjFWWTfC5xjOUYP+2IIsCdtfhzRS2Mb
AIdwzk2dA5u5tdv3L4/sNaeMVZD8cihnp2VKd0JOgMbaPE5GFDqeRiuTrAsU5UytD16tF9uSC5g+
em0EEVXvVs0CA7yEwu3RkWU7rus8c2nWuSdn2BdmfWE7B5QIJ7TQ1SM6ricKU7LDUsBUWegh7/hN
QBG7RGYdNJrpsWWdSZXsUyxarqTHXc0gjcMdBptxOesytSTxkywButYHP3HiLBNW1RkmNNRtNnM7
6XLjL9SO1bl/grtDHGvDbe+2baInYWXWw+MWWGQ6+gjNarVT9UX6Uxn9WFbVNWpB8K9qQNGQYyvj
nmc1M9nORaf10yBpi6Kc356b2cvMGNrYAFg0pecaOQKM73DPpMy/sacqv0IXx7fopXQjDInWGMV6
8JLmeNfol2zNjtrVdMA0X2QHN51Ifi9bp7iyTYmvz9fJ50bWli8YUcZHzyy3LOqCRAlef+Md7Nrt
3nLSZXYE4E33mND0tPgsPgW8DpXml/KAbMAe+N0kRjayovnp0Nx/Y1btQgnpGaqf9QUXb13Bbzp9
vgCQx7NP7h7n0n0lGCot+YBXzZOBqnuoviuOtMkWqAQY3kGdfNx5XtSQMt2ys+HqnNmr7tZPgJS2
JgfYyJQ/Q5jKwYO7NzX/WaWw5wCW0SY2UTS8ZFQRForIQOsgN3FUwsqS+N40G2B51tL7QmrNkZ4p
tJ4Ta8IbiawxeUB3tKZc1VcMMBeIz0ALMZlVNH+tPo23XRkPQcgKR0lZqiARdr1z+EXhbwfGztXo
qSKJ2u/C3y+gXeDGWt8RW5FVM+JqIlbjOdxYmphmf8+UpxuqcB4utfqaYbbuNs4uvoikf3xgY6V2
gWfxzElDAHSL80isYkEZWONk/i2QsStAukXjkEyIYIFBr5ZUFS8WqS+hu6UI0UV4VXzeZYondYez
Ph2U3UItw0zt8QX7u0ZzpSg67j6qELd5zY4uRft1Wr7dr9bbunOFnaJ2OIAk+AgT2u+oEjhCbhRM
QG1PnRYsuOzQQcntTKTDLBh5C/NSSyk6Yikya8FoFhasjCFCInJpG7Vvy+eNOFMkGnwUw8iH855T
Rh4EOzZCL03jWVgQo2NQrxFx6uClf4viXLN8WLEEijc9nU3wHJ7V8co7j5VeKMn6VvMHeLKPuvzz
ZSoZWBMWXSdD3p/tFR8NwasSiL26nO5wERrp0zlx5oztsayg9w1YoB94h2N5A0tJsYiz5QrUUf2S
/zaybkDQ5tTM8ZJCVg+H4xCSKIQYrwY2M53UCjT+VvhbXFSW2M+kW+zzsBfV4G5+PwAnNVZFrRWp
y94D0vdQIeLQufskEFNF3J3saYNHKDZsxx19c24gPtmBrIDNDfOFpU3pPCno94y273fLfHxyjn2P
thWLdlhJAQN8pFHLjnno5vxEJWPJhUMCHO4Wz3RhFBGfOsXpnoQdAOcXtBFZv6HnrKyci+uy+hOK
WsYWH/owiaAkp1Ts1DZ3EipiTEfj1v3EP1NiJXSo6Lm7N9vJywV2cDq4b4C2Buh3HgownFlcO2lN
GuWRkk0vUsfoNbahqikDJDXUs8KA8tZOhUqLazQ/qvQuvKzio4xnHg1NiVuuTTt4fJmN/XZXugok
9IkKHeAdyVheL9HNvJ5XiSLu38XM/BKuuXl23mPGQl/ZKjIDLGUI47Zkw7Fw+WwtTkr2+Gh7ZNua
zNG7uOVGNiPUj3w4PGWs5MgTGG92/7sKZY5yF7dilwk3ZucEXg5tDO2CSzutuVqL0PdAf6wSlf9X
3WHpAEfID4oQ1J55F7+LkzbtwySnKEi7j0Um5rvrlW6A2A6JB2RLlyCbJmczgTOAn0vtpivQY4In
NyelPgj3k2mF/s3C3LzD0NfWekwalQcH8NeY3effyu3h9UyLWPxHvpfzGr0EZPeUZM5OPWpByZ56
PASn6s/eOvraVcwxLgRkWz3JdBMpPGEXJlb2SzHAyIkJHLSDrLT4Z5pfxiSAtlyQbwlMUEg+MWJl
5XiRcN8Ld9ORM1mA9HI81k55Yxdze1cxQkL76G2TXq6X86kjFpkZcNlCwI3S+pBrKsu8qNW6LuxF
ZROTBXsk2QStJ+mhANgSDWq2B0WRe+hBlMabrsseiuvEQGq2hdHj8aldiyUTcW9EYUoLhjm1Imqs
CtVoy5tfjs5F1CNreyW3BH51P/l21612ktl+SRRNfl1zlqlwzj9tOvwqSSSxGCQ4s/irbSYTbkdy
i/w9xeYrcImH6Z8GUhc2EZwZTSV52wpYbsaIvCIDwaAmeJzIcJwrmicFCf/evMfKlOckrr7ijRYU
niMahsAXmZAUw2uLMzFJEX3/Y1mT0PvFZ/aEEmFThcVJmampdXZO0M2sAK6WpAHPZVkIgAUiP5zN
BYHCXP+Ibao0bYIe/+/0pj2RSHM8vvIQ4qXCXn5y2TNRppE1ab8plP+BanevGpKZIVSdT0v7vQSA
duGkQx8M5+btQxfdq4mCaboH1trfe2bM0MwjCooWaorohvuJWxKTnrSBJyOTwuI0pfpi4tqJjOj+
Br0AKjWD6EeT25Hcz72fvXHZ4uAZtknFOb4ufyCArHOfjlTSf5adIFd4trp1Ai5oBC+ImffKFUIa
khcPd2rbFTdZNCkGIMaVHj1bCGsxenxTLVkIpnQviAsaIrlWIOsA2zT2nMuJT23QtxoDY6myUedp
043CvyaM5M/YDlGwz90DmO0y1iy2dTMA+gYFlXWpZ+i/gbOsNInIy5Gxf5BRHjczvb+fGi10XX7o
xBMubU0z3XcKWtLjcc8znoccjEdx+sFTlxTF2ULLJhERXACAvWSfFONlS49iChtN2CTim0fRcDDE
4yRiWw8WLtLJxVinMrcPp2QcebPeZmnyCU/xXaFvX7J9HeSXX5EOAE5WiklzIgSfeVpcj8NR6s1G
PPRS76UQxCN+FrWoPhhbZ8JkKFiigaa0J8cIgfCdrSMHQTDywI10Dc/gImGEtV1s7hDQ1u7aDN6e
xwaEed3lXjiNg7+wTjdQLWglz4+gD6N0dHzallXxI9JnR6UoqJVQkATcc49v3uiv1ytzzpz0Siq+
w39JQjEA3m2KAcEJVYJhgpIPFgu8z3AScGrUqPZ6/MM3KHOQnbCk68w79vK+6s/iHlDmel2PxotO
YZZlgeqN1GJ5PPb1TtcWUtHnqPkjAHZeWTafD/FpkWY155be/rXqIH2M4Gr3ajyLLTlRtHMd44ny
tXmQI07fGFlNSKhVu1pKfKD5ov7am5blYvsFwWRq/K4v/PVWt4OYj8yQ20iV9AYdOAFuHzKbWRof
6r4nBuwt4Ds4teDfwQMEbQt3CUEWJBSnZlAV8sfQqAnAFxIQu8DGQTuEUd8kNDRR+gaLU6rQbXOc
Zmwl7D/4+G/kczj4L0JUQNNn+sk8IXq1i6waKzQCdra7cvC6W81Gg3EQMLS2QGXkEUINDXoMdf1b
Fug6nSwfBnmBzd+Tl/DSUhOzvQQ/Cg/mi5Olhd53opyDKAqyZOmjI9RrFmywQBQ3ugSpT7f3X3UM
alGLwxCp6WwdcR1p2bci5Bai1fUdpLMZXsn0a4+8hcSbSb879KcVAI8ACXZ5Q9aHXVdbbikrbzw+
LHR29T40FoI2A1Ew2p5XM/SbpAxSd11hrRIq0NrrTgckJ4w8T8fFa+YN908c/uie21eXRarGcq48
A9qjO1ic0/4yi6cLqe6aGuZ72Dl9RmR8Udw5dM7jWhbQPzLiVHHnTW39ZTcWUL+CBK7weugHYZ3B
Y6Bm3/0HTwHJTkVt8OcJacKwK7sAhyoK28ig1BPOKsyc5zZ+tOq3BY1ZQSqGoCmr63kJVuG3fqeX
4KRgezvJb51FWGhID7a64U2RR5mHBaLQ5TYEegptLnvNrp9Ek7ucYeX8amUwL4K5QF4Il1kak31Y
GXD+YgYBzqNgjE9dCEuLyBOlszuFrXhsrCnQJzhZcRA0K7DR7SLB2Z4BidO0zrNjcatjDPDB0R15
pfa1iVGh3wI1rwXgWZhsPp8iKqBTx3Sxbg0sGQ5cjCRrEo/9jTguMgIHL+6SyrOgHXMWflNy4u+V
meB+XZYt90CqGbC3GvoMaL8SxIpnA6EPkSYD0LzJWm96KKE0jBIEIJp4JVEwkHAtwEi2Zwee5hQo
QCpyCNbFtd8AJ/HLXn3/9j+oQuPUw+EOr2gfkr+IkdT9WEuV79W/pFXeiiSfIXo5ccTuKcw6Y9uf
sho/LXSFdzJYFANeG0XWEZ/qUVX0y7Tjyw/RvYpZXre+xp0nTjTft9PpfbLXD5vO6ODVoI+wDD8e
tWpWy8g9+WN6Di1LMUoqrVCootNvGxMrmTXm4EtwvZc6xFRakH7pZwG/3RoD2TmI5C6HZBa1XTEc
/EeVemNjbBuyjYLylb1uSh7ssyodErxNFm2F/E6WtTep4vybBBMQzxOOxn0HgqNVvrX2YQnYsWZR
UVd3VRZ+EFIMvlV8WCV7GEz96rAhYUjDYPVZZFtXJDkVrM8Qx57LGe7ENDqrodJ5xzuNcEGQQD7J
azrjA1hK4Vb+A5yapLRiDghgHAxSzZwcWOWoj0CC006+sRb5ILGs11ESHOYPV8xKPeIQ1jcCAzPL
FXSc3u9lL9DPZ/sw2Kll348WWc0YP1oW/an5AIiNjCEpPaOevzce/eDE4aUQ3JF+4PEg9ntDfvll
BXKYH0rIo46HovHPZ+haX5frH+qymXcAKOWKx99Ebh6Sy6G9k2F+z9gXp/rNlUIvHID8HsvHta2M
Jj5JVqVzaxFTcER0ZuFp3VWubZijJYm5KvtmzVbC/JPvWU9p4a6lkFv/tFLvlGOtLDgloK7zCu3p
WsHYlCJOgmC4UjNeCq7XFvF1mYcwmJ8XWPaJdTjKtHWQWRAuLvFZBGBoVooksEiSSMZ3yQz4rb2I
unOz+7H9QGv7LAPA1lUczwxf/fGdYae2Mly0NXlwQ94X7tGr4/+xnAVCT7wpIVGWT4tAhn3JTtdz
LvjaabmHkrgoV6qVehU9jCk0zS2yqSg1VzmTB4pFnVEdTMePqi9AjKZnrpjsB/GHcxXI7f7aD9cO
32Vf3gUxs9IQhZi2M+VbEFto1Quw39avLi/aU02r7R1CO+bEuRzzDdBcydR/aB89yLfD6KhrOuKY
SheJseGSo4XqPQgtQqvs060bOZq4LLwianH5dj3/heDrUhQGTaHeqLMURe30v5YyoEoSa3zweBq7
sja/FbswQ1Vf1VqQDga9hyG7HlDV93PIfnLZV/QJ6J7a2ExdaglWyOwytWLqH9jSTeWH3CAAxbfD
R46A9h8SIa40fmH3H1F+7ClFed2F0srCbgOoERseGzw9WGFywGQ2JFpAuT3Gtjoxy7xGSoNGCzmQ
UfSGsKW+pQayJh597cCKK37GZszYdLMxY8IKLSgfCeA4H5NMhLZ9Lt5XXZTqu0vBGmmytS2VARBi
Wf0GqdQp9i/UNRpg8Nut0WRzxyfNz0ePGOey76R5uWlegsuaEAeAu4yb5//UzS9yBTcjz/mbJUj6
J9nrfKL/4o6LS91mznPevAbS1nmbco8m9rwyivZm1nBNCkbuahdZ5njv+2KibPj600qTsUSEyqBN
LPu8mzIqoeSuX4S92r8LASp76MEMkti2ZzP8mHtnM5GaL8/ci0c8u7zVGumvmsFIaXIGTUOkfMIS
0PjE80ONhGeoGAXaymZTIUXisqPUEl8l/JcKrH2MVjHwNfAqfsD46JXDx5G/B7FMCSwHbH7loV/q
pkNrsgEtyXOezB//e8WWeMVPJsT4ltYT/xIJJlI+LAuUtxfFnFvFJUZgMHcnJmAhFu9EGPApzWib
CkxCIRuSsqc7nhYyGFYt5xSRKLZzOtpj+EFzLqX2VfIZhV4OmfW1Gz18ekTkgUY3pyCa3UNNy0Hk
vswS0B4DiBeN3/7bAG6lXEvzGEzXBDZ5F27u1bq0A6hWyuryVvRkTFQKBjpUJLSCheQ5v9+EH/ZZ
mWDN9gBCXRLjOW+FG2hp0BQXl9B6EXbjs/0GgkBBE9HGcuhXRDf68GJ3FmH9HgV+TePRPpq6840U
vzIxTYgKsxwKwz+tTMJ8IrWr2KoWs73crrfxgfZRbA6GE7SsdmzDuB6ZxuUONHKjLgXLOzDyxUos
HbOkHXFP1CxxKPnLtfAEzm12ZtGVS3ilCABRUw+pvRR2OALJJ7UHlwa3BLPeMHZ8kFYUC1USSqfc
CjCE/Lty39ktoHjrOqVOD9ZoNG/mvM0bkD6xdRXRHkBa3BrMSX3cw06BJw3sXEr+e4LF9XMjxphF
45HZUhYoPdk63+pmcddy45PYJDUETiBXWhFOmT5Rd8EeOUQw8VqoF/TcE+KC67cUY1ZyXj3c7AWx
RkffrJhbENQ1Lp9mxA3m7XoT0l2uV0/bu66f8jv5TH8Rz3yb8hx3lh/EU5xZzJQJ7LocfEQBaOb1
VgEjG59pC+0SUz7BzPb557h7faQwCaJkq/HYEha3kcEMdsI8sfgHrzlwbOo/X0uiJjwVws7g/yyY
/NHrfeV5nYIjQ4AJ45T20eM2UahL4gXpDrlYZzTrhFk0HUj3rPy4iPMtJOT4+eD5S3cmq8YUHNIH
Diz/qwu5ozIpJyJATpkfwgCv5rGIlTg/xunDcIRvW1DT8TZH/qUrsmYgVxnth5qz/h0eWFd9xbEP
YG5C0MowVo52RHMBzTI3s2iU7WwJUhIWnGswClPhM2uqkUVh/mFAQ8GKHHzA53NgEn2hYVg0lDuB
WNwllzuTP9b7butbb7MWTyVS3t30mughHHVMz5eDqVarXScEBUZrA8zJPrRdFhCiOm5b54ty9axK
akcWwBmioGkg7bAgJbX9dyxCfhOliXJ5r0tIwq9fiLQy1jqSITmcuoaMAoEIqlet5p0GMTD+KZmA
MIWcNKqv/H4cB6DDlc4YryHcVwfXTFptv1TDwUOvWcbee0t83BfIPl8UTYTPg0q8rB1NlW/bngVu
9w0j5fQRg5iJWgyL2TRH1OmkIHnylsNhiS+enO1Dhrj7DzJBqHL4uX+RUnanagvLlv8HQXfLMAP2
O4So8u1p/T/n6mEe72/+rXV91KCRQ+cte7+AsUH1xno2Fv4VmQ391zbOfEyKN25cG4JbS0SzHYAW
kTOID5HJ2evpLWJvaF3M/g4U6TgLfjBC1zfDElByvQbBjcOJfb8ugmvc3Dol+In24O9CCVljeNav
736CWdjkmuxy2Wv97NbTPGK7rLEruDd56/nmtNlKcpHC2xfVqUXNcNwg2+whPlb0Oxv2Bdd67PI8
+c8Y2uG5pOOvynAYfSBMQO7YEyIywL4xrdxRvMagsPLKErHiHO2WBOGulh0tDzP00jst5la2dv7e
gbMqZSRPX8rmX7cXVvFVmzQeAp33RCSbSOZ8szNayEX03E0+D2PFaZGNAm9uC2wZuAm91AH32EWP
mwfTGJVU6t0LXL5KAD0NNcTIXNWpk1OY7iEu4kPwqUOSS/ElsePC4h3QXMc4ISUvsdYefSyED6w9
oQwpbNqYUevCtyhNyxf9WfYGpkYcN1wOm2f1lJLPl0ONIsYhqeWtFmV046LAJkflAtDTHN0AvN2u
z7jX561SdMrt/Z22nwy7iywkQs7rfw7wYBicw9/SwvZ3IC7+6goSOMOo9jeWYLmr7DOXMuzQs1nj
+kqBpS+i68g4NAGmgd07GWNOuChp9l0wEToBM2px3bhSo+SaCffTwd+aUmCIWSjcG02XHs7s3la5
rm+g0oPXRC407f3BOe3zR5WxT1ZpWzCqQ67kph6Y/gPpDSx1nB4yFg2B8z9ClOfTNaMvsrXf4/fw
DUu9zOePPfQ2CoChOFqhTBJYNK3GJPNNA5bfxPTvPc0REpkYZO/CTLUygepNTAe8Q5bmvq0Udxm0
q8Msk0FIF81mOdLVsDhk8XkWg0WRWzj9iWtPcWZ6kXrmyyP412tQOJ6I2VtHclatX+1sgcuOw3z6
8TF6UgyhflB5WcDv4uEX5XC7PnYTeVp4iFoZ+u/mCQ1RN10aSlykT4lFA+Usvk59pZ65TQdZmeqY
nfOyW5vjIRomxqhd6gAReaZwjOsXuylpxsf1FjRFhMvyN9wg9IrqDf7B4Yw7SRwSPCusM2AKi+Qq
r+380QdoamUowRB1pMUGeFNe3yxk0WRqA3z0T3ud1sjeIfhjU8ysTWDqv97TEGoTlm9FbolHiP98
qJAbzucBcnmi7rUi0t8Gs4AVTiz5xgzHOegHtQdMMS+xlKxYxro44pHQKi4ibYshwvMXIIDRDB2t
XnWiEAfAArppDmLY9l0OdSiR9Xxf6WoLZXm6JVijpHnD1RZFzN8UqucEWHNBLwH6Fwa3/FnxCVyM
iwTK2OR7VKSdXMTtLmaVEvYmcJRG/I4Wf+S9Kd3bVXBHAa/7sDtXabNzUv4F/WEM4hoPxOSyQND5
6NxmbKQfnv5T56PAhn6Juhxqn39UboUEdySlRseMfT7IiD40+sU96PxbD5a+v5DTp04P2IzYDdGF
9vFeYOGXlgQZkPpHjPM4il8R86orjfAm5Ns31DuF071dOfooSqAfJPeTxYYXHob5eir+hv+ZfQGF
nde0RaqVhtLp97NQBERWMu7hxmENoOeOe2JQg2LOIS02g9x1o4j7kEjoXbaJUepJeZ+8gGMskcSQ
3HXVdX6t5HhhW907xEris8IMlCmthl7Vv1vwyaA1U6uVS9y/2EQ1HCCFD+yFDQFTCHhxhPEnZN1D
lYxJum5YI1SodoiCSbd/nKTOpa1XP0eXteR64S3/h7FeiSE3Tb00g5HHLdUWH39NeC3Q0yM09OsQ
zo6W5LKssG+AcP81VaALGyfh4tFDRU1jGv/bh+mbN9IhT3Lt7776ANSTMe0ECSWXpVLhNNjl4Ctm
i1fowm0v43XUEy2lc1gKJIMzfjdHqRP4OQXk0tgUP6QAbaFN758NRBzU3W5e9MjM/cLFNpPEZh7y
ml0NpHuMHC9tC0ZPB3Zpe5CP5PskdNryPdYiTFm+h+zTQNlT7MvLrKXf+NNoXJ06ym+RDLN82otl
0RX/4WRy7NzG+S+sgnh7N6XRFc70yLzmAC51Y7APamzwJydcO7uLJWfC57eyL2Uy4H41L+/XGhtn
bdRAkIQWdbJjHSpCW0qSBStu45sWlipBhMUPeTeWm+Lg+LtnUC+LvN0lllEbax/c/R7geZ316P6s
lIT68lVel3FKDViEwWuk/1Wgv3MDvp+098Jg4T67am6IUXrZqpS07uMMKrTTdEJrkawNsRP6Gja1
rRh3KgI1jDPzJu9+j2kwnMYhmgo3ePj50Mn/v5QC69h+BLFbgCNgJVTjLbt3/dq+CZL/s/MUECEG
kJrXAAG56MxFBUlbWu+5mxGUpAuDI6NSSPrRMcxN8GDPXMjw9dgzZqu+UNrlhGEC0EdW+krW3x/p
GZsjPDPDEJDNhuszWI44p6MmMQP5/ismmXjY0ZafpVZgYDeymRE1/1ihtbzlJgkFreyOUHospsX5
O/tEZrrzko2i1R/cocK+seLaHwH6cwsxeZomBox5A/8/k8WxkazFCWX3+WBMXp4YvSIWW7rIXy1Y
OoOjUj54ZBwLIEgnG/1KJZa1iT0g5uE+tvYtaWWGGZzRoCSzciVJSh56FkMcqcr3NDxPSPOXLDA9
k/u9XjR7A/HGGKWo7kxAli0TPYEjxRYd1OPO42XeStLchiWYByCyIK/Brrl+uo4d3u0Y7FagF9NF
QbJhgp+HSWBuaEzr1urNSgRIjc3IbyoNb0gpoV+p6G/hg2Qn+SQGVExfJCkqoE8J4+ZW98Nl/Urz
1QP+ScwRBxPotfqdz70ZgzA0UUYC6aLmcZ5w1dlk/3e1mc/JhD0w8aRe99C8FAB3iClgxUkS+I1S
0q5u+0rGEwuvgaGriwk17PI6DpLkQwP0E9lRyZX4ujwsIj/Rennumu2jA7JBOBVp+eUyCnwAZ7h3
VM4gAnJGzK5XEE+9zi/jrRVM4HOr6n7b+hh7KVZT0+3FzWaJBtwn6+gYYXhZMowFH1ORorNY3pCG
m0m15IPWi3synMHS0LuhLxgGkcXChQl278E2SjM/TAM444/dxHidaX3z4yDeoOdPt+8vOWxOSDRJ
DEx0SzEam52/28wE/S/K1U9rNEc9imBq8uBHhNiYOzp7Jbg0dwG7pcARpNeCtpvxjN20pfLV0QEh
qXX0GLXJ+sf35WZ6PrgE3KCmlG0eeVdiWWQqRjx5FVxnzscI2vfEDfeHbfPdrNjoTR0iTlkKjkus
6RMN/UzAAzWJqxrOrLy8u1kppA4VsdphElW2RGNZAZJLVtZIwRk1fHDQnlgXlwEowD537dZ8e55v
eZPeY+xyDLYSpGYb+HWYI5W0Qc01hayzriwBRAcaMyqXtcOdw7Fv7DN74Z7wtCKXxIh8bNqpVhxt
Q+uJBUHFhRlE5VwC2iJTOhi/QYyjhCow+/mOq3IwQ1fCLBxi/oytrdbP2DFelfNVeGpe6ytxzlEL
gGS93b12tXAfllbi0y/r2r7qAi4pQx2P6Wmd3vBpNhPfo0guYtRmdgqhEL7eFfBuNq1Eo/GGV+YW
fZQGkQ2EcklPRTyaMA+S2Bp7VGY47uKcQNPmarHi3inTM3bcPMuO64Io6BPWEoLE46LjyVnrBT5P
kUiU+NpNuYUxTtA7siZI/zTP6wBuvG1r9ToZzBhHDXY0rQH85f5Bfn+FdEgcJf8bIbiVHMWXAxHO
L60mHpSMkixVNbqPlgyBAVNRKa90+Gz9LFOHJghezuK961pRs2zayGA1BkxtLPdeeMDTRQZB9TgZ
DFr3H1KYr1fcbANIvCo8s4sU+kTO8fnlk33sop1cn9r1CPbqOTUo7b7nbYkme/tGmWU2ZY9PrFaP
Ycbwt4J1N/5PcRGhElr07y7AEX7AuLVfoMDuhD7I3n3za3oiRCf5QoXNCstmF9YWXd8CBhf1y7Zc
J6voizPolaQf2WZb+YrhNMIMrcEDqXkZgvEL6kJmjO4MsYfVjTE+y7oeuasEXP1XUSj1ikFRriIq
4AL9QLONU+R1dv2H10F2JE51rWTHgLMqThVoYoDMzir5I/82h/IxVLDqphPdbhu9QuNLpE4jXxF4
uv2Ks45fdN9teI7JA2CLDCzf0n+jSZptaoq+day1B2o9nlev3KhqBmDUzT06/p/KjdMX9naXVoG6
rcD7OSA+qk6E1Y7gBNdPm2zRtrFcCtzvP5quw4f6Ln5qI1j7i0aa1PiKls7WQupAwsOk+SbOF3J3
BZjvqmZE1mlmlk7Cs6ak2HqMCDb0w0wJAW9OsQ+Ybfvhjagow2Eu5ItNP4CmcyQcB+EFU4g5rFWS
CCHhn0oGShFuapR39nrC2ukjI0m9/fVOna00vVyeqx44AsbhmzIXyslnAZsRYP5qZkN5GRL8TwB0
T1bekVbUHwbbit86tYqMPNsGPs1tu1FtIbgXCqXxGCNT7XsD3ryF3r2MkQ1MSg7Y7j5iaPcYqLON
G2Zn2qC5zhRqNo4YxrRyH8+JO1FWd+tkYhjHUXF0vJrP0HEYP7VYjazzYfe0aGVeCOYXjaJq6fDv
U3bOBuw8f5F/zCQmUwD5xJZDLD4dGng0Qsya/ShZ0F+Qbj8/xvxNVueIeIvKjj6dSTCVPjyQH04a
pnWXlwQLnYKWOZ51B160oBjGo/RU4lxazPYLDbGGNgPRFzD8FsUdcRsjlVAXDwXLBsyzWVJFVKgR
f2ucDz3++iGchfGdUyUZCPIpxlphDAhaNtf42Gnri0OxpLp+OGjBwVEspSySuM8iuGZG3Z9PKL48
i6ngrn49WE3TaeY+kPctZRAV9RkZ4oGRnkKttH3gp20jUPSoWe27PkLV28qPROvS1i+rD2yVi8ru
wdeNTN0MxQjVQ0+dgeJ8J9YEyB35rg+9+96VqvkBq899xmkpjlIoVeJw0u/oUjjMb0wL4qct57Sh
R8jlaL+zIfpFdP+vXiwulkXBehNWw7I9uEJ1LK+iYzq1qYEQpv35/gIJLce0r9fTYbUX00qobhDP
S3i6jO800p4HunaKAg6y98Rhbc9mQLfBeSsqBQ1X09xju1Zee5AoIA2FADA8oTC4BJW2KB3ugGA4
nrPKW+Klk4NnSJ0nBgrBkvrvRJS5HDAa1kKBIibQEBRk6MYTn/8kqhJTb2axRwNydn3vEkywoTw1
webmlS1D82L2DDAm1kev06AIN/Yu5oA7ToVcXZpjgM/uad9b5a2N7m9UU5YwBX4jXMGSX3iuTqTC
BitVL5/jr4MrSlZMBXEgERuA8LWG4nZU63h3FBRsrmJ4JyOOcBMOzmf0pCXl6yZGCDdaDiNVlfa/
mQeE3KX/h9t2OEi82YEYP22DQkSHGmhz8BcmmM1nzxBaah5Gr8gXfn6WHx17JxYF9edFBV6VbgTx
OWTatCg51SKT3gx5v5sNtphKBLKrU+M2ZcW6ks71uN5iz3ZCOIzsiGKUZAvuYiJVGLO2rQf81I+i
pp1dI2ylaESOSVrsrDSDZlpuO2i4VUCLGOxdZA92936MSZH749svbrutO+A3IsNVWVWJP8XUEH/6
GJghxAIgmgyrGFLOWfQJcDi17tS4U63tlPW4qMCfG5Jzae68TkrWEMtykjsGUkdX6MCDWEVG/ode
VPu9rWps+0jGqwbMR6sSESi3D9oI3VJIMLlyg2XOElEhD5LVfY6Zrlj+6KBFS1iTyzKd+Cw8ctcy
CXQBFdmoIEgXyI5n8PdEUnM5auALwSApcMMwSwa5uYK59CylRZ7CvyLazUZ0dqCsOButYhHyvcM+
WopB1wxnsbVXFeA6z1zocL2bERQ0bP/8llqfXmyfgjpoNXgZ04GSWIBi9UEWUUK0luSDZvWPmrW+
ECLLGliTqED6CDrdXDrdy6y8cLuGUBMAo/piOoKjsuT2GwrkC7l+1T+2VVpenhkLn5LcFW8H5Z+l
4DERUgZxEHDO9xOR7suH8zueY7h/QqbMsmbYMn9UN2+j/Tqof+ZOhBvpu4i9xurgL7IxmwB22wK6
I7PUxlbO9aFB8zERbi3WkgNnoRvKsUP0k4BOqRQ9AQoTNFTMvPZg/z2Cc90lk+RBreEnF0m7S/Hc
03yXCYpvfX2w8bTLfgnkeoXtfi0fzbxcKl8tqs3hvp8CkHJXH9rpcjyLs7JJtiu9keX8hgEqlexW
ytJTz3sQIBDhi37m3UueNnVsWEjUcmk6y6NXDTmfA+1z0ok2dyWHgSAeQ9P/o9qD/auezIeEOoNl
G3cqABBhuBZ4+1Q8wZ7PHvFPptbbiOpwPFl46eImpQvnTNBM/qDgX4rPeIY/9cNgPMxnEwpyyzCS
ex21mO6zoD78R2xWG0gp7ZpG2O/8rolPj6ihlzaIpxfe6e5Gd3peOXbb3Ysijlp2pKu+BVQ9oIS8
uyZ4vA5c7syy0s4FdEjzPzGRAMuGybDeoeu1gSktcSdSd5+Y5HJ3lj2Abnnj5GN9Qr+6SiuKuirg
+s1afOaIl7bKmVYUR3MkQzkJvh+vfOQ+0uF8VN4//ytMY0kZtftDHditSrMEtH6K3Z/0pQV4+bNl
B/FT02lkhQ5rDJWl/XomKtP8hOuJIL5C3RzrZ4JmVocC7NzcMxAjvDYpLXrOiwjHwqAg29EAIywI
uzEohhimDLnG6G5M1lQA7E1JZAVmuYJJWrdL4nVjjbzW5kpxdILMOuq2BFfqCABGw6OfhcjmwHr6
uwe+Kqx/wnP+dr63vIqSnbLJ9/5AmOrjKLfEbcLwfR38SKq5FOhH79NnsHQN0wEHA4pSnqvF/7Oq
vXDRgM5b8/JLzrjczgIBwlV45VO1wrXhxTpIKomK3GOkwzM2ZRLU3kLgGUQsGEW4zKCb+5yNErJu
B8ojl/0NrPCABihM8bHBVwUz+Gkdwa1lCcs3K0zcCwXtW4m7Z3eidhIcrRYveva9XepIg0Hf1iP5
m6wl8tDgnQd18sI0oaGH/NoN6hBs9zmO68nfzf35RNo9uigTpNSR0Gp9oQVaTBGuHTcAGPz7bmAV
OcchR0krRdphD7gJIQTth86HazPcm1QXWYmaJ6TmlV1SsR1gw3B1yKIuWbtB2YXuc6GdL9nZ5YB4
oVID0I+tE9KKB48x0ymRkTbeOVD81wwf7l3p0gsrdw+sP0d6UyPM8RkbXjitkTtlWyGw14/bJ73D
mjePAn0wHIOWdJL5sEeT9QVhMH1mj/BlJiA31XRlXtNuU3lIXmzbMrKS0hOatWh2+pwfeSAS1qnq
G+YHrc9r6vMTu9nh/TX6NIsqLIt2Gd4xwVLeMWMq4CZAjuncgmecqWZd1zXc6OeiVMaz7yarpZOs
KTIW2Ekpe85oHjbeZsjJtokRb+qLtVqPsqoq6Myyot8Z4IeAJ9girNymnZvfXaHYO5QXtAF2APNv
kXd6SHfh86bztw0/0IxWpAZWav0VNPsYQDHiVvJJZsEZcL0scXfoi44bjexm1KXbtPYgN8XWooca
JtZJVRW5wQVJg7U3HYbe64JZzcahmqXMUsRqwDbEmKB0/ARUAQ2tM0yb4VWshFMNu/0AR18/RqMn
PY/Bt/7VBlWq96MK7jQ4dW5Xh3RA3UbQxK439osn9epLgaeGUkL5SeEfIpI6q51Zy7/Ypd/ydc7p
w5tV4l96h/Yb0atbPnxCTr6YzEhVY+odl0Tl1WaQ0KE5v9fmOvJr+BZEhKTMTVY214re+ZLVUHPy
lerAxBlbP/4BVWEavlkuPZFCqFMVfFFHRjN/uI97soRNpgsovaKnxFLGRZE/pIZn2MxutSy+Z+nf
UZMCKJF2h1Rs9k6xIAFFox4ZQpHu2BwddCPCVrfJttH8q/tQn+lqk6E7n3Tv8fR0A5H+TrnmtxZo
GPofolXXgU32Gi5l11gFfZwo7HFlT4BxW7hrCKohX6Oy9nw+sfccSfrjCxG9r6doLftz4d2iQgg/
Js6uuf+T9DNtCtG85x7Mr2L+fkwbIg+m3p9gFAseMV3sp9VoChed7jBQyeHYBNSFvrexuZxPJ0PJ
5Bdw+hJTdqN+cnCK/xF6Csvit2oSpJLUlY8B6BWBCM2588loQO9iJFGYRQNjYzCS4gozbIaQTim0
oVxBqRdEKXX49EYks6yJPX8JMStH591Q+FbwXr42YeTLesuemmhBfImcE7fCBZqexZnWVtbu7tBK
48YWVzENZECHXDKQsqvdqvRzFbKT+eOItLP2R00oyWvDLtR2Q9/xDgEsXfjDTLi9Y4u5EcZb9kNy
ZMd0HHLeFF/DV+IUnbMEGCWbDff+XvFF2mF4JQMw9H5tZtZK5EDiUSTMiOPOmsWec3rI+iwvwjb2
sWtI6NUnQzKf2vOg4dmTB0zuaLqJcP949pgT+0s6Xf1JCTwSatXLD3F2bC+Wtesm2NTsIGaVD4tY
5LVt0/L+uclTiYkxHcQesC+uZrRPr/OILdnT+YL8PcV1LXcZ7EKHCGmcFg0RSJDjInNgJc2nHFcK
1GSxzvpEJhKIW2x7wvuq55jOP7AZBl5BK0OvUdhoetvgBo6PEPm6BbIySPrQG5fR3KPMIeiPS4VW
HQSLKv1HvLRbmF5iZQoPMrf+n6yPrZz9qtYYViiiLVCcU/BwSUV4ulRbZXl+UVwqUKK13pB6yPVX
DYHNP5JOo6lAA2dRk+f/X2BBiW0tJ6/+/Vub1inSdR6LlYrrNQkgVudXuYtT0FrAHnAiYExVopxn
1eQBN0SUF0+t3NxHc2llPVXlmcyV9KBsUbMxlw/cwWob/pfySrBKeEKXnBMGae3R8PDul+YvbdLT
+AOkpoMBR7CkYGIm6RktiUiYuz2/eQbSMhYYpp4qeQfdXIlNDKBWjnGNSW7Ree3ncj6jwt0erRzw
UYCZqKgf+zw0gwfSMAFK359jLDVkDXMXb9EW4ryFqD93MTsRia0NS9n1rrEDbI3HPJbAl25AroMC
BKhqHiDAVViVAlD91gak52rqB9VjsZKyFCww68JOb8wq0ou8FUZeQzdM7jZ6ZdNB2nd4GKpAHr5Z
I06Ea0K8g+TEZx6iTJf3K3CHuZaUAZ9oqeSPr0bzJpnOIe5Gui06Kp7UoB3a7jKfxXP83m5fl4Ll
jNNl045rCdybEO7TUg25Jay9EDsFDvGOaPDX0a3kays4Xvody539a12j2FgId7DcGQWPHA/SF9VS
Jgk30pIzlB5gSBK8dvpZGQXJI+F6P+PHAnRPl5i4YvRQy/DUFqPJ/K3lyGAGFJL5dUkRuNMEo/FG
ENylMkBDCjgw+wfC2VtY2puQADD/YW30b25jSxtDHQwEcmQK93280YQeuF435uPAyJ0TpR+8FwYz
8KTlTiYFiD2Hb6LxRDFzkzwe+EiOgUKwYG8s8VdwgAaCldlc6l8znZ36MP73oB+Y4WwuQn6zUeG4
VU8zKLc3hIaYaDiNIriQG/Mzstc9xjOpzkf3j1gc4xjxk9wlWJ/Wza5liNwn/2bVOu32ye+fzl4l
Wv2IdTy761Yf/AQQ8M5WfyeymJ8GwnxQ1oXjGU16wwWFPJc2TkOZ0+kPng1QlzIAKe/J5V5phItC
KCBU+mlzNoc0lYn4GJdgMhgdznH8MedF0s0taIURGrQ9VGBqAJcUuDKOw9GNz7KU37nbhqbhFes7
314pODum1fyvMkI7G9TCQitztSfKeKlhmrgQ9BKxsJTHPQvU72n4/badpfaOaHGgNNc8tl8hHC4n
hGM9sMekeLB30SsYEtZtnBi4tlsNdEQRt+sad2Ak9VeneeWI5mtLBZ1CZeZK2jt/2wH2glhitPbo
46bhZlMKdtJHeQe04sc3iD7hzL/6HbH1r1NydVwzMU5up2qS/WbHXeVpzJ++NMBUH7EtNlFcjVVY
yP0faEUhBO//NS+2VkYvnrECJ+mnx9d+Gy6uulzrMFlR9GonRVdTcYwLsjEYzytj1G/2ZygCHc7J
uyQCElTgrWjRuEpMJQkyHwmDbuHxtg1kqt1s2MJuqwSuQ+RYyJsEhpI/l+LrSaeaBiadxWC881w1
TfLj4r82tnctNxW7B+QYOiG1fUqa4syNXRjtJl7TSoO0NsEaV0lafoY7V1ihBIm5tjO3fsNDYBAG
dH2oKp3fv2Bu9m8QEAD6I+pRK7UCniInnQnK/KTrMK0DnhcQOsOg68NMa+0Dbut11EFsDB0exyIp
hX6DCm/+1DXqGi9006A+gMo929eahZCCbbSbNoUjhdeKgDN4Hi4t+O3yFJntL323jkEBuQMmXuEy
I1JWl80eIWbdVXVegn1s+3ncmo9/6i5MXxQQBsb607iJTDQ3xkDz0gQZg25YQPAUXi5ynAH8MM3b
J3KQVXNTA1SOOB0kcLY6wYYstw5R2zbvEzgsmThkvcq+YvFfjUgo85C9AV8MPGDrU58yHkVsLJWG
LNHCLjzUQYE3yjnviG5gC9OCdKJ2kOKHRyy1ti9N8i/R8YrNfwnxtnXbuZBcx1JhceQ2GlEXsqPL
2CePJ9qw9irM/X+6pC1hUAxmxJUylZ7WSqsqS9uR5LZmg6cJVDXtpoUktexOSaTc4lFT4iOb8JM+
6bN8xQGHdN3qpMWQ/4fhRMF+PeX7rZka9yHFrihOU4zr+ch7CTOkT5iuZ1D+y4XUHG1jPxiKwuzn
hquVSSdZtxFj4+QvQAlzndOUCnaXnC0qm4t4x5gtlySyopNIRwqFYUIRqim2qr8KVC3t1yDbS2qy
tal4a+ePSFkxFElgnJt2AEKXat3JaZmrYuOQB4E8/2aoUFuwoaBq+SlBZsSJd7YzHnnLYM0e/Q9U
4qft2RYAjo7uFgID/yAWC2jiNQRAKsBkiYGnadqfW56qc5CuumHmLuBE2sy2xfLiFuj6XHBxOiCS
MhtPLXstMcDJkgy+KpXrN41qyneE2KsmjkjFN3sptHvoBRal2Z5tGvakDrHG5s6PDXBLFuuyReny
WHzmDT757/yZwSyzXWDIOswJgwJiQFvHrLpunO3gw9ppHK78XpAzVDupIefvSibtenAtN7YrGx2L
7C9890LJJ3ppq96IBEbPFlJO3JwHFetHpzBZgS5YGgG+QCWhLg5dNOENDlYLE19N7e0iOrAyvkZL
jcgLyBS29BIWa5kA2b0nzLlxdJfkpvMy4+sT9dQxZS8uLdtPiPYPT+udiUnwefA9URpjHk7deNN6
7FGyAXYRQZbiTYp9K2/vtjxShYpitW7uvjYJ6PBR5tqcGO2ZsJe69HF0w6rpVNdnGkKqEMnMSzXz
UrtQapTjtmZsuiMaYd2KRkITUvJAewUvBup4H1C3LFpWldzcIC9LbfJ3QP9VUjskYg3Bu66DxneU
lK/8x/RndbzDo4WLBKHX1A1kWfRgGiIcXgeMrEoimCMVd5wDZtWEL/1bCEWH3Sk3GcR6Wk3ZGBc2
x2AT1vJHVePKAbM3KKTti8T5gaP7n0mSrVqEOCuixy2BfEgqEpj65Plkk6IcBGDv6oAZs5fA9cm1
+x+alP2TL9hM5+3ybTm5sVDSS6ktjrkEzIjH0e3p1G7IxFeJA17M01QTRJ1aShT+JeSnBB9d47sC
ADNtLoQ5nT0eiGvXcrRdeolQdPfaocAH5g4DwTxJWnHnzHJOrBzuAIvOkPLboEXZE85PP8x6d22h
1VRam6u5+omPrqUZS5YTLcuIaXnTjTaEWeUd73cG4jHZyf9pDefwfxxuGC0935FFqlSiJ0O6XaGu
KshOemL1ZkgRb1A3atXlFXMvGAZcgd9xynIesFD3Z/UE2JZZ6xw45bOMAePtrt3qIM97VSqc/yXq
3ll1W4S1tZ9pJVFyh2CrReHfUGbQLzpmsvpNXt9EuqQcQQwdGmu/s7du8OQjxeovvOcxl0WwJoZa
nox2HpHfbZCyWUtjQ4fVLbulWlUHhzT1uR+RaINNl6S7Sw67Yj/p5/D+Uk1NP/doAInQnRHqb8Yg
9S7VeVv/y4+Mi6tK8IgFhaqGQM4BLAnr2gk1hMESPeqS3p+IRpl5WAkNX2DqHXppDyvs2+FHbb+t
jU6ryeI8n82+QrnM42zQzFapbPI9TRr5lEqmsQ9sNVhMYpDItwV8cZJ9WSzfpDz3tmMKg4UseVav
2UnabRmjFt3yi8NDKcnUM4EGWnN6+Cc1btwHJTlyNbQEfApuqc0pfaDMQ8a6WJ1X9rl2bc8Zn9Rs
NeTY9x0Y8JSfHoEKrJcmpOnicaWVzhT3Igjh2m3E8WFTBSHHQBfqXnS66PLMSnKgEP6lsAEzio0A
d3c8BAcCw/z87V+ukjgBnxpdBWqwlb/Vtzw0gXzowaTzYjoeD0TaRNMf3vJbyAbloLgDAH7DF4E/
s2ZurrXdT2LxXIg7/zNAqBpFFYa6XRcdE6dlct6J8fPZaHP/XC3CyJNTbd1mbvqg1YQXydugexT+
L9dSldrV/s6Kj1aEtdIF4vwlFZbZ21r58daJZ5DJG2oiXMyNz54IKbKOYRtj/JZB5BA26Vmi2LTE
8t84mkxHLWfmaBtu2b2MI8RHSSzPx3hynzY1dITeV21cE/h3JJ+f1TflFBy0VTF73U3kmmuUjX16
frZnBQz2o8VDP5285RfDXtd9ObG0eIJP7mgRRO8EoshccGEb5/cCL/KftYIXI7IrpabnqwHxSRXV
oskPggZ7u2lMUKGODlEpiUqXUuaXPPlDyGFJGVX0n9+AcVfHmv5Awk07v8NXRj3Xrr9cZaAfH60S
WyMZB2C7UNfriCtOVZJ6ySW6rdUpY1wXv9yCFKYY2PW3Cc/+TP4evJXOZ5JS7lamqgY9hjdGaK8a
Di4mkgisB3NXYa+vpLeb6X/W1vlw/BEpm2mVfGWvdtgu8zPAGpK5xY++bcSQAX4PW61uUtuepwNV
c3XWbFhzjCSbOxj1FuiKAxON7XFY8zvhTScHWCMyhhpOV0UwmhjiXUzZsZqM1iNyPhtbJsba6AMs
p/BPbJ8KXCpwNV/k2IzhhhILDes6KAhnke9c9xyWtb+XOG2lb2/6UXuiGZ9xOQdahOvVdtgwMMK8
/bysKJlCNVhTYRZ1FdDWW/P4CS9IXd/fUh8i57L5sbmmmvCtDYzSXgWbZV55iy4h9+aKTEoTkUH4
B/WPP3AFpeALDMjOCSLYn+U4YXeG8zMHA06mSjX8oK/T8FE8CyBix3uJoCu8Mfu/krEBusCzEY7N
1/dHIzODP+uzx2eHSVTrUi7wIXvib2PAkSPh2MD1qF9F0xdD4sbb0SbpE5/Blka2uhtixBmw4RnL
vWHGAXdHUAWBUudUi8vOPjTbO1P8P7ioIu2GOgMtnjoeMy9yz9sDcGzyGWzvUj0I7DeC6WWEiBnY
Ou/EcquCDJGpx+TR7sj5eTI+3c1paq4pMv0hJgZ78XQMzfN1iaeaM9+7UqbleMSsLNt0zMISFMwU
cyJIM5NgPUAehJJHlFVHSOwKV5Gs5OPATYnVq8Sgo64mUWPYOazZul1e4Y5flVZEa83YQ2VYhhMm
TGTuS/17dyV4x7SBlWCZ4nfbhzvt14vfAOuzSBvYQe0SMlBsz2HDIU4bXc68dDWl63CRNN/yXoVI
kuL2TsOQEKTgJ4AabyrIhZ7gRMtSQxhxhlPmlxwY/4Y4bB9Vqw4lPcRp1pjX147m68ZkhkQBSZbv
Gq/8bOAbKJ2GXdQK4QB0w7UVxKJpCuKEGjbqtTA9sWHlfMkbuxHZeuRJM7KgvlG3v0pMC6HbAoPA
ktm7P+WShEh/WeU4yRGCfYidq0UUbw9TNoYophHRoxgWzaB0SLJqBCPL2Fx4b2kmX1IIaz5lxTtI
CToXUQHyyPXFfQ7+yV+dinFed86q8e7HDuytW3ewoXSIk9jP60LU+BCoJ9IkbP3ekQ7M3H1/A1fk
EnDaPH89WlV2n5tjYwn/qiZaTQxe6HHO58sDTSdZdFMzdt0yA/uYa0hx3zU/yolbRcUL/P4P2WXA
Re0cPcTAzWrzYuOticmVxKWlfCwYuCAI5VLJATqiNddVZjdR1mhLgFUx+tORivt0lVfAfT3w/qvs
ZMSQOobJsQJao3aQGdRytkH69rrd3AZyer8erQnQQrNTxQ30e1gwGiOghk1ROEPgjZz1wrmEzXfi
FUmuyVVeUvAcKmUcgrtevSsHKyNRTw8bHzwY1mnHOqi/QporOMcs7feX9rgOCKwiUpGWIk9PxNQX
mIPLZnssXhctg1jKR/WqA1WNX77TKgOA0g6cBHhwVoJX3RdTyXMmOqV9fyXIsxxK3SLBjivYDB3M
X10FkRjesvYAKIHYOsl9/QEAOhgx4ivuP3r+o1lL+fTBYthJpaqLEJ2ntisJsidgDGV57RYJ28Y8
Rz5WQ2VasYzkkjavZF/7P0uiFSn6PU68hXWxX7kh9RynhGWQJsJv5qZC/APCuJBhH7qFWxyyCBSt
XqK6SnxXqqU4TirbLWd5vOi52AyT0ur0p04oj92rQr+hqT21iSf66txd5oggMg560Rf2fhaqxy40
V1BCFOv0zg1azzkaZ3JXojUTrPt3ERtPPEtKVvQQx7N8mITxgBxs+TCTXtzEL/yFfgFdMnHIDQZX
XRclEkK2ODRFo+XOJMhvLmjAI+ce+7/b3d025Zl2mvABjBRsdb3acFb2/xc3N3gN7JM65QwaozJ3
Z2wxElPrZ218coKDgXIQlUJvL/YH7oOZcAW05w4jWyiadzgYriYoIWY9iN02RTWT4PVGd0XHjFAG
5KU4Q36Hj9oqOl/7CKJATT6tSbniYdRgvkgQn57pS1B1cvo5xjieobsdbkCUBqzBdyIpmUJpmkMw
ruKf09xurFVOgBUuz5tJus4uLpdEo19ONDl4czremAtcI6pZHV9H2k8eI9qtG9sWEygra6PEJ7NN
yKr0TYFLczY0P8YNOUzBBafuVWi7TbqWB0ffjyes1n+UIpf6wtXsaatyzY5985kg4DqLaQYjujEV
++OzbIQlciUBCPWWygj9jdnrn1Tf/xguqNoqpfSsa6ueadOQzoprEdS19KewBye8ywObU0uGVjwE
ZtKaz0YITWrljbPwBd7zBIYpAismJDaDwap1n958JoNlOh+Hj0kzWIeIjGT3WG2zMoQNSH0anoms
twVb/QZkz5iowYw1ziV5VdV3MFxbjjENiHxSpAzyHmGjyiF37xgRXVNxi7bdl2qSq3gTlnhvW+yP
grbFJaoDbF9dOJdmXx4fnYXYev5kLPnDL4jKxR8f0bsaCQsH1VDUc6HirzGR3wRI456ebr0md7qo
Q619NU4bM+SCE2G8szuoP2ncgAmkCERB/qVW36Vik+py50RxCdtgRgiSMLCACFwOZ8lLAGmxJ+Bc
rOCo/V/wpjYjcpzBKZB4R0unR9N1p2qdSEXRTEJeQdR9+fvl3Ap3+GsJ4nikfKyUMYm9fne8AWC8
Nh9rn1RHHAnSBEDgsYXWjiUkCMS2GAv4gNLQ24KPjL32oehXTQXciHjcDQZWNKJCin5NxHoWUL3T
QD3I4GTQv4Ov9LZLIFi2SrJq7TJy9lYum46xHgiS3qaH111iUoUKp/w3l3FAbUTpvVueggKGn7hS
fNG6WWpHlsWA9etQZiznMDu3N2rSul336mh4TjnXB3RwDnT2dBr91Ylkt0NPK6cGCvzi8MPa+m3f
FXf3MVxOOBBEXzsS6rSkkUQrQSKaP3XQ94/er7NshLLst31YE3hdfuTUkNnpujPhoxJAuffkiyjt
xWkqVNhyFi02Uh7nOWcCefs2FOFR4iHkj9NVf2vfs7bp0/3Xs1oRM6N8bPUSD7inMv8oaRxExmNn
Qqw2PGnC/n80Ddlc3yOCC6JHhht4NYPryhpL3tKVrUpQ0rznntg0XOJoXFp3pfzEW2BuooSDPnkH
80EQZ7mfaI0lbvo4Nj0gdug6cFLZ2i2q7cUttsr9mdGwh8GNSbmAdtPBHOMldSAT7rpS3c8y73tm
Eor/aXLqmOwhGy1nT29Y+mtpx2Vqh9qoaRMASeUxNdc3nxbYMzP2//Lj6uKzDCiP4GQGA8SWNEJ4
uH/ar8gySVw3UkASgucWNSx9Z6SLlT8Imq46QpcBpAHML52bRSGhACqT57iob1Av1QqKtNt3BcvF
gValQBR7edGN0IwRkQnraL/5U8S6fZen7JyspyCyyxjG8GhLILVfNwsRkgOT3+77/BJXv8y/Ujko
0MYXkgxA98fQVOIExrFesb7hRIVgVHv2Y6cvXsBD7JM+R2iWUtmn2oktQgvDHN8yiCOVLcYabiuw
apsBogpTBwfMl4i3IUUpLk7rjJ1WXK3IG4vYpb+dLNFjxu+aSiemlWIwAIIPe7H/Ky/GWT1l1l5Q
8eGHspeBQPhUY+DVJH6kZzu/jbMs40bvtRPhx72I+bAHrlFeKIphbNbar3+g66wqoOt3aRTCNwzI
7HcqkZKeLTbS0oyf626mlDHLgp/UrfW37zHCsQ0FmFFO4MOABP69DW0cG2/htSv6XgKwoPsHqPR1
8HcqnWYtA7kC3Dml/ts0Qta+UX751OiqiD6GhO+IHwXq37nHV9n0bV6rIbw+yfYuAdIUpPxaJqoF
hf61mK0dJ051d4kP97UglV6ilsmqfnRiAZ7tjQV+v+PNk2llsJ2qginYq7z6WN2GOeVTC2j98VyE
CWsBPI/rR73yxemislWYQRFZejG+5RT4OXCVFqhr1+FyxddFxKpYAENRbXhWTu3PoW3jdEwdU1Dk
oFsj2IMOMbhbRMtYsQvns5ALetjAvCTXVV6yhU+4+ShWpzSDAPnGAcQKIDeSLtcO5qnDQqxJFP5s
ozvspDhmvZ3RbpaEwtx61jGbN5KfdweslGdELySX/27nfYDVQWy1D2Q7FN3tqyEPPE9OvMnksLOG
4qNmiI6ynAgy1AgJd1n6oo9TkzlJaf4eWV9OA+8coY7lvcOIC2dYs94HTuJb6naAzX5kg/6JF/ma
Pr+LNKAUTYmdDd41W3RBWBREO2Up2hGFbCuS6SpBCoSx2g5FSJqGjihN59pVHeRcrxx02DKpWXXh
5J7PQk1orPoBgQeFaSoS4L+ea5AS3OHC4aeROgoBWYGGuWCFRFmzlSthcG1gNu1xI7QKLcTC5j0l
t4prrbk7iqWX5f1N+40uraKd0v0YApnClL6dlDStLWQQ72lFFLGCu6Y6GU6+JwyQIqBepRoaJBcg
A6+p+EmjyXYcPAvxysUNtLxhTgMFTITrQt5OFIqrB0gpHQHWxwTe3XzFtFY60G2GLNIw9pJD1MP5
vQ/A17lpT9COjGx2wdN6g9LkKHBBH9qg3V0OkHpjp3qtrgobpTAFeK/32jl81QsilgC48IIkbInj
gi47VNFdktGr7Qeae4L6SaVBzo6hhAbIZ3tDGsUS/47zgUpRVOSIvIqmI1k6k8wOaTqlzZNlEYs0
UPEuaO4fq1fGuMM/c3rNMx+LfJ2bhAyoqLyzeK6h/ziQ4mEyitRmj15rioVQMAWw1nRDPN/EHzYC
WACNlXsx4C4pn+lJNdJUNgadL5C6mYlYN32YgnT6MzYkWlosehds6ffmCUFjsHzZ7Ya8W+0LgfXb
RBqJ2uEqFikGR5kxFwyH1T+C4NBWpoL8lG9M8msLQwW+/pqApJXB+QhzsMbEfkBOp/2HxPWrT3Rh
VIHBKWIQjo9/5QAup9uezHId8mYZ/du5fF8cL/kgJmaqtQodcJbrdtZlA2V4el+jpjWxi4BxGNd2
L0VRHOtvuBhKyyuqBwdxXXuISkNn4Cy+lMt6K6lw81oc32ZGo0FaZxORqigS/m62kgEeSMhnpobF
xsbCqEBsC97Uw65cihdP8DJAfHC87yiIUF5GWcWA601j2tbIyAyTrdSA1tCQ3oxyojGLBOk/O3y3
Ei3NpW63o8bAr5y21yyLLMOsW/3krTQZBeu9zHsyoc4e/bQbuLlzZxpXuPNCR7//q9fF1soAiBhW
ME/M4RGq04b35Cxcmgwa9caN8VMuhq1Q1ozKYMjfmkEcvjsMV4xN7+qOSoNMMfSwmuHkwiHuujDj
iTIaAf8bEa4jRp3wVi33QVnK/58Yx2beEIvJDjzqCj5Cr5JzT59q49O1sQCxGWAddfArgRSglCDr
5NVkp3tRD/9E4QsmvFOdx+2HPF2miwW26giMGLnRkE51gaFVhSyy+okP9dtRDQyiSYunrcaTqEKX
xMoZ2Hfbxg92lV807gDkMNMvW9Kyk4LmRf4JywWfcxxB9q1oiQCv16GKNRYD23Au62U+RgWtetQG
kaV63FqWRt/W0Gan/z8lJfxTSlpDpBEbIStFUoQ+i3eIRzqjUx67XyTX9vU1cx8hGOa0sgXzVVyd
YqRD60fdFyaHya0LEIDboGaDX+j4+lYtQBS+OircL1+sIg+jurXmgb+DpFukOQYThjSFcm/jwePO
fq4glhENYikTiP9yRtqY6etpe2Lqmta/JzY08yNk8QgYGB+aRElII7UGq1TCy/s2iYgdjSmL5d8Y
Y1qgBihW0bxCy8GcA1sNKglp6wA4ndKHj531m+aYv9yJ2ZmFWFdeAPzgvmj3f8B5LEPPPXGgFOfq
+vVvxM9NGSLLao/HLv7yhP71aQUV8ELmvWUN6uwq55VVuPFW2Fr3cT9KNYR/MaD/jzJhd7665hDI
J/x4zhUxmMbPTuoLspQ1d36viqsvRRX+i+sQZOtDKRrcboTsqY7/vEiO5768c3Rfv/U1P2x7YfnH
LcTRdilzlIXAVsR6yegsg7XGrcG8AQaCiQF4M7oT3Ya0veqFamnYRCBeKfRzs+wnQq1jACYEuh+z
rzeg3ReTFfTpoKPLt/175xSctOLt77cpA7WbCiM0vTK7+eEb25U1ZAsYEhTqxw5v4ggQngukgDO9
Z3RiFHr25DdGTVTJgiQQZvnQayWIPJLOTqiBI3GS8ba/ewmjXH8WSHyx4NHinhgNkzUAYnhQz6OI
iAkAQLRtpxUPdlod1XRr0WyNo2jr9LEbgI4uf7iScjDwJw+v7qkDwk06y262ESw3MvIE/2fJDUcB
s+JL9NpIvyhRDkKDaHbJzZCTVbR4LDavNnOiTWFfYT1FTcqtEhWKOxWg3ANXT/pzRY4DzZQUtXgb
j4/EJhHWR1zlRTHsaWXtBUahUqJbUcGDSpyFZ+FrqD3q4YmI2PNb1RkNW8n4cxKsqAkBkXg/+kpl
W4O090CTagwx92nzM/YfZXY/FrhDtXUrF/yU8HGi7l0NMQp8jnjRc9fYYsI65BXevXyJOkwII4Xo
eEUiOwzy2BS6+GM5KPuwg4bnf/qAsg/h3X4emL8HZoeA8BvaqQgmKyR6ae03S4iw3Zzh1eue936c
Gu+eAWgi6Fc0GetxZO91onBgK/CD3sdwEIvz7UsOwuIFmZtGZn+7RMaYRzKI/0PR11PlRLMV0hcS
lWQ4IUcgH/A/0jNT+o4Lw3qd0IrJiaLJQtLE7V5mclfbZ5wfDNsJsDfn8TRXnn/Cv8sUADHST58f
kuCnq4r2Q2rMx+8YrYJtLn1AYVpqkv7ifBThGVOUnXN2DXmtU/haF+AzQ4sj9/fCfi+7jhT0yP9h
YRZNzR3sHrGAz5lb/Fa+QNTXammuPjmfGRk1doLsjioUVGcpu+rneOrQg+DCEXmLAZ7NfKhm/6b9
K4wQqoFtXa7w1nyHxt/CQMsnuVgXqzrA1CJqxSPXjGkPYBAWmUnFhJ14UsXb+TEA0I+NtJHyX8+C
3t9QAAYqF76funC0ewMpMnfRM9+WukGoUsoHWWoNFTDzHzGxY46JrGlg2Kc+xWpDsT2Sutg3/wVA
D0Zu/0iIBXejj4uUPs30UC61uElk1lZQw5XcqbJw7sFVlSLsdRB66YHwUwfgw+qaLVre5d8qx6Xm
MVzAIYAg3JBCYwimN82eVZ1BxGYZbW1er6z+f3dAvn+TJs6OG4hQAzMIpUqKpe5XlI0Hz8tkzqn0
+Nn8mKrVUlY1AAlnl0R6IWCLwyF+cxF05MIfSa2r0NDDHOPm5tp9wNEtgDDrY50qRMcHQTwhOoBA
Xs7ltrLBrmLWUj5bjKoHPLp5iNO2l8a2OTGWwww8PvQPedMSJbUAbQNLlO+I6zZjRC4JxaFhQIaV
4lWd9JgOasYvWZ9sGtW2QOeIvyarVjJHVtND7fguov3x+HW/ahw7L+z3M1sUqQQRdpj4tl7OzN0u
njfrkfo5vW3tV6b+9WpY4zRC5SZNMJsM6A6Ym+gtUYORqP13ZdXdjvZQ4FAbEmYCHtVLDiA5X1Xp
kAwjszkRSJAEa7BhCbLd8SAtm9R9r+700B+04m3m4Jw9qT4/sVtajeQdJGyrTUys40p9DPOj5b8D
eJGKNj72h/eUsOATrdo5zuza8oeIc8GRWLXlZbbBNWLrLQ0kqwoo1MylH+ubKr4DMioPseB27qG7
7ek3RwuQhQu7RsvOqH51EOv4uoeCUrkyG4xTUb3br6hQJ3Ph+U4Tsk+LV4iV5scE9Tt5lOgTB1+X
dTOcmtL3dHDv6rXsbeT54QyZ2sR+kZBUeO/UxTByC6vJLb0opHSgIud7F6NBGc1B90G0qeMYTkRj
Kj9K4Wiso4wLpMWbsAoeBGMNw2Qx5bejtQeDeS8d0iQgsT2X35hZtsPbb/dBrgAytIJSKVnin5hj
OBbqWEgpiCtUOse9F9Gh/xViHgvL52j140KmTAM06zmwu7hQwPPoUNfHOsIDZqNwaLQCqURHZje3
0uqVrBzPhCvNBmhP/F8ROlIE2Goe6aaPQKicWktIm1ugUXhnFCzc9AgftEXjpCa8NqbV2oY8IeBx
SXdB8WD1RXAtqS2hQ9h94tH6rWdzhKmuq734CETcbzaGL5l3gEhzAf1rtKZSw+dGa2eRBnYAu57z
pN8P0oSPcanuAcfdzi4XwJ+Xk3MCYiYi+pw0hTD7SV1u556sxvERk36hbGRGceUmeA5Ss4Dxj40f
O60ohlJ2zb4WwqPM2MaULnyU0HzC5hEo4qH0zBhDG2LxzlL9izoMAEZzT+IsuI3Ca4JXqAOw0SOs
fNh5SAvs41jp71PmILr2tb8UoiNbme4Qfj87Z31p7bd4KyONlYKq4BYoHxcYQ7PcGDXnhQBts3S3
KU3Nyx+sBqKsLYTi3Asa0kwZwjl5b+bADoDlWA6lSY/s35oHUwT8sOM9bfDML8TB18einWHiSXkE
DdiekQCtdWVMQt/P80bpyQikkiqXGB0JQ+3DDZR2oCAcFvff4X5oJb0BAKXGTmU3M248Du6pN7rJ
MmBh6SMMXSn0EUupnuYUEfa0nRRbPn5B3fyUDF9CIs/fjPUN5vRFgcWTllZFI4G7hBwYKg1V4f59
qtH1tMAFM4gTg23+CfZT/Qjzcn6Ly3yk87L32HoZ1CvAJ/00G1q2oW2N0ty7KTthWGfAxsAZOWMv
bwlgTtZmxEOvohZn9iKWMtHpMcOGOK8cOkML/HvnUiZdFAWk1pw8Uiuha3wYAFNc/VmPADrnyoJI
VtGJg7xvBYXizvYlj+QVCXUXSCgdZRHueI8919/qdTactI4hBpX8BKXb3EzPPO0Zx5ro1OSlX4af
/FWoZbk/AiAlE1CvDk7gjrvQoc9E43XnXR6Z6LFIbhEAnL3KRSTF91UCmKJLqcBcWS59vCEV0MOH
QiDi12RrQZtvUyPOZIys2BITDk8SNrEX2ziONkt8lkte6qHvb231YfiZ4kqB7YVGFuPyRN2QF/3E
4DLwBIwJt7Z+zVZyhm0ByqX+zU8KRuE6GRZJ14Xs2nsevyrGqCfwwsPUDgZMGcAigP8O354NcxQb
KQ98jneSU2Lef7gj4g5p+Y3hzgu25wwVIQcQSf/rDM2qLK8fCwGUkBgtzuX225WjzjJPJDqgdr5Q
LJlh5BIvC2szTw1qMczsGET0nf8JcZMD0gTQGa1WNFUZ8ihS16DkwexpC0MGypBvhAMN7/0pv3BJ
/z+nMmWX+Cs/1TZqr4+zo4W+JzISlNEOF68NL92Ua4Z8DHKLo5+5PzQrH6h6hXI9+dVffo0095aQ
pr5ihA4OTtSl1YG7w8x2QQqnQ0Q9HxqDJ76THjZaywujSK7MgS6fvOvsP0czWDq6NiPlWUbd/oWH
tOHeUTTCgKxflGFEd2QV6wvfV5KHiZPuNyCfJmRGJOlBHh9aUc8RROr0e6caqyfF4W58N/ZSRb06
OE5+dMUeY5WS9WrllRdReDiLZnYO8JmwD11aQqcxv21iAYTiqI+AWfyhZqe0Jhl1/0nbDwCTd90L
hj1aGs6pCPbje0SyVEr+Mr5VwdjQLRyl4H5StDZ8I9Y3+UZbqtZVn4T/K8oHbigr6qqN8BGdmPiQ
q+ZAZGLkJfI7o3/4BwdaHpiGR+F7LWfCO7TQgj3O1xvZ2eQnTyIP+DE8gxOF3dbWjsp20iOBPc6U
uKaGrFtpV5qrVEa76e0YT++udRuJgmtOyfyB5n0AJqXIMjEsxfngMErCX0P4O+UbKSaKCqMnrHHE
20Dw5vqezr+XXTU18pHlnwJljaBqyyLEOUAkvAF9mTS78eFJz9gzAxYHEDm1dAfYxtwoQXdslHJv
WeylGzspnloaCGr/A/0HU++vCZntYQlmENeQ3StHgolfFI6NMsz2zgkQDOyQrqTp13VaIWDQdfO5
vmGx6OOazIfu/ae/yjNe24MANSIPkSZLYIs6QHKn4CF8ESSMLjVtUYLI7kG5h/5XiYaip3nVjUr0
fbwLJk9rZ8q2TYDtoAvJ7tpNc0oNb91WSCV8PoLeLQAu8OqQ+t93Qj9MTjl9ZRvJFLRxR4h3A50g
tti5UVfJNT9DNlOrqJD6kyB+Bq1v0RJdofdhpm1yCq4h6efWnEltzSHzyNHBufKkzJCfReO9CVcE
8pWfJ42vD8mhazdKOOC9484A3kuYxl0FkoPBh7YNqj+yxXiR7PPpssnEBwSeYti6snqEoxB6lIEF
BbPMd2WqSX4eZkg0jRwA4w5J52JYDx+YW+LLO52L9n9vHgobll5LY/cFElz+ggxtW0hPeekEMnNI
NKcqQHSmZdo6Q5muLfek50zzOvJf3DmiabMEDkNfqkhqen0DC4J/O8ha70z+scIUvj+MWLpp8gjX
AEZCiGfJgF/o3Z4784YuX3CQRzJ8ZCXgM3k6WIOYBYf9XTbBgMhrQ3Fs/yxnkTRCccb5qKGpqOUV
KHZrg6RRtL8PZGQAiDut+xShLu6tWqqam0fwzlZl2msvjzPJ2UhOaMRFkrqDwVSrAE2AH8TrcvT6
kvgbCtXBihnR1yEQpdwMIM7/wXCNgGUTi0TIvvZtYe6c5uu9cLvUGLNLZVui3LJ0LkmxMkJ+8Gpe
orklVgSe9mSudGZx4dXkGrDLdS/uYUKe17uX7Fpx2A7aZL01qFMLQFdT5vuul87c6OI/u2moOfCG
3gE0e+GrzBU3qGpdK0oKaOr9Xx67fFhlLgjZ/17xDR1yhYlc4S40njOxBOxbPO4FZUo410nxuNjY
lLDtvlYwIsBvDY8TRtiEcdB0yO10k6gEsqsmU99KV5+NVoARsPz/vWVCKAgVjXQ4M2sTXJ0kyCqC
6lVtv2TxVP907n1m2/BpmFkFL+vB/78BQOZdhHCbnOdq80w1pBwHuBzM3HC57RZkGwgsoDevTX3f
DP4PdA5yJ07xMyCDG40M5SrLrvLf+yz0v/OrrTjLiDmx3nLDYVEV0Qr+UmJyq3CZrp+R/gFGMdxf
W7bPo05UjSZBYT9aze/NlMt/9p/4h54TV7ZGT1dg6DYmuKG0Q9Uc8qb+NJ/V9DJjPGw/8pRbHpEQ
cDRtZEUkOiQzmsJkLn8Cs5+4oirIbNucFSfYjqhQJqZaKDOYIr5z+6cKsgAMFWmlbn8SAW78nZZr
pNswWCHVk2sMFV4Tnpdf9nsrUvJ2wu8LxrnvB6YrIe9DXrG+ohYiKFdJXnItoGytxBsfO945UGlD
HOqWscZfJmdj9zcPY7qnavCyIfWUGuvW6611Ph3c1eaWEijvI78+/XUn1t/OyS8cqz8KIGwn9kaL
P7QKMBWTN5X8Clnw5TOTbm06eOQF1I/liYQKk9FWKmTM2ZI588igLd9m5c7JzgQKnq9bzLR7RXvw
pN1UnN0RiRdqpqzuBAEH4caMA3IkzG+408s1y9F5wh4nrt9GnZBbqm2dW7ms+DRDoGhmaS286XgM
+2lUuP/ucIQg+b72fHBg2Lb6A0SvHHuIyDxKH82Lz3QP8vyWYi2q9HhAdIANvF/w9qBmqUMac0RE
tlevnuz9hvxgGPFN+cY44sDMkEpBAOQfpR9YXkrVa/Qbu1aguU4NvUN2DgQpT/zBxK1VzWHxoj3U
HUEv2pP8cBntS7dnYQq3MV0FNxJfQDQ5TpxFoa8YvKDr+v1L9d3UW0YZg+fdATNW5I6BvXOEyQKt
sR+wAy1xm9x7+zg8tKiNemEyriEqCqv7Psap+ovSW2kZtkuGpSmnLtybzr6w21NO2m02hLPF7TPE
6M4NaSxEJ4Gv51Yi+YS3U0VLulDmmYEDXZcqDjhiJ6ezj03QSe+c40G6VMvFOLui2fztA6DCkjcS
l+tZPLiKIqFBcQyvf17SKmYRjjdp8WPCZpQbt+WHsW6O+xy++emFO0DkgcoSmqh/urVNBtEcEwwr
58J2kdjs9Bb4NDDyRRNSPReNpP6p04QKpTZ8CAzr2WsHGX4x3pC3WBf/zZ2yqsmPWiQ5dPXm44Ha
Dvjop/lOZFR12L7dfOf75viYrND/mFiwCbQzakZHzXTdEcWXS1tij9vV4raWS6RgjY6AJkSBd2Sa
jcIwDPmkHl0pPQe+wsqw3DvtlUd9ekUT5Vrbh7de6wJW28hDsBjBkLXmMgyw2defqUullrTbx1KT
23+Sgz0VeRjR0aAxa9Dvi54OA7gzYi3aHJ7YcgZ6DVJilqCfIYnUjRd7nyGQ0puC3TusYqWZi2r8
csTC6fCH5GtjT/UUA2zX6TytvkQgnerq0/Qwxa0ED0ORe5OQYC5FT5mSook62hzZ4/l0vMQCOlnq
Yz7RRTfntIS5vukRFXaO1RhJkpQeBRXbySKq4H6cYEMmELhe4p9jaQlVaHTo+3V+d7wOaURx+/gW
LknDs4pvh/9Y5TNnPyelFPjFCObm3xRQ5uozebDeqKE08Z5hyxymuOTditkHc6qD/mWcfxA+02Bd
a32WNivA6k7aDZkNSFeV0Xziw8zq7PXuWWeAu6tLKhnDciEdBoDHQHO5DJJRoqIuwcoMp/hN8NBA
YYLTbzr5MHvA3TpJSkYqPoex73SybfOLtdpBOllt7JlDP/4BKZbbifNA5TeQDsiJNhLReMqToonY
O60zvBNLat6U/6MGgmDEfxlFuMD7ppHgNUkAl1RUjRTj6m9Qhq/SArUVXYl07C2BO2eOp5jf50Od
puyqeDV2JuCFaE+B9ew/lxw3ZNKKP8v+qodBqqrFvLCsACrP8QsB1/4a6SEh7BnuMi1+Tno8JIbc
+hszFAhC1i6BNf0r31BShA4ILc+77X3rVn0ZZRBTwpP8GuuN3Arm7oXc0jN+09MvKb1DO+HZbCsq
wsC2sZo/vnaL7U8HKUlD/ee5xSJefIEPdim2BS5RmeoC6E8cRa40d3xTZznQk0cJ8i6RV20Iy75E
sV4bvWH33dU1piYTTIw9f1VLZWFEqaJPU0VnHGRwNzUGXQEPk++ROhSsuNe19JBzsLCPmYGE5XfL
i8RytaTlaD5eiUSpisqUwi2vZIs0yOolcJ/yKqNwWapo+phRDziDS0JtRI09KIe6TQSqraMGvmPF
ay6k3NG2R4TqxputIKSKC0CCUffFIFa7S/ipaZDo9WHrdQtSHy0WdSIY35HUVqvsNlzkIj0tJWK6
FR23g9YAzNPBLe57ag6wmLogpj8JTILt3bZa5Lc0SLhpqyitBZBHFPqvdKLHkEXC02wnfztzKAmD
TgotxnPopOmrbwf3EDUbnj1Ma4ncf08JExwIhhJvuQtNSg6CFqit+lw6BoLF6/2Akq5MpXq9rX4P
REasWVQyn0wvnt1AucO0H06svFBhlBGLa4/CgSar2xOV+1ktrbaCnDpKGzYNMlZmFH1SUv7Y5kJv
HoNAIGOy11pD49whg5IGIBRR91ON5luGTA+iakFFtPFHvftmnvGIJQNjNMUnJLx7C5C78N3ZNKlg
433kkoxzugQjkhHG05XhUND0T1jtQ7vf4rgdTxhFCyu3oAOJyY9lDzqLv06tc7cpso+8Z6OCGm8M
BJovOcRlTi0Y/SOObRcLLCbZbGcCFz4oA5TUaf4sMk1tKNsu6O9E1DmrtxhusYT9/Q3mzojqymWA
O6FkLkykbLtUN+16tMX9NgB14TXDknHXu4SVFG1J8HGzkgkCa5IJ2L00m8AzEtI1WXi/ZAqsYez6
cSxGCVCIiwvnPcTTMb+1uN9RSN1ZcMZfjTKBCPUs0mqjRwPNKpatyibPek88kZfj4OWsikrqCtsD
UjmQeJM0fhjneutvbkmtjqemCDxwqQuG4jtWnQ0k0OTq0A+QykQVGJFVk8kwhayIX4oZdcTOnfhN
VUSr+HMz6JMqa2GvGpxlvbHJ1kKopZvGpc6ZY4YeH1ubZs1vZGcXUy+b/wRVkNhLRZoxoTFh+qgp
9leWI4DsuVRuxbbiwPuNPAl/gTK3hc9sdmT9QuGyjy8G9uSnwrnpterqvKzwogSIO9IBVTwMEjn8
lSeNeKWUXmj0ws9Y6uAcNSoLEoTDPgAfweFO73Vq/gtHPL+32Q+qM9oL1AYv3MyUMbamCS3QN5gr
j721nnHnC/IJtDWfA179zFu2BDDj4dcQQZ7a8SNyYp6vYs/Z3fzg86/c1GlmDXIj1eBeeIB8z8tO
eCjk/tVHq3+lTtOKPE0rr4Qiq2mWwzDdQtztxhSU0tm0PyPMIUmT7/oyX7Qev6svUTgnUcgu3Oou
858IduFNPWhl2tQpZ20oJ+1cpWlHIYs3Hxo0VwcIYYJ94rGJtvpCVBkd3iTJAES0SCJGgTsDmQmX
gnH7wTkAxaTxnrwgwIeojmrPTg2trgh8F1KGq1xs+igxfmDRhTFQ8CxpIx/kxHFFj0oluY08sQ+o
FmCAJnSMzgQKdH/8MmMyR4G+tauZdU9BkXjjjqMDX/aPuGUDAYu6HaynBOYzuo7Yvv13+d5skgpm
nlPv1y72Ej7fzQ6QJhKdwAOLsFiVjH6S1CnFdaRikpHCwmeTksx+krAIDMlerN7p/ujWkUmoT1ts
F5xL0hkZMVhExWLsvQ8s/Lho006+1Z1atwYqqrsAKHPTgjJYTxCcCuwP8zNQuhmOhb3+SuGa4UkP
IGp5QvrOLe1GHzSVEo+T/v2tE63swoSJBLvNJ/bfxTdgja+VgMc12m/2HePwKvcUPN+yw+vtLdN9
njZ9pQ2g8AO2dBq28BRSOge7IEcjtmZ9HjIuArqhFWGHbvJLnofIuGG02+U+K6ajcSOB9iSqoEtp
oNjRAthJXXkBxeI+1rFGspxF4wNyvcoNsMHjMHydOiaQqM31WuyyqXonEi2HjEkNYBCEF4uu5czW
mqg5H5I/3mTVIC8M0Wirxj055LDTqajm4ypUp/S+wR2m5v5a3SmMJyFqf7sLiZXumgvPAR6IYLIZ
XkS3jTf4Mujqgc2nDT6dg7N9XpbXFjIbUBegUf7IAzcbPkqurwJEcgqDygM5zLQEi10G9bl3tecN
XtHZ8KBoETSLIPERN7s9XhANKphp8oiWFQodvBVAgbwsqHKMwNN8qtCMW4FKf1EVthWqOFvRgewU
B1P9C8CWlyG7n12kYXuLQdHcYGBjMsHuTR+tnLFpJ2ywNmZIlPAadabms8i7SrLeyJOlMSIrPhFj
RWy3YKKUQSRhAqNlJ5eQTshE6jhB6dAWU0LA0/7tY7mmszNHOXRYhJMtoGN+AxRUjct9Ri0Ir5VN
XoNYK3MG96vpO7neJCoIRrWDgpyVSF9BoqUTBFJxJWK85W0Au4Tjgx2fduYPa9G+IzGI9h1bKyyX
g18QHzTBaJrCSw/1weLSlv2ofCkZ62MsbNM5FQmBUs0k6LwdHKSuQc/4eqjKTTlAayIqZSB9MiwU
1pGpyH7pRgVZ93kb/GpJQuGHxwx5qu3Otwt2HA6mSAto7cXE0KQ1oOlgcZFp/9qHcPE6Ps+uuuld
K6/ZRhTnjQxichM+DqWcHTBiHszaVFQAfvlFzSznA7r0obAkd4dEuz4v2hk58HY/f6kKpgNf9Str
nIq7CMXuWT5h8dZLVP4JnZA6ZIi1+SCGpRPtjxxYz+AZ+Y+Zb1AWwCvAC5T0znk6ax0BFZDHin8L
bCySeyf9qnxTH1gIlxkUxggh8SxD6oaxQz8LR4PphJPY4ndJUXbS5t6ZfTGSR81J4dpoAVk1NLnu
ZHqZaO6aRuSAGW8Hdx3yp6zX3KUDH9qozku3GjMrCJEYZBlzg/Wv7iFxVhb7HG1Jn0HtkmvTu21D
6za8IRaTiHVyB4MOPcyQ/oEYG+xBXvhQZYnpu9h92AKcc7qAPFgi8TdOADRs6uHuPtDM3eldcyeS
dZ/yT4j+faDqU5EtJNPYmsh3P0DyDvtLq65W0Tng8dukhi6gvUWA+cwHzOTV8WEVUasUOiNa5wEt
dQdiWMndbxqGHC320dhgLKogRjWJyyHRafqbvpR0DujKREluebqWP9qPQKi2dF4trCbhOuft2/Xb
yve7ic03bYEJA3pKQIfn6rme6bLdKpSAZpI8IaQLuEdIQAG8EAM1QlCOqAUPSYTWi0UqUwRlaq/Q
CaKJAAsiH1OhQKZiEZOX4fpwoEafaMuaIV1npXnkv/oAZ3JGVRsZiZdXlFn03pgbNh2dRacluXIl
pPzKfXl8Mv0yBz2E17Fct7Ydaoj0XNm263YJYFk4AFebxriIDFPnHbWpG7E+2KdLQzQk0zSZdrIp
yNTn3HbGe8Q36ag2FA70iIr90Ec2xDiO0XzN1Ikko/PVFgpv9znte2KjD4MrYCF6bhvMnfRZ3sfx
bOAwMdi6w9VT2KUKAkdUPpmxISBH65qQ2hphqLaRutoHKhLwW2p2PWXE373q81AVGddwpstFzCTd
VdCj0wgenI1IOGRp2UivjPF9ittL0XqfDbk+voP5/wWztAd5E2c12q+oDcH9YjK28/CEwmJuH4uR
PTj8EmfRFUgTsJerl+t3vPrshE4XD5G/CvBegBD3dqH7Mon2OUYTzUgd9QAilFvPVaTF35YVXuPN
9kpEPqtdhPZFF5omPhZAZg++zqZ+N5Dlizxz79jpg7r+G3mi3XDNG97aEPZknz1aP7McOuh2aqk5
HVrVlalz3Qwm5feqrhiuXJGAjui7swMjvo/cJKICV/b3G24IYOrhVU/B7nLbSKlorp67vsmEnw+e
GMo5F4mpF6KFRVeMaPi452P5Cx/Hj23sSPntveXzNCTwJKLV+dTG5oteIkyKJ9iUEkwARiCXye59
usIWu+KebPjDB3kKKQKh4coAgFG+bYCR32nsKa2vQltJEW6Yq+c/94DdXiHggR9WF+Q13AaeSNtP
1U1MIdjJjLKSV1UOqok61gqT2t3ScFA2dTZNXZLr+k4a03ae4PjQZ7wN1Xh5OI+XnE8FZL+472g+
6JZQkf5J1JXVOiEmNyTO+Q9KB6Rszu71BUiVxnB//ndq03woJuE8PGRZhbA94xDIAyXfkHL/MrxL
mVxvChjwJfW0lBtOtE2BeSxVlemhjHm90YJiyT/Cv0VwpAbUkYdUcWBF7cOPoKMEeCYxcMM00Nqa
nEF0QzFxDfKET7cv18lqDq63iAIX47Oa9xYWAy4OhbqcYeRkCZqcPQ8pbiqCeHEP0ZhDmfZcJyTk
VmiWUTNIhbqq5infqG6v4YiO7EgWE/vNItQBxITtOCmTDKpJLDvNjUHi0WmNHf3CCvQzP0HsOmP6
Q+Xc/LQ9cMQpO+NBBZoi/pI6XnptDllo3IKmKrkM8N0lsvXWf1r0QIoGJrtWbXxRDCQ77rIXS6dG
adDdG6cZEXQxfU9tb0oZ5+G55BHZKMiFvIpvlGlQkCsd20ZSDIMIC67ZswIialTsBEm0G7cXOWnu
XcMjGLJmnRYKhOxHC+sARA4+i+OqugYWBfUp/7/YugCgGg0eiZv6oDPhdCv5q/5EvCOGU6SOTPLl
JdIRAp8nQ2SQKQCS8aQtJsPcaqvJMLQyUpdPq/pITHxv2HwGlSqtt6IQ0qqgHTOLZDloV96whZ9X
3DUjRHD6EVi5xQ8wvtjD6FFZsDRZJEca4E5HTZ+PRC7I01JjQqCQ70+53AuEhYSB9X4hvV8Sj+HD
5mxKMeVeBgOdUNnwA/NfLEDbcXSAXVP0ICQxPtyMDOFLG+xQfv68g0K7uPqs+EylLTdcUYheExwX
8UQzHBE/mVN+KMZ0iDlEpqLVgk54v7f0gHOqce3VTF/ld/KG0Ka+NQRk8BzsycXkSIR78W8H/EhM
Ifn9gmqG0ic1VLMFwghJuOARLhLnGBVV43+wak8cJZHvW/il+gkKAIK03AhhJLEpqltZQ9mofdCv
9iAjBfUS2nc2vWWHMGtyzpwfwVX7KJ499hoBuNbDraZhXQX2UnGhA3kftQMf9K8yIlKAfcCWxdQR
oj+MY1PAIVLqcUjq9N8K7P/xqS4aAstrn8ntFgGHP4WSTDZEsS1gytj3n5JPIAKQJoU9Q2cy8QOf
6FmvxPECkNKoFHSdlfeT+qLXDiUwnnx8J7Fzt6+6qSD/z1ybHk96m1cyj674N62K9q2HlTE24wir
fob6iNyCSU2rp8PWfZCl2r4IAHr9asYEN6ZUN2kPfnedFc/gda/xOl5p0YFDMiE0Ha/PoY/Gkect
HR5ZpANl9om2nJc4v1gpympZaCd75bYIsqXqG+mkwvtOg8t4AGt33Ft/6bCOJLwaLwIxzxJ5Bc3w
9+kiNwTndmbedyz9KF3+mtOg+6xnf/SfNv/7w+49nRRnaW/z/pB1I1c4FQeiGmI99yCV15CxyO0I
FL+pvwIzifY/yVktjj8PfjrVPYG+W/laml6uSjc5N5+k7pg9R3zCB6TS9BvsO6S45I1RkEguQ0FA
Dz0xwRUaEehT3WMJS8cLdu7FdIZLTSs3PK2sVC5siir7l+tVmA27Zp42cAUnNM7NFspvdj6rP+5R
6m1RfVr8hDj/Oqzc76aQR176SELkmxHvu3/dnhOsPvBdyy3/R0GXXCggZF/Q4HPmMz46EoIBXGsn
dQhwVR/x/UXKP7EdYRG2+T+mf0QuLxy2rJuo7ulPtJv8ckhvIAIFDLjU41fft6vNR7gKeW5HM1cD
nPgvaTmZ1WaWUNEws20BnaLh80HaJ2eAYsPesxq4NOD6IyEdROZU944Yu4r9yBaYijEK4ASlagoB
Xv7aFXLsogiLQLhZHjgayLnZj3GuIevaQfxagbQBNW4T0g7cyh885mTkssrtNZp2Rr4XGvPmbkCH
vpAdZxw9xySmEYnb6EA9ysJqWP60QwcBH69Zr6PzIwjkhZ5hlLZrTaLii7zrBn0mXMB2jpUxnZYe
DEpXDB9fd3NdbvbW9dSY+bLblnbowYUNqXJuD6CNP+nNC5zJAyHRKM5l73bAFYu35phaARTAVyqH
lPbK152EDye37iuj18YZTFUT95E0jaQ4+FHwDF/rCL6ftfqGNkajTOef3ARBYyTbxX2E56PIGBwW
3Dq/ubFDEKiq37EreBCTb1wGQfSGi3l3BgRjlcg/ll2z+bn8LS7Gi41f10cjcEIdqA7satby5rld
6R9tY7PntF/QAJPulcbk8J+Ia8Z5czSH/ofKSqqdouB9BeGosBiApgdDc+Fd08qTnDPfI7xcbscW
gHaiBRxBRXX1gOjP4c/F7+3oid9vMZQndMbpTWQOhH+61vyAiCSmlIagiOsKuNVSStBCmx3kHf14
588OR9MvOWKtIeNO6a1U5ebyXO2Yd+Hb0JSONtkyPic8d+96/PGMfLTphQfpZY4xHgB1XGiPdp5K
tzHheugRgcAqjo8AWJa2sqre7s/2HERqGRoMcBW/eRGsBGk8iosfC8KC9evBnciEVH3MqtYoDTuh
iJH4KycWe6gTg/d0GWmiaJVe2ukyKl/3/ip9kYtZ8b0giT71EMWbbhgnyLCQ3Nu/2nn62CNykt1J
RThfb0bduVJdjwMjge1amanvP+8xpHMOdeQJkP2WsPh8H9wZFvivZzT8SQ/8TpkZ1oUpJXZpJI2E
0HHVGEBAKQu3oe4TH5k+ERYe+MKs82neuAmwmI+eU7g/QGMaNgziUkdeERjFoC89pHze1AJlCHpB
qr19Z/+yEUVhzG9F+lDjHYa4MoLj00ETGhYTdvbpVEOSA4zOiNtrg7YmAYJpMNraLNrD0NVOsS1j
sLr3SWa0x75W8Ii+hO875JbRAdXPoyyeFmn5CsdgoOeqzPzQ3blDwv6vkuVmri60tTPPwx4zb8NX
UFE+tvPkIFLeyFqX7yYFevOhiJUVpfz8NF8pGhGDbJqHRDnd+ODhBi6ov+Mg40q5lQpPgA1KnsZh
Wiw1HvSp9RKyfDl0x1e8bRJm953KcYgrzn90GdFuvl2lqNgGfws9anmveur3ZZ5VQaLAcs6w3mx5
UEn1aHehTCEkHUg45ireoiTbLICxJYbLWKYGYIYB7zZSJwX7hM1rnxxJHG5REWBjX5kVvhwB2lJT
1A/Tb/CYbvE8ezC+eUYhb+HG7dmapW8Ig1pEkwhVtcmzMLyH2Pd2F2Pn2h7NDJtDCAv/B8UipFVD
8eZPQ8qn1SNm4Pojk959tBXm8wmFLJvQYskDBw5OdTrSsg/0SnYRG2pbOlNL3spcUzWHSS7dtymi
7QkT2DUpCqGmnl4dm2egScnRPVIOTv3r7ZV2cf3MT3pVmTeQHD7JAMyOLOkF3lK57FAwcXg3ddis
oIw2hRj7u9jM+Z+mK4FDxEvJztXGeCsE55/Y7PD/iglLY59BROi7lr/AXjITLMpodexyBHetsOqi
iGvLlNkXqfsOQ4I/3eu2F6MDBhucRCsUNQg57TxxunJLdfd2dyUll0JCsTddwhoEQu8Umw44IMRq
gXqxXZwgzRidg2jOVILNM6NfFgtVQhuXObGpwLDFQeGUjhYhH95N5cNV7m8+UrMrxzRsVuyevwwT
rRsmqpzqkIxeY5Qfe80XvnmaBvJtuVVHLvuk4RJEh0lgL7YXkQSG2RDw5OO7N4N+7Q+yTXvZBX7D
+eTcraYk2Jff7DjE9GIYGTgQGzyvt0ysh+ZPnAETAegIj1vyzlR3519dk8AkP8oUwCEpOpDeJMqT
GL3K9QNh8SUYE4zDCzFe39hLHjUt0oZVfbyAr1Eku+qgbDq0w0Ab9eLojOb/90Vhu5AQr2NvyCDB
bx1JEp1bdaj+86L9Y1jjxqf2UL3ENbvlvDO1cTxJ+quDm+PCZlOks+1XtIPeq18yelpmrBjPVKdw
se473Jd661gzfie7wEFvYa8DzsDpSLLA6WpfOMvERB+gjgyUnxFTctOqcOKZt3BRjaj4I3GQWLJ0
fyeQ0ehSiTGaH+G4gO/MgD75uHHxquNsI9k8mRrF/A72XnhY8FVK+1gCrOggd1QjAFRXhRx4PvMN
tlSX7oAENn+QSfYlpXuzCAt3BteivPqB+t49BDCT4JaIigHHnO8cV/I22s1ZmVFA0DedkEm8+RSW
yAry44dmjNMhtEbhFweyBHBLJbaGbddiUZFJ+QywYZzM5MaAMqaa5OP4ccBRf8N+U5+bBJLi4xrp
bM0MW8KAqOVwkcmCWU6N2Pvi1jw1Fr6eEBEf945rXK836uS0FotRl8FZMG1aYgXIPJe8BbTOZ2nh
u2ZV5CzIVvPDvrSCdSVu51Nl128iiyt9HicszrwIiLGNC+Z0eVs2r5ReG+1hJ5KUdLFu7yDnHmtv
PYfqlA2BXx6a4DIotGKVJ0jXqllHjgMcRWllej7iQm+3aQKiUWCf1CdCKz2dx+f9PWE04Xn/zi5e
e1yiPVH4YAXKv28T385vN3jmmfZln16WNj8wc7MFb+7vFIjazOjKhblEgrfKUGzYSrvhvOX2cVFp
/aMWEX069yUdoLQfklCJxSe1QR8PgN3kWr++clpBN7bNTHHZhlGjtdr2g4YLxmayajcrbNqOBFFO
7jro71iKv3IIHS44NEBGQj+Be4ZRE0BTQoedO5jPPJGKixDG3u7z9qgmqKJEJGQQA+YK9+7FpNPa
QzCqQKmlyXjppwkwlUsd+mzBtg+oo1d3fCrz0VK9m2pMtQgqabMRrMBQ2wVFDc0NZ66+LYPkc7T5
LuggONaJcuTJPX7wx51FiHWHBD4ALeU1v7vJjaqlXvif+80P+DRnEYzwyk+mEFnqEPbSnEsREB+x
my4y58qflJ98NJtzBWDQghnPJBPQXUymUGlf5XRGYFb3/kiCCWY8LQl/FdiKkBpo1Yg8q76IHLxg
YDthaNAHfJbXYcKYeoQ2UDmfOnslU/HZGEBIzsxmTgrQtBtfVblETK7UjPz3XL3oG9J8vt6q/JF3
d+08QA6umO/WXbk5cAFSt9Fn2JnnVTkXZffMAC88AMih/Vf7ul3hfEWI6kXd/mCV5Dx74W+14bfi
fpelOCoMjVsO90eMENsDBguxG73xkn32qBReeMAIbN0WX/B/9SpBSy0mltNQtTG+obZzt9JATxWw
zvV1P9hR1UxZuxddwYR+q6oGUiP1bnLhVMnPOYYGOZmJc6xnEZM8rgEUaUjUOntbZ3nyCJo2aQxb
l5R8sOVpVGSuQh0mhg0yP7yos2iC5oC0Onzi4o4snriD0eqCogtYZCe0S2Dh2Sl4dcHCd5/rbLEf
cibx93sL5C+PvTjcVnYrynFS3VPVE2w3KA8HgppOqno9lnuTdBa/8RTfqab6PM3EXqdi+j0TXCqS
lVwEuxGJlMfQlbKepPy4yOJ+60y9JxELDwQmFMqDm7IkNbnhQU3yid42BtYEegsTkuTfYJm11+y7
tLpSZMIfxC0FLcYrK1U5ncGKtpvoSTji/u2mO3ZYkIMWZ/JRczt9dvVoHvbPM2/j38vCSIsdvYg+
0m8KIuFo9Osy/xr6YN9MtkyOkoBFczR+3q/c9O5oQ/PdyG7Mmw132KzxI7e4lNxTRaNq5AdfBRvx
h3G0EZWLB7FiUyFcY3bHSjV/wa+Wlxxk73Z28MBx6J9RJhw/XmhRP51BT0j9K/rdAlEk0FYFI0dt
3aCN/4qgpik+6q3Z/J8K4JCnhSepF/Cg/zYvh5lx7/jA/qK1xg/2qCmV+ISEPpV2I6Ux/3abbVm5
Bj7tBHDjpslTGr4K/tCaHcPuh+nbwIKQpTUtCPeJubIgrqPMZzkWUqLceA6ej3mwDQFN3vpktdei
+IRlMU2GSCvsQlqv5im9Z+QFo7IpBq1QGwDdIEDFi5G2RPGWyv+n+BdLCmRLxzq5qWPrYxGwA67b
vgBb9nuhidFe6MK0FzcQO18i3cqlFdeL6t4/vHlB8i7i1Kf96WW7ShOF4qe0xDTXQLizFw/SuRWu
fYAG2Blu4MlrnVmQLuvdA4W1S7NxyYZtDyVnZDMWoXlucTk/6iLT9YomGBqTphPc51mtUBwPRcjb
dwZzrYpxmc2RwJRQbfkv1PNTSfGrNWrIibDsTnUwYGVzw5w1zmJcPLg8TP2ZWa1rcHrGyoBzOir9
emvr9cE1YySZ9RiDbPAYh7Ts+kwQXrsiAV2iD4qB4jSxO5SPPtPBqoPyBfSO6JrpFR4f9lOhwTwU
PYTcf9GbC7e3q4S3ilSysB1yVRS2KGqSSEQ0Vgle/j9JEaoJ66/ikclU6CA1O3HaweMqA4/HjJbq
l8XGb52CI8k7fsgq6Edc+y/NH+aJ/X6QEAyqF/awxZwHUQQV8RecLIXg0DwrrUBCZPyIBWFTzBm8
nUpupZ1ZApjwE49JMje+Q3Q0s17YNYJvIKhASQOLuekslBXzRT01GcjA3sJEoYyhvfELpzoTfNFu
uZzP5eiy1Qqv43Gby96RZGkyFbH4EaBnK98lGu7fQOgaCqFdwImjHBQ7Op4ukHSWCtGM+XP5XZ8M
F2UoLtvvu/Lo5nhG7T5wp3HinSq6MaSpXue32CIqOY8EbGVhKyVL63viaXAs8HgaSJWGKEI3vaf/
f11oNHv9ZuaiNlvoDDN+1zOSXEVtPTGKqULxPfFwP7DyjmNDjlL+AxF1eXgTO/0KmT07DlCU88ru
jaKgZSzeybFYKqxbKSrLYWNTyhdnIzDz8Ux299NtZZtxKb5y8ED6rEkEDH4Bv6HxGotS7lLJ5eOH
wfr+KNLJJmRHH8sdTLiDFSnBfDLP4R/eeBBg1o/Yz7yCWM6WJeR429tQ5qhHoktKeXhg3kWtR9w4
JRAY0zIReIB62vwoOasA6V429xNaYlcZR1E4gDDXmPamCwzlJzFCG4/VNV8jlqw7J556Fyki6koA
2POtZLT/x8uynjW361iJKu4TcRmKiABNjWj8XVsrnxNlZJb2s7sDz1GboOFOWf/dcwGXP2HDzAwk
NlNI08QpGRdRhDkRHJoUlOOV9HGf89aorXPz77jyMzcFm1uN+vZmqrfaOTiMUu/D8Dai/OVvGp8Z
Zs0YO5EF5JftKOPTvywjelyE6LHZqdVZGydDnZg9g7LElkZcc9ElqroBjkRVIEL+SP8SmofCGtb+
r82EI8cwt7irZ6QbNwVLIn8W4hrYJmeWcs3OOXEwJ7/Neh4il4sPozCZm5s2k5JTRyV6uQZTbwqc
X5CZgoNypCjMa80xR57jivfhicB5xYLstCeEKoNAljScDrXnCIBUB04C6nbKrPLol4MuX0zEl0bH
wrf6nQGIqeilDswqaEXzK5fWScwifjQ35REUUKvV1vshO0I2ODOgUS/TEhxnu09LaGdk0X6n3r/w
BWMSkWH2dRgV+EbFCS1K7ozpf2Cti0ytUiVmnLSYsC+wjJXpvJbGAC7BngPrvRU2qR8E0lfsDXT0
+6/Z3l77rG+PWYVrjfoXdUZdRUcE6P52SuXPsnFjbqdyrvRTczLJru8jwi0zEEvJ/NytwQmwqPFa
9WW67k99t2TDXmWyYsuf/gPCXqWtJ3NtlSoDceR4i8Ipz+bymE6Xo5AJ32b7auQ5nHfiIZfqGP2l
tXDTWEeH/XMw3aMdaNSGqPk9VjJN5SgQfPZjJ5oTjOQNkC+qZY19W6V8dCbrGQWNVo+ePXNOP/Wv
CIFIXEx0V4B5pdC979/2p2HD6b3N4z2p6TRpRO9SNt4FFKefQ4qD2gvnL5FzCoEchO9v7GS/m7wz
+xiMXZU5tb+mukDdNjmPiRD7aJNNg1g5HOo//WC3INfH5OsnY5tUm09U9WxMTzFduB7BwWqyW3vy
6ceWoqpM3PeVOqqXNlE+AnOC/l70gq2HtE+MwT2O2mxpWBH+D6nN1mzhMWgbO/L6Y/ZFuzp7x5JY
hvDtuNmjnZNdIzzpc38EzTJ7zqQtkqyEkL7O6MarWsf9wow2OTlLVdRtjynb1tPpxz+dkKBxqVyH
NJZOep7O4X2i2Q1ICPUq1Oo1cTarBEv4NdgNyYUgnZXfUzMyZnwesKf12VviagbJhXPC4IOtUSvw
Wrs1Uifzn4MpWWIgVlFLjxdjTtDm58X88j6midhqXV8xgcV0Rl85yJ6InryNE++blOOzFsmw3KMX
FR1gO6mHnjQHkTWHykHF5sh5ZT6pR6hOMaTvvgwxmRImEK5+UBIj0OJ3o70lg6iHNCLoe9RQRDdW
25U4PmurlihV7m1oOuAVNzkFMtiE0jxrrFSrI4g+JPRmToXprcudIOBon3nyhTCDsQsKFyiMBdv5
tik7enpIMSj0oSnSzfz2OuIbY8kJMISYc1SbvSatBohtWwmq0kkDtRSQe9zJVUAk5yh39esrXr2b
4jgjGryRSadc8TGwz4jnKIiua+SS/R952twUDlf0jl3FDunI9a85m7wY/VgxehdQfT9F+rguHcEs
UYbfR2PoUfkFPJbrAE69ih0lbFkoHNWWmlrzcgmuiXFjBLTgIyqWluTGqfm1636lPLhxokc8E6Kh
J5Xfj1xAsCrj81lz1R5K7Qlfwk7PjLqGencB/peH7m6qXbQHlPDyS1NalralBOJj78F1WyFKETBR
oSb/QIXVTDzuK1osPjAUDT/7v76a16nF0LZgSr7z5EPgGwCfQOZEYTB9IYp+aT3x2DSC7bKWZSeB
vUNYcb225FPBlvqZJ6iP4izeCPtyQYLV6ei1r/O2Ki68CgJX3lGi4Rby/fUFtl55YXU+db/ofRGb
nxm1AAOayAsDYAUl2H6QY/kNjGb33bcRnIiEbf6YIUg383CltCXmrxFD/gjsm1ICz2KAo7DD6zXD
dqai14ktFQNR9ik4BSp7IfsvKSymT4ViCp4knvybAsCcdsYsq7tsfZrRaXTeYHld59n6REBkTdPX
NFYlItuFLbba9y435pzRLpMXCMg/YApFHq7iD4zr4ai9C37RakEpdkKr2Yfu5Gp84obdH1ZBBsDK
OsUSjLPP57D1EbOq3gsCNqYGxKrqwQEakWkUr7oWv89FfDXlnW3SkVt4I5HmYJr99rdcKKeOzyTu
QG+oZfQBuO77S6Qrs5PsKF5BffH7ZN7vBPokS8xG1QSz0XV6crDaHTL4ErbkN9rGxowx+Ab6LEyj
3C1LlePdcczJ3Ho//Fj3XKNcnlZJKJ9atDjqh8ST+ZSFNmgSU6TSdhBds93ibhcwBX1Xe4ED5gdO
hJoBRluaUMYTp5OvHkfHkgd3PCI/PDcEhJqeSEkdUHpSayIdBEKSQYrnRObnBQC/UcQZWmdJPrUW
djXrIfYFXupW4VNW46N9zdAlkdfZzLPN0x7j9cjopxCaIf9/iybFzNycRxEwIW9qij3pbh8u4TM6
EqcwhksL8DM9esqNdsjyrct8IMNbx1tR5bcIQBOF5sa+Jy81g1GZWJuWYxDUyLzKDn+DvzEGMThZ
uTf3YC8Wro9XPJ2qgCnc2D1a0UF3/sQvfBXqPj6d7NcpuT/wIfgUN3awUCkh14EgSh6KJY3ljNPm
k6sVN9VB+raL4yuupoL2rkMi8eXACTBD+aHFP8ZSwn9GFe+YAQJcRSy+79HpjnBWKBdeAk4oTP6X
v63fImOw3lUw4Jlz8xbmUSKaSQ54tXei0qbOxs+ZSnkNWhKGqQp9pIQrJXIUw0HsjvNuSbQyHgu1
PsRIqRT3SusJTIXfJ1pK8WSmLkTnvvFHs++ypOYtgSfEqzYkWiOJQyKrXVsQCHTv3foui5PueXWX
WG/s0dAUa1OppW46f1386oKWFIuMcU125Y0ACAFenWyeqAk6YFoptlXJ7St+0x9/5ndCHuuCG8e2
d3r5SXF/97PGaQKIsORBGTRn7JxVBD7hCl/nkh3dcsJ+cTdf4gwZN3896jRhoIciTykyLWR6Tk5o
VUnGFZGw8+/KeO6GuIGQkEAnqNSObu92ewFKz9BpwMuWKa3BxsgY1h1zlkWeF0LoDSuNPtUc6bBs
B7m9OacjWmVbtEcDdPtxpGu3wDxaydViHADQFNVCoo3VVYFy7LLLcNAbWVjmTdsz87SrKyOmGHCF
Ov2OwGOYmNwsncqwG26X/ieo6i75MfO95rxOGoST/WtJJeSrR6yzQ2WCQooyWRRzF3af2/cpGu+d
aOGFFQj8gz7L0pykoN/huQOJOJRGLno9eOx8jjOPWZSMIXA20fHkM5Cczs772a6pSS8F0SmPpEyP
rU8LfJZDH8CeONVEvazwld7gQwrMSscWDPqzlvUCrGqS103xMxpsSap9mCvggvJ2ajw8RCCUI7hT
z7i8RoRVIkjn7ansJWisFlrIAzbbmkLfv3F2uZVkzRJ0ZJLvwxpimwJHYx3Kw98maO/XNN1INPZ4
75a7YUFQkrQPeKyE+WLO9nQxdy8drW4XYebGbRaRIpnvYkaHecdwLu0/C7M6BdK+aOnVJlSq0vJx
RdKW0zyMa2eHI5DEBQoru0WvjXWOcwIpbsgxNd816XsTD6JFSa5D/+voDc+q/YQnp63gxGkm+AN1
q98a00GaKvXcqXQmZXrfrHZ6jy7E0UsWVG3TkDzq3YDI2ZfNhXrA3WwTgOj6AM0wmpyBJm+G/FiB
IhktrSkMtUqSOmzw/XClZKJ7vlThydmnDuuw0U8E9Ses5rfYJOXLOEwMSIBv6IJVP2tFIskGOIGy
uh4Zjw21F5NGdfh28QiR879yysNJDDmdKaVBpryJOrY3Gw1ZEZGL1wLUFulxdiuIHuLf4P5jgccC
Bglrgu71VpsBAzA3xJ4LWy5uvsgekaxxttHAZKj365aZLHBXJrGuzr606kY5yNwFRuZUsK9zC1Z1
gx+CDqOdDAaRc5qYpRRYo/RuaQpT8hDEn9wD2IoOtRq5B+wIo0uiF30dptJ9yKyJ4m5i/dAyGmcc
exzIOdbJGEetgWKccfpFhxefOtDWMw+p8K9qMDIReZ8LlDe+qCaI8W+1P11BLGnzuRSeAwD6svxK
rRsXuss1SdN/50o4a61OhJMIJP9fhEXz2+H9gLduGXUkpskSIIh2Fo8NtuSj8p4Dq364Q332t0kM
/yT7+Z+hhrq4MV5pai/QuKCWQAPM6KcjCLUZFl9j6pjW52mZI6oTlNnkT7SKa+GN7Actn9B88/u2
yuBNYV6Svdm1otIFi4SPwCgMMrkCNchNUj+hALmORXLKI80/39+AiHlxWqoQbTx9GGoUYSeKo2gb
jCi2GLzQaA6/y5nesWg4Q8rkRzsLvR6JT8dWQZK002a81LL01cznno2KNJXYMu+Snx/6zSEW4H1h
J1tKY7SO8wM3zA71bOjeZLfWJr2phqmz5mymzF4rwxZSQBeCRtIQSZ835+4XFRumMoG7SLoPSMaI
gQQbyohOuhYf/0xE/y5ODR4+wz4i9E9XSdoxBrKT90SYM+8XfQxPaBjMvHVvflrKP2i8muOQAUFI
3MurbMZTd69xUf2LsMZlpvd+d7EjOQree3vJ/cDy/SnTalCEbAWrfjm75/QmJyij+RJGkuAOO8nU
gVdZLktdJJcfjEJi8+x/5bwszpPTkNPJ/oM8J+EwipeTVc95S3NJR8PgEl6sMif9WF+EuXXT41nu
VgiAHBoBNsN0D24Y5Hq2HfbRejpTPhTlI9re8ickYJ/CyOg8F4TyejUBBnE7b/TjW448XoCuBDzK
RjQJwNiI6pWhjLYAC+t4pM19AiLzhbSIn8nc7uB1292yLxrlZkSAfnFiwBbhK11c9bpXFrtVGYON
aMRpkob/Xs2cCmEW7T5p2yxdaPElwq5Mr/YVkfVDooApl6/feUhH27GaHdzERRDXDQ3s9y+IiP0Q
RgTup2sbInGzpGf3XmFOOOW1zIbgAziYdFXeRKxdpKQAJngwry9UE1QaGpU8gUndEIKdd/gf4aG+
pj3CNEdDJVjK+NHFs8VL4NIzBy1TAdpN0ebl1QKFVBoX2EqfxwDBA/kDwa3DHUYsTADTCvTcnLmj
+CRECePhKmGh8/+8H0GmOsATKtuu385rOlX/2dnLB0oEf2e8vz2REkXzEB4iMbQGDLYAmr46YyXm
KGwaGDAGl7xpdazy6zq/Im4FpFshyQLPNdZk2M6+7KRsM7IJimkmOWq0XuzcvTf15NDqXhedHKSB
qcMIiRPcLExoV0Zv1kVrwI141h+M4luzL/tuo8bdGKpiNw/CuXDO++pJp/qMogonFqSf2jWrF9UB
FWcZS6OGenJl8dT4jN2sfAOHKqaZNRPS46i5DxcHDNWlwV/iwCRILufRqs8C/7PLkADA3cKpmZPz
386+XDRZ/v9TkHl6KzCSxlDnjtOZ0FxqtnVmDsPCosSDHQqPFukARNIiJNYizbAz5DqE4WLKK1cA
sCvth8iba45sXSzqcbLXDAYr7jE8lqeAbB0zOOkHrVX9WWzA+idX0c4bRk5eeyO1zj2BmDXHmmXt
b7mBLsjoHSzGTbI7/9CkgVBjiwy8+hU1MboqSxZikP+UBFzmsJUiUgPTzbMUauu8DZvSR5xm1yWi
Sn79E5Y38ctG7Sxiy+e78TKc7okrUmZJlPHEAkq5R+pT7hTOKmXV+C7DgGDU/MoBxFGY2MhF3byl
jjTAlgnPTa8LFEJftw6szqQkA0wzhYSDW+OPJbtGn0anpYbPXta+T3Ut9sSPBZCA1E2iVS0oOj10
uVQOqC/ysQ72C2N1Suk+tAmLMTc42FXiruX+HLmHs8Ml76vrTGm6LHuPRCUBY3hlIweBmY5J858U
uh/Cyk2JvAq/fZBo9zc5XBYHeWfnffN92D9BJ58e97qZqpIWLgyi4u27engmupLXigvZSAgUcyAG
lMbhQrRSDKnmf2YfcTTx3vA+Vfkg9JBL6sGuiKSyR2xgaeW/mYPdCvvPKg/iS+1f6RjsBJB7zoTs
eVFCM5EL4C1hThvwKcwqcszTzwUDbtBd53uRPQeJ2L5Rw0kdfZOYPJlRDVf3APOctcttfn3J8cqy
vFg/2lbaDaNKpBUno4WMeL4gm9kXdHJSWHz1WaXgCOg/O6wbBvMuJDkE//gIiJklqOJhlE9Ir9jJ
DzPZU8Z2Mt9I45H684yV/ggr/P4o7QJQ774t6IHK4v8hTVsrcvd6TfCq0fjtmJ4em9+faqEF4aeu
0Fb/AIDDgeBs2e4GOjxce7t0VGE1F7mZ8XgHzOcuKV+UrfEQ6qZ8oFD2O7q/xU+hx+VZ5A2WL1SI
/XeWiMtP/1sPco2SGIJCndFQbOY/XA0BEX20njX1gprX6Y9pQpxUGmslTbngeXUfRQVybnFnRcZ8
wckmFFDBpm9mKBP2Cm9ugJEZauRz1niYEjGxhVug3YKw68pTqURs2KlpbIvSB+zoB7wWnLfFfOtV
RggkomHBqGGBrH2sI7wO4UehSUT209aYk3lbi7APV8Rf5htQsoL5rZHcpkyT4u9ipsKE9+Vj2Jdw
YX2wd+fhN8j/Jb+EDTXNFNqyjiTuJEXWABuuKrg9iQozyMn4A4ckUyufnuTk4SD5KQvi6+ERpeFa
1bSdvOEoxs+mmx3VgwYROf52NK2TByRC4Ail7c4OkE8jIfVM7ASL4+5lytn9DTdayM+2td0Q0NZZ
D6f9KNM72YFYSvEwBBq87+CO8idMm11nIfscPDnAx98lxCyKv1QVPxSzoZR5oxBMy816aSpf6Dqh
6VusBzCu81KH+aar/n6p1HYKw8DXFZfYec3urjyAy3DbvYnY3TRDbTU7JGbxUYOty/e6NUYWvCeN
vcdEO0f+1Cr0Ja7rz1vU2s+OyMWdDA9x0R5fMjSd66KFRwHKAWj6onrZmXkmaMlF9bOD8xXLDdVq
eB3XmGTJXpl610vTiFKjz3IS4zlmvlWkAedQ2HNWwqNV2fwq2o4ENuFmR+9BABjm5xSQ9r5Xe52M
1b8HASJi1juQfJSBiHEkdihd6zqc3UZBsKkxjYSbaNZ2dwgl6KzjmpbX3VKjPd3JW6B+U+fcECEX
J/HgtYDSfBHBCdWeF8UYHybGAEtJG31ByfhGR8LwBg8hz7eeotwUYY9LkXAR9y3xFvtZHsOitzUo
ibamrXl08TWVyqj6ROI6GmGV5I3K31+noOUwhyhwREaN8xd+DjzB63OzF9fnXiF4fbgZeghyqOIh
XMe/yzWGr7At80cfyW1E3mQVH4MtQVsrKReN9yZJVTlqu5fPyeqf2socEfJhhH/2fE9fV75H5bTI
1FLQwOAleWb6lyuxkSxCuZaNU5RO5x/VlIywBP4pNGlS2ZJhOWu1b1A4yAiWPu+eclAB4iEf7tf+
xrsdNQ6EgsOf2VD9QGoaBxR36dLJpKpJ4XEQT9/2HxDaNIfQTscZeE+CwYz2cwI+RNOQhK3fFkIV
jbmr3B6VeOSFvB/G+a3yD4NEtxmj8dcY1brOVo6tEKsyItmkoGK+aTaxdrH7oxbshsUjJQmDZN1d
XIGErQYqitcZ/jbBZVfDGcE+RVhjit36NzMRXijxi+hTaH1Em8kP0TEcqmYePyezIXbXj4KIasyx
WibAM6v2LCJbCOk8DXaZ4OpVIktsHjTEupkv3GdTTCO3ydgDvRGTT42gezZQD8+u3Ciyj9UhqBZS
pprAi7lP1MwTXqaRnqRd7NqoowJpzZ10e6wrLqaDpZZhW/5E1E2NRYpK14ynMDGYHO98Oq48bTo/
EkuIDJQJFsDPtrUZ2CJRTdj9b7ZNVgJES9xkxd00aAVQ+MGqDSdjTVu8xagSBmiw6oCS9B0x9vFt
vbqm5BVjVty/PhJc92YIavfdiFNhNoleO0ZTYzg0wURIDiiAtovia0CMpNcugaaX01YcObx+Lr+K
q0inYdhxoca/LL9Khan8UjM/TQt8ylQ0tp2xduW32RbtR7Z/mqZArVeU4AuDs+QY2KkS5CkiyMTu
pKJEdjze54LNNB4RepITOtLDxsqiWgyTYX2Bg1MwSTV/kMzQL0GeACD0/NqiDQqle6n6e41Ga1NJ
y1IqDm1QUcSSV3sA8jfe8KW3OTa/66LfGCg7WKiyqzDWUd1lJV6Suo6CswpJZP8Q1UIii5tJMjbu
wu9GNg6yUpDp5f9cUgQyAOmYoufarn8/UKUiFA1cNF0pwq44lLSPJI0G64hxV+VyA8/VJfm8zfI3
Khdql0lC0a+7WAvLp1Oyv9REPK3l3GZKP1peePmga0W5Kxyr+67gBHJ9eJUnIdSDCDhxtnYqCinJ
J0ZsNGOaZvIjnJVkwPZSuT5KA8UO8Sks/Q8cmz4RNtLLY8YAxExZxnj1kdWrU/sW2nVVvIGKwj5C
Q9PLHHFrxhtCxExoDTAzEwWxXKa+DdG248NPeEntsirWO8qcEvWBIQn2p3gr57JfgDdwFCDYbVi3
Gum1dWGaQdHrwC5CV/PfuKgxwsN9zxwzzdyYewjpDbK7EDd+f9FkDg17qFqRmD3d1wt+U0t1pdLA
nvjOTu848E/hfsO7VwaWvIUnWMcIAS8pTWNAeZuoj3yT4tWLqT62fbEDJ+7aheXEDuVBnmZfKQ/Z
gDG8CA8zVMP5/L/rQisiLW5wC6DuLeyKRcA6/Oxe6VyDaGQIQP3nOLw+afzUCF6SfQ564SrEsQ5q
RMn1P/WrKtB0g1pt1hVd142OLyVt5P37a5izqfTucA+/pHtJ+vzStuwfboMQd2Aw2B31c0WoYHzR
OR+qIG0qaa3uol4/yiCxIH4eTeaL8feQD6PZi13JYVHOUGMgnUugiwamGpBpsrgE2nL2TXPvAi//
uOYvXGTipwoTH2U/oI9PQs4YiI0PxAryX6AY4BTWPYWkstr/cPc/05KoGpl2intzQR+WwYjpvhrd
hHZgWzwQiPopPxJyTC4Wn12zI+U4UFooyGWYqFvSlGa8Ny6DXOQJyVMd3DXXSoLNjvgEep2YnueY
04ERhK15TG3ZM3x11eaZmTJtUbmAWa8jP6F+hisP+zMPGAsC50vZ7naHJoHL6HBLZ49GRsR4lKLw
IBJz+e2AxJvbkRTxE+RwV8U/obk5U7ZiGQxT6T3bW08ce/G68CbLPmt7YXl/OCvYdoVbZj+Pe68a
2SMIAUU97vbnFmr1HqNRC37hlgns1VALx2UAO4P7PCkASV9OdF6DOn8GPvfNuKSbXeNcjSVTZ+l1
BDbK4JGAffecBzDzy8wG5E0KbJ/auh4nYKRA7qdrJBTGMZ9Zk/2I1zJlb4fVZlCNBTrxFkOND8Ye
F4h/onmTQJ51Y/W1Qur/fS2UjjAWLgK9Xkwd12E9r1rTjQ3jK9Z6CGmCkRtTyTfUbX4+GBvnwBwm
2FuMzUUvnqFvHvvL+6TDf9LTkXS9WnjbETsrPUk88rSxpqtXJwI4nW7PRJguvTGnli6tDSnl7L7Z
kX58fJEuix1Fc1bzVy/H0VFxsvlAaXK6gj5NiSeN4Q/NXGnkaotQdIrdJ0rxjfEBFuBHU7el07XD
JZ4ros63Gbs9q7140QsqzzbWTKCuuzR+mgeJWSw/wO+892apFuhehYhKdK913DdnkNFTzRpwpbaN
Ng73mxWmW606l8L2sFJJbalBA/LLDcPRPQx9MLmMg7Flytp+VKiQMjDS8n5Ol1rKsYmrz74ykeWC
w55vUrpJZnA5D/vwzkDmNosIfuDdpKOASeZG77nThzHzoY3LoWJf5CBtwB/Y8ZV/vlwL85HwQCgM
njpfEEPaqOhMpXsNCByFV7tnqlQTi/dKJDlonxnxZHi83xWhixt+xoQOMA/VPGbEj/e2ja7i289D
FogegD6/JXVbBCxTP4GW/S8H2nV4KKOxxmAeOtK7T5DCrD716rd4vjPOZnZZJc3y8QsLqLriO6Nq
ShmSUaKWkO1+6MfWgyHsyF/ACUylm4vtpp/zNMCW1Y4VUTW45fUsXzVKysFHzl9n/YnQM8YeUiMI
++kyYOlSWp8l/TfYCfB7x7ppAYSkBH5T466mpXWPfK3bIA46/k2V2ASO+58CtXvQOCCpO4983Zso
+WMkXFLbWtsDhNpp4QpqANno5THf1dNkYJ8l2EFbCOOXdpm6Ps7IY2ZE5PxcRi2S9pK+imVGO3fv
Yg48kJjGAVvGmJfPksHx9bFOj23y+De2DTy3KTaVdAOZ/lY9/o4JeXLHhH8LFz12lB65Pw/2UWKT
T500YJdKd8Gtk2QS/+hzkktDPP9BVQpNy7U9kVOEyudsX9/1n1qtr01JwrSC8DJohy2BQw+7a+0R
gcizwqSkqbfBOlFW4tjOEfTbtH97mfaCHwDrDjmWmEYH6Of9juUBPItik/e9hmbl+vwp1lI1H4q6
VgZBr76YWVr5y+QQDpt6wIlD3EtnF8FOANAxSkG0FUN2nhe/POV3814O0AyrzC3nNqWXKEguH6jy
XF1Zc0HcsWvFohN1MXDdkEBisBaBHpOxAGHFlGRqUjONOGm2E/pwQJ5OmzSmUr7mzmnlUHpP3dvy
YsGAAVkpTADwh9kZv4CMjjWAkg/E/HeuNqVPPMYmIbMLe2aLHcrcaf2AHxhIQ/z8vwgDaL9Em25r
HKsEcGmKwBajUbdfA30uvb2XPbRVxwxlyQL/Lm8aB+I/xQk7XE5IVaD/gET6xj7m/CdCt87xKybv
Opmog2fNXfNXJ4Snhos6/6RkA/AeEeeKy3mO7PzA/lV1qqmx/ay6NloVq5CAPltPm9f5wjPO5bXe
B4FM3+ZOje37evMkOmk0x3DC8j3A/E6+GhB5m6zRoapN9DJ5oXqlleySd+2Km1e8FL10JWIYn7ck
/nC2yXtXop+01+j4tRC401MC0Rcx5L8ixz5foi0utRX7V6QKeLkdMPWLPL347s+vtTlrKi+doeMP
WJgPYaEh9pkNW8unCD1QXR1OxoKgvl586kcECQCZIYN7BhbnZqY7WS/vG/yp/RM6tnh1O4At46rI
rJhin4pGInNeiQBIqLrxuOJly+cGhXn54hT3V6oBIsW53r75o0rIZ8Sxs0RlboWXufx1uwHery2c
x0lN0TO8N2H3D3hbGZo5DxQYl+45wpHM67ENxCpvnABD0AUTj0Dlc3pVA5fkEXhuZIG74vcz3JTa
Ff3ewm+vTX6I1cMAEIud4qeVZuMvUsyBCpR68k9RNVtH7eplBV0gI99LTLo111Ick876lPgrpTrn
r2G4DEX1KNe/I9HR61l1AIsDXFg9BQs5sVigTbm1s+lbOOA0xhSZnZcNJ1PZjdAxJpC9oNVBhI7L
UuEAU46BBBWpvNWmeSUSuy4ZO2mlX3Tf2saYWOzf3Ds64ige5BsoKq9jYerQNc/h5wLIJObqPeP7
bzFeHDOjsOoC2iRBsUjmzan4BCcrkSoZFo+LFi9nfjbwwUS7/SUw1j8lnVW+HlMmOV85FNTRfL1G
J/qMSIty9Z3lNOPPf6JecW6neGbXHVAdX7KivXSqCM0Qk2GuKiYzgl2qOR+yZm7X94smeliFyejC
kVsVFDXX9JEC68L9Ws0ppvgJOUVTV1x9gbbZBqBKkdwjhPKFEdlmPiYPICPv+HysHamx8+nfWr13
o56E5cnnocpK7ree+x0sZPanocdDy244qfxXS4lcbUdnGqAg5dbU+uri6E2oV/o0XOO1+EGlMkTc
3U3JooZXtKovgvj8ZcKlkADpmD0uCvoW69by0RIUxoepo7xlAC8TGRUGqNitk61WX7ij7Oz24xo/
cXzpBO+O3Ft8muJBYypkWVWxfdyEvqwn8maQndjRkaycz0yHQr2CweT3KtgXoKlfCjKUQxwHvHWd
iodjPpgW53OeV2MiV4Xt72jm3wEyITqLMHeAbfxDTfboWXDRZr9KexIy96/rCjXtGvbdgRH2aXLU
jRtSA+UPYZFshDGThDXN5Vw443oDsJ6ARVdshh4KskWc48fet/jw/MVQEdOIB5xkZFAnIGYErYyx
NRC8sNEih9S9ydFd3tqw2P1/M88a5w9VZ+uWfDIzn2BQGaHITJi7xIt5BBySG74l26+2lnkUrBW5
nFf6ts0q1DMZX7SVeQkFaAXPWn4nk1qaTX5QvEb8K6NkFzfvB0S1LA2n1lPnBGIDoIX86/jldK/J
JbykVILxssmp2R5QKh7Md1KrQhToxPQS18xkabbXAOQM5ywfRnYM1ITtb/4GM7xsfHuUAU6JSnt/
a4Nxc236CwquMUxZ4e/Eyi72KJylcu+g4l4apJqDq6rX0d53XLcaZd5erHXVyaMy7RfZi0wtnlHA
EKdSXKga6aEYdrd047yEXv5622TOinqpnv0VWa2ebkk+c1qTdxhLJHD2ePsZdskMDq9Vdo9LAiTL
XdR+9vOX0bBzEn8TCpUGlWW9mrz/UrDDMVxUNZkpZr5OMEcKMvhN/Xe6uDEj6K8ZgijW2oqYbCSj
Zv5NURtiZkZGeqFjWuEh8plpspUHKQ3gJxQ/7sjRV29yeJLNOUnkqKLm5ZR2/Wh3tiZ2pdOzANer
LYkS7vm8v4Ey07ytdV37J0GSptfigEPfbqyiAsbFsrGhYN2pTnyLpM4SX/wQOimu9Zve3I4vUbGH
seUm8KOsc3BjiudF03RV8z7k0UOsKe/k6ayJc31Z4B0PAt6RJgZnSgSsjCkduejk6zvFX2OaG+gb
kzaReLK5tN1RIB/0uRgqypugDpLQt0mzRsXAo+G6HSzIFDL0zijzNB72iFv/r7YDfrZkyV+DIQHg
EaVeWLKh03B9vdQRby2Kt0vbWHR7L7Gp365dBfOAw4D2L6DW7UjV1ry0JVlvL14t6CDGla5Pzwtx
g/HbX/mcksjEdaFZYFCYNnP9i/wbK9iS7Lr0UmrF59vGIRwLoCfzqkwmvXEih4e+yVF5yKrzuPyQ
s8JqMzUtdW1wql8TcHh62A+fafl6oLNxqCTmKrtPtNjuP+p4P7n10jyCYNtSRHsp9V4G70MKe7Ek
6qJKPs9m9Zm5KotDYvKRa8ql9XwuEnMkwmlNxYG6Hp+s8Lhiq9RHXkVH0tJK73OYtyJhgxCYO9Oj
GjO3kJT56xSMeex/HMObt/Vcwehxly8B403J/QbjvKh2nAO/ixLnxPsXN4H+BkzWv0iS08Qyb3GZ
8WxASir+jY7aEinz3t+0LiAr/tYCbtnR++y10YzZiga+WEHSFJuvWGL6PB+lDR/tip11HBHZgraW
X6pbKwHHjpR3duGx1ru2JVOSjo3D0r26z8WUOUWqwqwvinnGc101cS4OnDBeeilX4hNbe4QsABq8
fCJHaafivFlwoDHeLZsdsXHMFg7Xgp8OntPXK6zj5hmgvSLGfKBW2eXeVxM9nsz0KtynJ9nQ/SD0
xv9T34sAdCN9RQCoD4EUpHUalDKrh3fH67RHVffI079rij3YoMMIYElUjgGlzBu7N7jeXdYLMh/K
JI4FdBV6FmLIe0E92piZ/2TuNugtRrSQtUh0rgJetMevbuARXEe+YKxzHVH7J72g86bHzMJ3gE9m
dsIO5I8F7yTRxNFhRzrc5EpBo/crd/XpKELK4Y+3OaTA+O0AE3T2W4YI6hNi+pOKnNL6pwLdGUsL
Fs6QK7qbz5SK9P8tOPr9sv2oiQ4RrTfy6tOZO/YrBhrFDkek8aBf0z8hVNH7VGB8ft7T0DIysCI/
Ac/UXdoW4fFBoXE3BOeiGeeVMzt++yCCsfm4e2nLOWQM/d7+SfezWxXaoNHUbLaem3x36T4rOzDQ
cwHgoCHCJLFAVV8KipoqFPeeS+iFaclr5smYQ4eh5vJUPfEi0rdwkpmwjohX4eEql7ElrNsu0UeP
F2H9k3j0denEB0PuA6l6GF7UfRHxRryGYgAreafOp2CsM0F0Y/PC370GqT/8zNjiceGBvoBaZGmo
wTG2fxjaELFo2OlRggyoX4B58KnqkV9wWCTqzJOQFV/klZR9zZlipQJ6s+M2psquSpXsSosODi1f
yD0bNK0PJDITeOD9ijou3TZQtm8uuSU05p3rfMWHBp5rxUviwwOcywNRLnihuKGYEiRu8YfrQvWo
Qd3iG7wejDXI0UXhJ7MyjaxVWEyLfXYd8BMqq1zksF29r/wrgg2JVNZpE8nVNX3kSn1U+FktDY0n
HYG8QXpRW/t5ZCKLtsy/H5dcLON8ch5fj4Z91STHVBmg6VNhUs90a0ifCvm10t2NZawrOe+acU9e
i9KoW0m5KPQ1ucqgS/lydgEBT9+8kiR1CFSQ+i+/x0KgjprB5CPROrofMD4HcRCRYtlLk21lP/1G
88CwFiwOlsgjcdOt6bFGElgk8ujlr5HOgX5eaPGfFnvF9rmpgi8tysaAHLeiOztZ0hLEhy8p/T7n
lCKq6ZvXDqbnklm91GUxyVbVCKwkK2r/3aLXnPCT0lNGv8wFz5JpLvgO6iTi1wyBE54LkjPbjf+c
34T3+gPDVDcFXuA5tjCrp+a084eP7LDm3GjHrKPlMebaYd6WlBsaO0DlgHkR5S/wy2MrIQnVBjCK
pYyFusXyudZnfPl3vWG+EJRwIlabaZWK6F9x4Ke3vGq81CB5hn0I6qzKD3ryFRoDnKgZy9BzJASs
/G2gM2dpVTbAaE6EaMRWZygXLKBrTl4GZi4l1V8zSSUjc1BTC+7P3bRicB1wyC342FIfPgVFg2yu
5b+wkL6X8SQQik9BzYZPvYz3a6b7E7QQ9dwuD6TL+ZtfAfT2Fmmvsp/8AKJWPA0dPoqj3QGVf7er
jfLIkaiwzgneFiXNvfRIUJ7FOOQ9LBkqwgnz74kmmEtSxvcNi5+ro49Mn0m0hKX2CgIw4S2jPihK
jG/nOv9VYKyJTGzNhjZx1Oetx3alhOXmpaAr0dSBcbaCZ27wOAlihgkrV7PqKoXafGoMQWJF1Ox3
ov+gDbv7oncFxZ3oE5kJKwgD02E2FEtvF84NawwoKCiVhHgNGQdk9X/tDYBtD3+n/o0a56XlQBm6
9BKdkGwlb/eXOtgYCrg2r73o+X5cCsvKGfPa5jEdN0h9kbI8Ni8dj+iFPkUMQ10m4J1lfmPcpG45
H+UmoqWlYyWbIuKLRkbyI2RLmQ25u9Rmmn275RtvLQl85VgD+SPKGUYkeNWFmuH30TDUb4pVFKXY
nBr+eiagJPEHtKxvsJYvKQGmWKQ0P43H7wrm6JFyt0yFLt/owngAVQe79Q8XYY/x0QylsEDe+nVP
nW/RGQXTk1K2I5AXOstjokTkjBAqnvJuinCHhlsI0G3CVshhaa+ZLSarrBQI2EkFsUNrQbWansWu
BxC5DSB/2fzJR9ZlBgy4AQIbPzOG4uPKuWSZyjh8vaOjtGBNbLpOW9YADqhdYWgXnPbs0WGS8UHx
U6kpWNJ22tNZJXIQmGN0vUJHLK84kQEkbNXvN2GvO1ozqY7zRMjkfR8YGQ3uoxNZvsUJlidU6g2R
tBiICccH+h6G/jjNev76AeOvmnu8YSvklWc51dXbuz0XrDkl4jl2ZQ6k5711XJhbfUUVO5UBRPbb
Tfhl+HtA/k8I8JnfoeryICGJbo8Lnv79plqJbV3VSYUAPctD6/JVcYMwYSCFy59jPH4P4TCAlj8F
Jss/7B/RuT9PeEPmhFEfBK6zmVJhnIxhrKBNqWbZEa/KpRUhltoDhx8kr8Z1bdnPohaOUWL0F+FK
5grbSe3ASAEwXM/p3dHO/86YfwcnVy+7buSA3mDQMH8Jn2mmfMJRWtRHSSahKQhxOY16uf9f7Ep5
9bBKmDjWrGj3QRuklv87dsi+i9CpDZzNBihmq6OqmgfqUNksu7nLwA7sF7GCA3EuWWyhPFcN9ill
Rb5RVdrqw9N/59e1hB2No6TePpu+6dywgLlQ+ZvllZy8596/7DItV3SXvPT85E62PxKg62tR+Jz+
NTIGlbEiq9cZOIZ0TdEYl5TwIn5c8HAhw5nDFYnDlB/Jx37wYAGwSzkvO8cQCX72F1w/RiRPGdJ8
urazKzssWgu6AFHR0DRG9xTC1bz1D3sMpcadcZcMcOw15JZGJfcm01by9epLF37pZke2D//yw+Ha
IcfAAC4qogI4o/HJP7d2Yn3NvtW5DZkW/T+0FSOatBV4dcetMZ9adWo4V3sTSkbSmCUYTtcxRYtm
IjTkg+2YiqxBvVLABixdLv8EQWQAF5jNUGUYWYMEkrIZWBgQRoqdv0DFULY0v0p+hfEKWbdP3L4G
X939UVvnLQP6Wn/yjY243JI/B5tJHHXmWRZcLW7j4AxBS4M9/YYzpX0ijlJNmhp7bx4oa1v9R0VW
btGFCvKEO1OVCzZXqmL4PFD0tFDaHaeO6gyP1wXBXl1ZfN+lKDnHP5mM6TU10gJS/WTllQizlmtM
AU/bzW1E4YbTDhIKIHaJNLTSM0VO1+CXozAbnetx+Tq/Oi2/WfQHog0to+LK9sWBmB6i9Lo+olH9
phFxrTdYkM/X4wVWTVRo1mxuG6X5HW7vzfUPBHsH7/9c2LDNAwa33hZujPgliuqIRRCEoIvA3waV
nWyIF0iq9dnYoH4olrsZDsZsRCSdx9typo3AUHBVjybYHvqvUQoaNchD6cp7tlxIiuaMtxVqIpvr
PfOeKBi8LuFkALeWuJsp8azgovGSCmyOIWK00mHsN4dnK74Aso5VNo2bmHBySna2toseiPJdmB8r
ApuvKc+/9gdgIKETa/KqSGs6INeJSRR8QCAMk17Ra2AasQdfdtqBikB7Iuf3Co0YwQuJIljzbart
jslt1kttitl+gurkt4sDy4WnwJ5dBQZfjiExIkbXKnITvu/e1s+JUTuvKA9we+4NZJGQ7lMN23mQ
yfxXLycW+COQ9Is20XTCOJu44NwazwkBZ0E6iCCyGaKA+bG3tJtU7ga6072HLKE7Ffq4CRWEDWrr
IKGkxVCNhcPT/pu1lCvDt+tb6tdsnMQs9Z8tTd8MsmNA5R/2QSBMcEDUVg1CJpFaNMJp+fPF4krh
oXWIyOJl3E1vmbolC5S2kYGCkW/x3tvVNm0rw9A9AcmmxMVBDMaiq/D8qGd+kNHvjTX7YxZrziyu
yjrfTFSvpV2Zpe65KV7+sAlRMcTH/7VdCc4Bo6jyDEjRieeaBhVEr4AjcCw8EpbZUzrJdZCLQC5D
B3byt0MfY3PVxA3f49aDCFPKTWBmbDokZAq1XgulC2GvJiu2N4ecfTUrYtrbQELjvFipt4giwobr
JFewyd6GiFqzppUs6i8XUc3AAnTMve1lg/P+nGIyorLatmg/jlWVe26H/mWQxkREC0ZOc2bdUjYk
p/wVOGY4r8Xu1pC85HqEoIQD2ySUdrQ7eBqayLdYwWaWf3ZwZNqATYZzV2sOBYUIxPai1b3LxcRo
l38e8Rw0Uga+pGrprEHophpx8GxuSkbadNfk5cRsgPEGiHXIL0MuY6w/tc12b1oIRWVYLfl8mspv
It9DBiwGg+dMI0r19+IqNMwHe88JE4HTE/ny8DQoDnBBdksIld85OyHSl+jJPEPyI+5lfhkB1Ttt
yfWUNu7G1350p+WOujMaiHO9CZTjhY/moOEfzP2ljg0XE9PwBOFE4vipeFvOuOnBmN8Oq25wod9d
9yvYcCYyfl9ZplSY2S/B7qBtgwevAvdP3HksUb3+LfwQpkEg/sjhPqDqRE563vKAnUUs8xD7fWCp
z4bKb4BylWOKa17H/+RN60hIriUvt0tC2GvKXrOKETVOsyDHSXBYe6o9KoV0I6ZbSm9/RDXEHcTZ
tlU1Mj1SsGGoHej92OoNPldDSTdImP+H8pAMb6o5nTT58+mbRVubTQ9T9ZBefMcu1ULDiuBoS0f3
khvFEpMAWYpSY8oWo02cfTUB/orR6Vd5bEi7UdKMQCR+DqLRiVAHxyMpe30/7ERn6pePRcU1ecB7
Gw5WUkAXdfGe3JphxIp9rU/M250WaHOIPlsY+PAQrK08FCR4iLxUflBoXKHLwed8rBYos96pM8IJ
dTzExJGPkxUcVDszmgcuqmRm2bjJ0tF0EWgo3Yg8bKNqbCnW9Q8GAzRwczOkweTVffAVu9tcOyr2
CiENxdJNSPdg1q1uxSZqnp9YSBsgVXhNwCBFiXrnst4ISuHXJTwy3Gx9zJzK5P2d6akgIDbmE2rc
YbnTklblT8TMbUpostGSAB7MaSuD4YG48OdESp2GWJVga3HQDMAaQq87m8egk+sEmkLRMEIUruVd
NUeMigxbNF5oaNlYpqksbwBJRha5xSUvWRZffxqE97QWBWPejf9jokFf32WgU0B0J+NG/xzkIPgy
mnY86RMfnZdLa1vR2ShvwqiT/Ut7NRxQHj9K3P+AlAiV8anH7VfPePFKLuhT+bA9mrBi9XQOISao
7fZItcW+uCLtdoAsInznr6ey8/coY3fijDknJYrlNpmr7GoQSpxZk4xfYa8Zuj3vmvDqGVTlTnJl
iXPKcuIQ0IFV18t3FCB5BW7g8K2HlLM6R8JWQLke2Cev3C2GSf9NceJPDiBmXwmLVSjLEy6PjjfZ
IdIrKxs0c/012aWSUfIVwAOWXRSJnoMft91p0BguwbUVYAgBHbHBvhXLRwQtnoxHYM3KBiOnzvTN
KRPb6yZJzn1RL8m21rS82hys1JqhZFYTyxRXfboPF8Z+u1rpF0ybY35egU6RygWSZRDIcxjbnZHP
vHxKR9yoY0wqG6p9vSwolpOkH7BDhHFTCKkXdSwxt5jq7EB/6YwlhvIFXqMis6RA6zViBetxf4e4
ezaVapW+jF0l/tbh8um6yFnVh8WNh//4/gg6sJwwJ6seKkqy2A9r/CaqilkCm/2125gQUifKFw4n
puXK1F6mc4z4OUcZOFeiCqjIA70rC+AbTsSbnYRjZ9MwM8cCNNIh0zvLnAYiyypUzf9jqPckgVQt
y+BW+VFVkhKERfOzJLj833qogLQpL2xjzl10T+YPcQ6NAAhUtutVmDoYWezRUMswvSfnt6efIBfY
yKBRrPhjoj0vS19+bPbbdboXBDF7G9og0ba5gMcrCpYQIW4p1I+VdSDlyaAjS+/hN6CNp9LTJfNi
mNfiVw5Yg2O1eGJ0kz6RgHPWM6BMx+BIrPOeRGaOG8VHJ4C2+aLH+nb/4v4Em1jI0Wf5lxvs4O7O
FsS4o1zsrzwi5+sPqc5JTNMrXqef6lXQQiALGL9UF/ymvJJiCskyBfM+Z0u+ngoVMo1KIrDZmuQz
rLprE6FZxaq+BElQH47gRUCN/OpBNF7Purd2eXDppFBB2IJeJBFE45q3Ia+54z1FPD/SGzLDLdQj
qthjEoAp4BZDY59gGFAuPXzljDVszwuVcip7FmkaACf82C4DahkF2wyfXE2q6oagjdfryBIXNehl
x8AiEmVeIrqjnWgMg1WWeCWEg7UgUhbLml3kDUEu8cMBMTbdooMMwOq0X32/H5F4njb0/vMWwnaB
fOgXyAPcyvFw4MkZ/CoTJp9GahymUFljoVKag1/eAkOtPeBbk6eEdsGjWx3Cs901Ye56Tv0DRIKS
woJHQk7F+AVwPkmrqsu/61Rm4c6AJll8s4TYWWqAVMiYF8sQyt8vcxUVoReUcOglx3SVTnNEm7b8
O+CgqJO9CecVTSv4ieKaNWdetMab3JN47uIlbGwc+7FmJtmJLHpLPgw7IpzinN4XSrgbyPup6Xvh
TxzCNODF8q4qvC4oKm5C1XLRXZpGAZTrWxi2Ns66eYzafM+S+F6Bu6jicxdGBRVI059dEXi69RsZ
pb8UJe+sKKNCgCndAsWGMYQLV/HIB43xG/Gg8RQxLWU4gelvadfwKwp89+p/XrLSrOH2fMicYR71
OEK64IOLRji6YfAaWFh1DqVaD7G/fqImRvdZgzacoqvnF9A0PTWHmiPjQuuT/HKOyDsryvjFXovC
jaNa4sTn3xnS5FyJR1ZHi3YOeKS+SEweqgAZz7BLQoyn0++6DOyn5PsgdPCKyKBDoQ+lSQ1V1Pna
1E2px8AgnT+/3Z69gt9UswCMjwLdI/oG7+cuRagMiK8uAYCWhzQ4cW5Evd+VjenaOv5Xtuj0v9dT
tp36KNQAT9TelfWFD0yjzNeBjSAYkSj3layRTdn4oj2hQX+tCcc3is5L62bT8veZ8cXoduIEcEOi
XjD9ZMScWvso99li/4SHD9ZwurMbvf2Us66dXerpcXCcPRf8023ITFqNF4sJ3Nu9t0XKEFV04LD+
utmcKDILIJQYGqeHF3qqc8F4bURTkmvkvkAmE6Zrnwsr5xFAaBr/o7ew+G5kGFOTr/nrh1EtJXo7
3sAmrTL9F8hwlgnXXzE6Beh+/ST8N/7QCj1ZdXtIolsuF+HaFBI9VeztPjByz5juNUSHHXgB+xov
gekegkv4k1HQJYWD+9CSYe/QzMBf2rGmQ2clVs33YC36ZjGvgA7LSCg2Ku+ZeG+WrSTTHsDIRXVp
Vx+qt61ZM0KQ9srNGI8llfNY0jUtQllV9bNBq7nPJy+ZDAEW2v9BumlB10GZvG+X2E/V5Yu/h5ng
j6GrziSVEnFgrVVcA1zcDqaBHRWj2ZZxesr1fCODx5k96kSDxFPKGnMWisopSbqHwnBJu2X/FL/P
9CRWtLlLsm7iL3gx4gPTV1rUxZtD7gt4QWArQE3GxOQEDu8dORpu/yEU/jMS0s7057B4KFiOzzMG
kjwBW2N6y5h3cLG+FH3RYMI32JAAXZmQNJBYA3JnlXaDbwTDxvDneiHF836NU70iNJpojDgioC9m
bU7rbZwOOz3knbaKUpCKDhxpdlAOURipcXvTxWKX6Ic3mVqQF1xtJSvOiExXZqKJeInaKtKBJpVR
8zrVH+9PUNc+CBE8+Kg6zHSv6Jf2kcbkwlXtVaiMdwQClZ2dMMgBmD52HvPLTKLF0Ac8yNJ9JHBz
IAb8APSsmIy2GQ5aaFsz60eHo7UcvVRmSf5mI5xQnIb11kNRkrswsX1YmcNN6q42ObrDOmAoU+/r
BHXsBFj1yh5ZxJ2tL69rXlUXwhOr6S1HLeXbcKbrZbqwHvpCpjMtAjvV8AHVEF6qeR9n5n+qG/x4
BX58dKmytf9rvZZ3m3uQjd7m7tFE+H67ykKt7fCOyO8q+jYDitkwWx8uYB4rJ79DHuPcMZeTvC7V
SlIL/ptJDhUEdt0JaTjWpvMPINOEzXIIcdnJoQ2Vho9c8bFxRmmb1gwIceTibL/2tdhpczAuVTGM
rbQdxezIVErsQkwIbZU67g6bTeTnKoaAdbOrrXx3e2QYnzEb38uGbNQ46ZjLGN7Z1s/Z5UBY6oIN
xKdXN1mPpEEamrPOYLw2i+mVXGFJjA0sG6ZhffjsVUWBM7s9FMrwnWdws0hLHssJvopHVqkOLHrB
mAnvh2nYYbZd2Yw7uVpO6q9T1h08s8M/+ke/ACeFRlvhGE/bmYbjOTHaPa4GdtKt4l+7diP0Y2NO
bdqsIdRfh9xKtFvcFDeCtyiuMpCgfR8GymRHQ8L3CTydq/FJlIA1+2AnIJ4fR5WpkJGjcajnu5uV
B+iGWGzBx2bVsQnfByB2XcNk8bLOC+muKaq3BWz7F/wmFF0LQpfHG69bZ2259je3OFsWgrz9/2e7
YehkGqMyMHgCZpsRkVA5dcJMKgxsf3XQL71Mya7xcEktQbuH+aofp6M/EeUVR1rR8B0jPe35BlgP
UE9bvqLksfIiOzqp8dGsHSB2SAkByQlub1ZBTppCQmMzW5RKqEsDjHo/WgotJBO2GBSqqmNTt6r2
Vw0KTElGh64Spbn0R1uppPtqxmzpWdS9+f5T25jB+psqVaxL2jeLu7jF2kfLA6jwPwHemn9yt1Mv
EbeD1WoZ8w9LJr0H/58NnvPCl0+1iGaqzjI6eN27VZQAMFhWQqcbES84ZlKq3bvRiQqJ12Gl4o1e
3dMMxCQooA8tWrmGoaUNH//SjJ3uU7LGLvf9LsIzr0M6wqKAnb0KSGNiFCltY5qQ/uuCIelnvuZW
OlAo5AhEWiT57zpJ/6oYkm1csPYnfBornnzT/2FezLxqHrFbMSZGbZ3rLNWJVksWJvSt9kGiCiPM
kNa7xp6AX3AWyuxnXQ9mJNsrVj1ix0uQfcvUPiPAFtoVJKnsXNUP0Q7mIhpPjZDI2im1ZxRTPc8I
9ysmz23fK9VgxEN8la8b90xZAFJK+vSteyg4y7s/3Xjs22v78bljFP3ir/U42ARu1If9wGG6s9QL
Y+PT8pHnKem5rOA6T3du51BRUQwIZ5A6EoI00aiDp4yTFtWkx/daGOZW197rmA9cw7AFkUBPbq14
ek4E3t1OW0VrSXhCtAh3uamsMubWx57UnI4Zh9GZjqZuHl7fxOJbiVpGxKW4sp5usZT48xTn5xiM
QJWp+Zap3FMjKf9U3dAQ0HFKstoTFyXUDcnkqXzi1ZMI5bkrClRsAKjdDTPhyddzh3fJvypVhGvJ
KU4PVDcbCEJoibIaU43ZbTobL9CQUMvNm7K3YPfa8Qgkt/97vFUhcg2eSQhHKgLLko2Yv8J1wh0u
jDfn7W1HEBHyZCUDYJck0wbsEB1oinMNavxXvQ/2sF54TjYGNBbSHmh+LX9eZftvG3RyQ4gHOcni
PZM0k+uBrclhPOQ+IKIDguMxBX+qMxy2rbTTTx1MR8zfM2hQj0aJMiHelB+mSlkcHd4rtAroLKlt
XIM2qi5FPWXVvfS/pleGYsHzAM7T+wd1ih/tb9jJLLqB6/LMcvhFDkQkemp/b92xCE0AYtDWC3Nv
BTc0aIBTqK0HytV5TQ6JPC3WOdEkpx/8Xi7S01gmS7Lmsz7RSBvjDYq6NnGO73JgG6NgaHEIg2nx
kOu3hoFPUCR17ftYkKUCCmcZx8qgWzKMmgO9u4rBSL5BrlYb5nDy5bphqkn0eruK7bjqQ48lcJYy
/PNNc2dq1UE+RO3yNcQ6LSMDAnauyl7LJjbMsrC9VZOReel6epWnL6fw9CRBs8G0lSKSYgiDWdSn
Mz9fT0au5/IP6Z1cHDBeysw68Eaeh6Ir0z3Wf+GLzn2hhYc6kE20TlVlYmiBf1Pe50zuEfLtwixb
uBkwBsNXiqxB0y8MEP/YZq8hb6edu47wjjblsxeA77nyJZsH9i+oRJ1TXBBo7j6ZV4ULbBYpK5Mb
qx4nekSGfmRbrdwdxz8CbEPz/oq7JG37LLwNDgpy7/NfoeC1k15ZL+uNSsx6Is2rV0sJvXrIgkeG
OEwVbvcmQLZZseu3hNoxy5tOQD5LKcjMMc1ZSlqOXHkMipfzx4KSZAmLgrtioOFuYSCTkY33uEiB
hTfihApqo1K9mZSgR9QULp+K4e7SAbaaAQ6kL2uhEEfzr+hBgx4HZVsMqq2/6Kvj8SkTHBc6H9Ne
LVH1jnXsb+dU8p64K+RUjEh2jLhsJUOAnkffl8Y7miyiMhzXiWcu8dCxi6t6Po6vRawvCsin4wmx
dfcUS4Cpu9iATTHq/VYPTbFiJZes0EPLI1IJZdxxq6YSGl68LXm8yYiVPfg7ZHX2EIkldud4yHmm
DUgJtVZ32jrqq/VgfuLXAXN4NbH2RyRizTrWh6+vhn0tv1U7RRH+drH9+a7Cc1nYe6PyCQu6eMCZ
XPcgf6n4pYrW5ucdZ1K3pNJQiYyI3/nYQccmUjKrMxGP4XLuzZfHBK9okG+FdZk2wN8r3G2Ik17/
ez+ViZcAZu650L5kS7tzkCeYFnYECYjJkfGcQFvNstlJPfcOxYezrV7Ts3TMN1rpfntDDK+nCLgD
CCly/JmfZ39rbQRaoDtHQqJFz8bjJC3S33pteJ9DyPRIMjhbFF2r2h+4KV6ZD5zni78WM3znMzl3
4jGZMJgO439S5LIFc3k7CBs+r/cEpvDEg5uxJq5g9Kl1VhtJp2Nt7w+pxRW3k8XFV0EOAbp9YFMH
oyFbg+Y9B0EgvCsqJtoL0eXS0x0KLsUEvhHvuoI7gxYBF+m6/sGbNQC46q8gTzP9HwJoAmGTMuYZ
P/hJrZ4kO/dts7ovAacWmF6OET1kblNtzUKEwP9EUIF5BawawxVeBcpPB1E6Xp90A0zFRo4qWWgm
0JAHYAfMGUp0h77pL3o+ZAksOYsNpKpdQKfWhgcXMd/UupoNyGldl/JmmtFVZ7afUgi14D/wvDdr
kcYhfVE1A4mdlH4hVSjS1so7dpQl1c2AXUSn2lhd7IYlAOcNRhFjeaC63rFoiN2LYtR/QrugD0Mm
ToHEjVoi2wTh/QKVTsmpEwFFhNgekqV6X3Vz7AiMRAW655QfOMAVRBKLA3D6s9SDaHb0XunF+AFK
E45PB0zY8WZajB5GGDvbt6CIA/q04xp1w6Jv3HAKmXUioNGHDWNnGcMhs8bPHKAGaPrBCzMfT8n4
AEFnXQVK6wTOlOSCwCwbVaggvErM8vKO8XQace7pgHpSwgC67wH/QQHgHF00yhiPQuS9kB+Rm+hh
AaLNgWOznuJiAEblGHlRiJ+hW34lCb9q/3exF7AjYhUhoILdohyHqSu84QCBPrhyU64XqIyAmgLP
y7/AbDAOri5lSZCYcB5Qkl6KbhNvemKNUmHY/6rgSWutRiZVbwEuRv1/gdfsTH+8BISxHgyB6wPa
CXlH1dtB59T790fe3kXaJe7UBmvxriCwfFikI/yzJBoPI5WuS/3RebmEMYt51f7UbvQgekzZcBYZ
bZtxU+3dwiDJ7B3qWMa6af9pn7WLlOhcCNvevHleh0OL8eFKOc+9yMps9ehfzaDRwVtIrYjIoGm8
V5wiIeQdOVrIxdHEJ32D721u1/L6QPwYcO0z/oIoK7xaaH0FWIN/kEL6QzicrciIXl4hXuwXIAOq
g65Qz3T+Mqez19bjlTi/qJi4RFkb1iuaJiDnE9YbBvPtyZAzNhzr6i9lQKhX7bywaYWQ2hFb6AY4
L1mJtqGz573vxkFvWdM3sMSbuXU2JNEfUo5NB62Ub4CX2CrXiRdxHmfVLSgld1QkQJe2hBMZa+lX
wtuDLpAj1DfwN7XxNfftcCwl+JuO6lTF9Y1DP2Bvl9qCybGMQg4BHUfBqa/65mt3tHbFNkQU58ft
eFkd/PCc8GmGcB1IBTenj9dgusyr2JRelifvpLwtUNcPfoIJbYdzRMGT82ABa0Fb+grBQ3UfZyMA
ZHf8K6RNia+A3ODdpI6SHO21XrBY5J6BFe5YK2eh/d0V8ykOmqFm22QwU/GfpNJ2wLs7+QwKnimU
KAwOlxQKEHdDeqpjx75V51m/s4nULmBxkmOJkN5AhsizzO2CKRD+NdOzUaE/sU9phP6hlO/SRoHo
XAK9Va0x5/Txrhw6zmP9U4R0gW4bio1/1ZIuHsYppsxCBrkyYaRvY1AALkBbm7SCuK+2CXbef9rB
ZNJnJnV5fFQV8K2bdkGKONvF/5makjWs8uOcXx9h9Jrv5CUa6ZS/X1pvgPQS7RsAo1rm5ysPk6t1
vca3xzCTAOLofHRAkfl6b6NxX96DBxOAZm7D4LDbpMjKN8pcM+xR2XITYgy2ZhA49gPNOqFH1QKF
QzappnaTLu6R5Oqf3t9uxTIs8kzYQIwqhjnYW3S6YhZ7jOHCb4dD9v3E+EMA9C+e8/zc1YqiMYPA
egcw4S/7cKpHPKz5ChRvPOq7SsjQEdWKQrj5XqQ7tmuSGQXd7aRMBJ/RUD15lLIwI9RNp7cQ+wnV
kbvMESfT71EImy3Di0z7j/PVNO44qSbcJI5U3rbEWhG8BoN7chZQeuQYbu/XbMalBD2QrrjL4IF1
8vdKH5VDnDR7vhkpNZGQAN/r4VQUA7ibX/MH7Gpc3rJE9YsqbkKAijPN8JKYOKOwyZDQ680kq3/R
HBWXRCdxpex+FQxZvbwZg5v817injIaVGY6BO5YoNKXTInEJbJMo+f2FbROQDpBotvmJ606bHUMH
MHew4/sug/sCHvRQKSLSes3uiFSoJQmtQel/yKBKAyAZ+yHyATWABdaZJWdAGECTooNj33GDnr5W
UFP1dE5dgJ2zZpkc+RcIEpEuscN7K+WFNjfpq1r8zA43M3NQtEEXDl8OhyAYseUCgGQsKMDllsIu
Pa4R3KO9g4QvtnRHwBbdsNjXGAHF7HhkGFJrmqV+LHmrVtwSq3CaGwH7J5wcZTgibR5iPm+qmNox
wyDp6nFm4CKyABvdxjqLNcvwtI+WZYjJCV+ZUuHnHqYlT7M+leAfhAW7QRQWIIrwCNaEka7RG4YP
689ef4cLlQi5qSGe5eJSRfeuP7+tJU+oJ6FQy2CpbkHosmI42c+STfQ7IlpyiNKb0dDuL+1Eploy
OqpZsZIesJuDx2AbA4e5UMqIpCUKVAdBK8V/wFnEil2PlS/d/VJH4FCqnkQ0PFp2buCUbKr29wSz
C8T9y/WyNjljyOhAh7CL/LBeGqnS9mdStsqRtHhlyH5zmtAoTvlYcZ7XG6NwfL2UD58fkF/QVnXU
G1ZEY5T1epXqZNGYrE6QJJ9PdWY5mupymeg2Q84u4qyU81Rxr1LUnPY7E5s5yNLEoFEpFL7Bx2kG
2y3Cp4VMJrj7LIq0fSmnPAzv/Yd/opRfq+HIS0FAvTyhdUPT9jKtmRd2npZB7B/UrE8E/Pfyd7Jl
4qazyz3owbifSliNK4VYJnXA9+S24nMynCNLdohxfxZGNrNjRGCFFv1Xc62eQrnCwQ6s6x64DC6N
Cfa0aINV5/huBHIPyOY2KSkZXmEx24YU7cy7uSuu4hSyWwJwt9p6/V0ncDfhOpOmI/RaRNnAqVHy
Fph4sg9yInmw4Q9/ysR5mgBOWaQw5zS989XV5QJDZTPpf2KS86fZuzRjwxtWaRQhoduQghBqZnMF
k4cuuHrgljpud19NByydjksy8yQ8kOdn9GaVxgfyby2pMESq4e5QkhxUGCHrgoK2q1V58dkxinvY
Dn53+jeN9Dmt3MMc/OsB69QW2NhGcJm9H77neRPo2aB8OmjohSITmOgweqVlUUx4kd6IbGUrGcIY
cCdctCidcqxQ1yt1f4J8zMjals59hZfYpt7ZM99rCqpV/N8/AC6w99jQ8nqpNcaZ2jzrPERIEptJ
Z2OjNufpD0qbgP5WXqt7WAIE075Nt9AgosHrOe/VjsgtnuQN428scV883zdDM8YkvoJRebDvyOZp
xl005tYY/I1Qs/aOeHsIx8NGCpi4zlPen3GkPsM+qXgQwB41qbHxjTBgp1j7pZJKPqX00ZjKrgYP
WiJYh6AsMEdF8N3L6i4fx9eA5Z1GA4qG+03wRHiIGF58RQ46rz3BeP7SWhUL6/HYEdTf8k9RL0fx
hkdtKTb2aVHPsc8aighhs/EZ+lg3NJzoaNVY0Df9TwhkijyQXghwV8nJAVlKO7fAWulm3DcrI4rB
4Z1g+xQ91v7N7gNAol8UOuMJoFUgTH4XemrZtHLyDHuETGIraV990IpSA+732vArOxjVjXGQWfjY
l5dC4GgyLblUmhYAEsd/EJgfxkBBVcnJZgNIrWH04ZlXGVCJpgOezRBOuEeDV+au2wm/ohXzc0JL
QcnPuR8tIFyDoAAgx3FHgsEoWaekXK9lL/RZi5htps0nqCBZEVKNLAY+kaX6yyT4/F6n1T2Nwl85
W0TloWClRQamqomTCNIr4qmIzE4DC6cLKfsBgHRCT+5wW46VgA35tKhM7N8It262vAuJI37cDu9c
NMAO3fGJaSnfSzpSzYik9awqCXADEKg/IYcBtbcRWAeEtncoYYxOfQWDdJBcNTtvF3m1BDZCw6ev
DfBBNlINkJ75xoNiCNiFlkEFo9gCduauI7L00BohmwS8N1VAhVFeS7tzux6IDMv/uDpXxIjmXBpH
IBaJHyRRPovFeQOrS1IEnrxOB1KeSMr6bfaH836nO2llUDgBrhVyfChbL8zcuMGCU3fEJsSLkmNl
ICtlaKL8DcDUhri6/fkdbTKZn2jliXX1ls38EN+Jll4nXNouD6qzT++tf6m0Lg4xMgZ+XHYbGQ6N
TbVR9NFAmxc0gVs5BQ1Uvf5tKgUcVw7+XIrLR4Fbp08KIi3oPOqDAeSazG98Eh+v20UTYMqHoCbf
k9TMoNFxJR07fGcXmDngb6ZEPZzBnd3xpaAs5u84hWZtqmqW4L3/XjEI6y9nXReMxH5ggGw581Tx
+g0LYYeKstVpU/6UYUVH3nrzEFSeDbm29Dw9Fz5hufj1aJH7kxLPUXU/SuqqGAFu3H9rEv30f+NE
8LjjpdCwfnRXIfLFJq2yaC/nK+docdo9xo6sn5WrObDmONdvZswTt1yARDJbtzzDk4lRzITvv5QN
5qSAoHre8KcTIwyJJjq+LCQNQtp/A1g2UZIzXxLReGTvhBG6rByYKIBl2GZZj/Zfk3Xd/u52aAR+
AJltZkeFmR7+q37y1PALI8EJF4z5F80J9GUy7xvXBnafop4UUGbL9sx85gNlZmM91+4PJlDf8SS3
ICm9qMg7qD71+pd23GMZZDrI4h1jNaAFq53qf7P79MmMvewECgVL4SzXeZiI1qvQg2F2Myhm250+
LIicsNpAdXrwEZv7VJwk8gew10RT8EW+wpIqvob8ky5pRz6dhri2Ns0kj2lyHGChOCeXsSwGl18/
RH9K2iz8qGmX2RXT+s7oM3z23QFwdDW6Jh/P8zZx+u+Hg4NwsBqGUSICltBpZXi1EtuMDzOgggV8
pRDPqn2Al7GGriXh8WXZkWHJOa1nqKcZoD7p7xxUBW9buS6POof/OM4WLmo/0YG08lABsvnTHnT2
rlDv5+L5kY9M920WdtaWmVFKnGaTi7r4XQRtKrRtvliGuZdWLbhyc0T6fS3i/QEogg8V0h5SZNTe
DVslunS6Oc9igrieVGHuZBFvHOJRcflj0VFigkDFu4fz8wDCEJ7ENNSjecNX93xAdQflMWc2Uizc
7kHCGy1Q6LJDAk6YoSeyPfC2koRv1tXpxJqeC94bL7po9ADErSXAXU7ss4TqTsbyVwsxZFk5Qeec
sAUmfOr5AiaNtaorwFs9D7ir95Gl1aEMCz0XvDkkxHBGb6Jm2Utk4S25pZWxigDzFESyF9YF6VG7
pi20NXXeumUgaa8D3TnzaRpaKu9B/ntkG8UJgz9ETijn6oDKVU80wbeadqYVjKnI4ZPExeKV32cu
6sURwESh6vPpRlKtsjE4GcE0I8Ar44MOnRCEij0ILSjOSPxtI/9R66HUBhPhI+jspFqbbf4ZRH2E
QR7n11u4YkkBm0EfA7W1Zw7rjf4GFx6qJYxNqht+fh2nK8aVWYsZOAHF18alb84b3dOJXRtfzWEm
UwHSwZhlUm9XEZn9DVMXhVfQJG0V1G76G453q9GpDd36NtjrvLrCv8nYniIsdw4/ELRV4MtW8E+U
K77f4wcfGkmCxpqX0pUFSHLlk0pUhjfQJiWpAfkWI4NIO9DTfkdRGfG5jgR+ZwskOcsnlIyP7KHy
iALjmC3dlOlfSfepdqMAW4QMqQ5Tq8O9nU/6To/cd16wzJdnKrmhfsVkghvdl42amA9LRC3rfuQ4
cO7pxbTno/PZjcyqNYJ0ZONI011jgNxWsYyxNt47mdez5IgOkmuRbzA33WMELevX9Y5z1R97Jtup
mYYAAxYEKtJkh3p5LGQmH4x3wbsZG75kpWDIyHVJ7NmOFW7wSfxGStwfcKrSHKL0iusvWp9IwiO4
NjS0ZoYOqaXp1wEaVajH6SxYTI4+yjhei6oXazHQKfIakSaHrSV4oLbmgMvIz8JgkBgN3i3j1dyL
Tkzg7WsTU/UYGlxwM64fy3cXtJkb0gyrPlF89gUVxgeaE/L8ShoTNTmP3+mgbc/sIEhErgNaMVot
lDGSWTYgqB9oBpuOtPIiftUtPHS15jV9VF+XiaUR8ZnajQVB0H+tBzctYCMzkCWZD6vucbTrS84+
tSxO56ObkS/5LtW3ABIll0+8mS07nm1b/me1EAgJtCNhZMNfQZgyp4PomHiZ4JExdzisAunnXj6x
euGzkE1i2JkP8g/3zfXYQbMfXq4ebwjSKlyLZiQPGM+R9ITznuFHfgwz8nUYLP/hFSGMTFNPFvZH
4djBKj2OOz4mbT7YPB1dQVyuES6rHjnSAiQ0JSziQbpMJt+9wFB2chV5k6UEqAd5Vax6yNad+Cbg
GGPeU8A/mclBRhVDbgnxZfpuX2FyI4eZxLKy7PJxdAPfRRAHn1KH6JUuExfD925i2NZ7abeiL86I
WSTn+iY+91xmAJILkipMlvJwGGKPCV03EqOICCy3HTS6ZWvPnfcew3NSCNsWt2EuSyZBGme8RTE8
C8t7fsEDH5AtCnYhCAl/bg2ooMzx6asX0qw13UX831z5el2bd74S4WSNQfVxRmAAWITLY3luMASL
nYKxkYpuoFyil/8LTB6HpPwWbW2EKpDHxR9NbPwrkprPCDUhpApGARHjJ56spXGhog4bclavwKHt
9pHt2Ji9y/9iLPyuBzKwnlrbHe1keEosuJEhNtGKGe2Pg8aLWRWBiUoF07RrU9HsPnfu2sqIWSi6
PUByr9L7ZcdmG9s5Wb0hqYmRtRrRHuZ8Ih1lqhAaeiDApJcYKqeuudPCBd8OBaT8KsTAIlYeXa0C
EJhWTyuP+U93Cwh6EKRuJIESQYAr5aFUFkWoGcgK8m8oVoJ9fgsBNN66pyX8AQPuka29BohqfRC/
p1b0UXPhKmkXLcZk0WTmeCsmxZdMcm/nhumuSHOqFXZUrK7dNvNakWy3mExFSoWmtpw6qtO41tZ6
7c1kVufGeMss4ii7pyZ45/BGeVellevVIlHOSt5+XGhS+dy0NUU1f/Dmro+ICfgnbUVvVJWkWI42
5jgLgegalbPNH94T0SWXiqRdVK6SI1737sGLPoQtFzIchJp4NvGKgRPt2BRi4JYSI8+cH448z0iN
/jUcVxX/sU/RjnXJYzQYIefZ5AsqCeQDadMFo7SvNHpucuPc65IiBc1sajZw9Tdhudgos8b5oVvM
h4qZsQ7ita7K63Z+rfJMby3eiBsZN8+Lf3uEjAQrxbdm3JRcX/eBAJkV/MWJAHiNpOB7/tkMkhum
u6oHEkyuFPFkqqAAhw4RJW65iUlaAAiNzSLX7sM0UwhQbKhMo/zTHcYMzMh9mEYAf90ru3AACX/6
N45UL7T+cK5bnM/sGnZztU/ZUMJUqudHTGi3RharyWb0WEBLLbNbTmlA61FiVhNL6EGPn3FHLqaG
ePciug5krSqsRqiEWdG+wngYczr9RlVaxkh3MZIJ7G6vVTNmfaUmCOVlJhnzYtLmB1Ks1sWe6ORn
szAbQl6fkfOJWntPN6j3Vo6akkx27WRTrXq61qRCaA0oazJ7QJ6AGDPq1VX0wivKdw/Fehl1bFyW
ZHUdNYEzzZ1kvDDtP1mnb1esFj89M0ONW2q2gR2Cf9iUGttL5lGBWhzayMbsddlfVNXC2jK03r99
ER9CC/bfMHYZuC07cFSZIjVET6hCxm6CmxufYmwENSJnK6kpLElipWeLtIOrRzEiyVab32jU5Fp/
iYb+XmPsiMpv96+tItO2aSu85WBlzDXkmLcaC+63ly9bGDqTNWnPw7F2xT00MzmZJl8hshfCj1kl
iF3mN4YW3OQ6a5+QyWIG6RxWvQ/Yc25WuHBKrPgPcnBhogBMlzq2GTjykRcKu1BS2AmVwe2882KP
6CXORn8RkrPGQyus35Gh/7mkRQdyw/RiAyxUmj/uuH36Fqg6xXERckMrkSnPVou0F24799JSgUIG
UvLf8IR083L1NGignWbthGtAzTUz3Vj4fYzWir9rjtKd1FHZRaZliVI+c1esYwmiio5AkooeIBm6
aGfKluqxp8HC08GXYrOqXB8roWYs8h2HItVr+QSY8QcuUloqEAY0j8CU0r6vRC5/U8MpvHTqMBvp
qyWdsoYwazpXvrUx4bwdfzm91kU73pWfBeOkTG4ruxci1UiRb7yJ0ImfqVgLvUbp7q81twcjeMIy
s7ZP2/Uhj1JUrym4XrCCVbNix1MbQn094YPncJTYbsgIrnkR+pxc4kexpuSVSoi/Tdv7zFjtSk44
CDffmdi2u6r9hbEG4t9dZ3FWne08ptYqNUceqEJyz6jKuNDYsOZyvUrubBzGQv7hb/lKW/tklZ19
mu1DWjIfRLAmuUfN62kcqE7ZqouoLODqdEXmKwq4xfh1apvR107cTnRGEsoK0/EWF7DoJH21Vr9h
+Rvk2lOo8QBXWaeRgzIpiQ7IYvnpsPzZbFgh3IOBVWUem0juro+WOduq20odNe1//Q7Lv1U2sQUB
MAWFvKAqRIpT3avs/hD5OhouWXN1GP7wetGpvx9HEWWIOgmKafkXRbkUZh/Crg7BrnF50hQzf9cr
wm6sNNpvMX9UU49rl+ZFnulIPfm1N9hn9nbCtcrWDBSb4T5abxs0ioIG3jTUE9aXaHUvllZLV7HO
yI7pCuJ5gqzUMfL3s4NnVUw2CNcwtdHnk7qZnOGuwNKLWRr5cWjbE0PN6KPb5apcINcinCa2i9hT
dWmR2fz0au3iX0S4x69ORGwL+XP6WJUqAbjR+4TwC9kx2H9wlAdFSXfS6jooENqwRo9XTireY0ED
VKz2IChOwzsTvMP4+ZcqhyQcfwsp06x+xoD8UCTCc6lLg9OExF8xG050Frb2nTF4hYe056OIIxq2
+KfWYJ8HKKV1KezeWeCCBYH5VatpWl65bGsjjt6sVoCfNbjMbHByEY/hGTT50hH37BOc5OfRheUb
0L+ANK09cSZ80bW+N0rFZBDUWBVUUsRcsOP8vHXD8cZTfpZW1fw0DC+SWx0OILmSPGLjSgqPs2Zx
d1XKuRuhVdIcdEcsK218GflcCK+1HFhY9Gbhf38v96b9VoR4FwVEd/StItJ+FAmRxxV/Ei4SAfwv
MtC8kLcT0sSLIvVhSl0rgZDVApmadVoo05umBQvhrF1D0caBc/aqpwLl7n3to1kYzmJq7OaXpmfa
VicfTrh4k0G5BWg1aIjvXydoukuWVTfmytqUKh1zDWyeLF2mJFCcwHuNkB80GU2rlvnPYkvrFMG0
KKumyqqa7l1fRp2H/BmIOEd4YgFSwDNcQLXdAGGCF6kBbqZhsw0PawVuINVxHUuJLTlYhL+7elq1
Dnt+LTt62nNHaeOP/n2wViBTD8/z1v5LjkuxmiHrum2keIuAOfOTXtX2bUQv1wMDyC4Odly6QBB4
kntXAxUAk5g3qreJjvsT8MH8WUnddf9sd2xz4ASfybppavlZNZW5D7JXhzFWPRgxgfIxuepEibz9
ks4QdWOSWqBdS1hCsLedYBfbZQT1jwLdsfTsvRZLfV87/uYsOTz9d1KkDCxJJkj5xGd7yO0qBeRH
PzN91jqQa6xHPtXCXmaRvZ8vH4lPk8uyhCCrtrRlra/CCjohX8wP1+n83nmjYeNJSEe+oYy3rYoY
qJeaRE+gH2x+3nNLLchKrI4OFohDSFj31fq9QD8CsnL29jZtZGCu68h7WoFGtzjXDYoKuHMgANtf
Xwnb1BJ2An+j5msLCyo57mzGoN1i8/tjlL+MeX0nLD+czdXfjcOUVBoQ8uHKLahnlxbs12Pdzk0T
hdJi/FifWepPOPR9Tvpa5ReW9U/ePCwps7Jtp3CJHDtDlGl0nLCo+brJwWQhd51lwHEOGRZQrVKG
D6YbFR8oX9Pzd9+RfpNCEyLHI1ecTDJaJYIu0BcM2fQUeE8AoV96pvA3wyg4HASyAa81/t5JRVtl
N0Sxt6qQMWFVR1/eeysO6oN652iIwQsJy1GLGvzVTujfG++rE6FZeBrfkAjQCChhJUB0Yaj99Gz3
DKoKgU/QCbpO5wlP81/rG5zTGBUnNBfwmO233AHdQTYigFQd4Es0rWgzEd2YTyW7dQmKHFZ1UXLy
wG3Y5OC+71AdpvPE45AXB9bBgOD5GApAdcOnfSaBRv4XK1wZARBgTrUSlC2DqX55ZH9ZWgZ+Ag3D
EhbVTjdbOaw55pE5byTKCmM4z7JMH9IJkDe0dYubuEWFS0K48TXBva+MlqEoptv+I+PIfqE5vQqN
SAhhvwex/8RBlPlvdvjWzPeXJe59W1pCLP1TL4EhOIBmjXR1j7yrLU244U9KtXfJBOFENlyRUMLP
Ra7fq6kGfNJwqQHgDOZCMV3/JEz2Bx9mAs5Gax0xGe7qh2jJ0YrKFNuFsjJB7flvmC/l0iJBgP5z
fMo8TJy0owOaSmDjjYjRnqxfNLRpFeBBB6VUI4NdLUVNteDA2DGwJeeihe008Kr+IHbAqMVlL3Xx
HYcnaZHMalGki/hJrEh7JWWFO53/I2SqcdOWt+vsrlYWYOwJd8I2g3Y2QYwotVovt1xuhVn7GvVS
4H8q40802yTgJtX6imqzCQzSU6wgrTRum4VOhWworIG64sHF/nmbR1a8HbqX1xYK9dhJvcHczwDg
vOb40KwadfXOWMD4+jVarssxX21ZYtu++4yIW2MB2c+dtRZTj1yG88Ou0u5tDzMBC9j7igkiGAyG
GUx395s8M7m16rxkUi27UOCvI+eTfnf73//4ZKs16ra3SDtBsuqkmjEsefT+s8YSw7BPvFXOFjpy
qtw2R94AQH9TNORHnpBFoLMddYisO8TozzhyJZ9bsFhiThwNn2BwssifEe4btgSU1ufBaGZnYFdn
iSDSWEFwZFSBObqxCNyToL+xNoS+jhjXxm50JOB/ebmFDtadh+LFGM8tbI69msTcx8XSGnK3ClVn
Dv/6DbKFhb9zUXr+bGs02Z8NgA7+ksVECioEYWDnlGkwsprM5uDGzpL83e7oKvbu9fk+aF6R6BGT
sw1OPrftYoXTmzO398s+Euc5wykkXiKdSY0mjdjNaPyComCGxo5rFJ00p2lJzuWZufabcS6KHclt
HmM4ngL9tQUrz+gup66iDcZ+DDtNMeehCagGSQhe/0NEE23+C1EM+T/4ujPoH2+QYqjxOkDBVgCZ
QqN6ZVPELDIT6IqfbaaMDKUpyJw7g3saKNkii+UCw117sfvqFZOnZA7KzEPNQveSZ1FeG8qO/FA1
gWkahDM7sz0jqJ1M4cyiHS3F7hcV+wqLFGs/DznWV4kfU1sm6rjaet5OwPWwa7yM3qWql+Ln6qtP
uILm5SksVTYYamWddMBj6sKZs7rbV0ITKoEQ671+2Uj8NtmvW+sz4sxJkVJ8opjelyGPdnWKpt1Y
ntbT9IHRbEvEUGVYDweEr3E0FCE/b/Nv3JQwGHrNpF8Fws+3tkfYjoW6XeHYhoeK4cWNPinMx58N
2Ea4JxLiTxg7NRi/K/JpHQND3cVWuOwMCWNcqdLADsaeZ+yrVwx9XXuwzHjZdpQ0iR5AKlymc1l0
DV0hiIXRnpLgsm+lCWpCqx56Yg0GR5br1Cj0Z8oHvxuBBBb26YF1e9Rv/Z1LAxRajsjF08kF1E90
vBqLcK1mZYJQdtjUvkG2AP+hyhvPLCtzdlEPSQxSjdZZQdUoHPJ0sm1SC0Imgk6dohUKsGLdioTr
175l2eY6M4usNq2e6tBgUd/N9f2Unn6LZs+cEVHDo+dAqUMmKaWvAOsJLpnZ432ed+za/DYqHbsT
g8BLQG4PpzsAKQczsD76s2AK2JXBYTmrmzpizIb05FSp8LGp0ot+lNCwrYp2mx57444LNctCsm3U
xtCWtqEiYSRD8aiLsWxoJ3v843igHThFQ0nxOO2TYcTSzDzl6MyvDP3SOq9pbo9gDTpmrE5Dm1BN
KU6MsYURe0AnyQDvufpgUFTjj4N/m5wrMrwVXdOyOZaEpKM90TT+F4LUO2ZKsMwg6rMLAgSIzbER
Vh5x37PMqcI2f3hnh5uTw+amWBb9JZO9mnXwfxchfAAXWRWu/dBHxDb6yBBPC8s4VmCOuRG0O/9F
oZSlNqosYe1WZEB3UK30sIQmJbtbh5fqVIJU4N9LC/f6igcDlhI7JXy95cqsr6ycnI9/o/F6hArg
HDVAPQo2zkt9Ih+N8n/QyFn2hoNOKHjWe99Omu437qeVBUA/ZW3qaYN+o5uofQFwhXomEBto9/E5
rLHr1VCpyWyrz2IMPoKK4m7nIiNTxW4twGqc0jDcj6FXhgZBpgdMzoNjhgCP3rmOOMW8Ep+ZhmEW
UcoPEOWvqc/vPKEhNsE5TlR9iV8YcJq/HClBEIAWp3SPslgMOqmRIMIw7BruHxc0PeylFqrBOa9T
s6vtA4Lk+iPI+ryrf868meanbIDqQF9EcUGly0+1hqq14AhPyZW6FlhU/l6m2rbssZnYhykcGNGK
JJf22fkS+MmQ51gbhsMAGfq4dIvts5wHi5zfCJ/LYTNazoc+w3v/SJabMpOyWXbIbqfX5UHKLrpo
XMOpqNgc32cfQKev6YPEyVMhiADVPHnm5pDTEA3HTs9qBtFVnhapN+UtTU8Ky1AFDzKuJF2Cc4QQ
8C9l3gjvacs27T2+ypVFylIZwW/AWiV6Jt+uACh4CG/yy1b9tcBRpq3DF2xhvrM5S4EBh90/HExf
4x0W+/ANhwxqSK/axHgYkMezXEBFtrfdJjYxoXKUHZQPSVRragTmdaWBz55IBC3fbt3vdWXku9Gw
bqsK60qotWsma9P3/OruQ25zmSDyCJ2hevthdhlaK3l/dAqtp6pFB8LVc4jmrsEQuQT0Cj5nx8PQ
00+qDeMi2/4Huppj8k23uc64eSJAqrPZckGvEvwh2n/Rhj5lmOiL0/dC9hDFtw7Nowqm56w9B7Ax
lIRBb9cUg09btn9HLKRXK1ZlZ61hO3G1rKg0ZhNNSxb769tlUpkkQn29Fk78c4ld+PDiHsrcbzI9
At6RnjnXHbtznaC7q3aqqa5w4eJ7bo8mvIgl19QG7TVlcB2Yfj5f/ulN4ipgTFcRI10KVGCHWAYS
gfUINRt/+aEZNzqpD4VYxcd3OlNysM4F7ri3hGb+hm8FwXzuKIA3wnku4ZtWamtntdm2WyBn1Hi4
cN2OVd0w7K0252UBwW4xHSHeXFxqmFP12iJqFPwOXw0ng2fRES8gcE56GOXrgDYmq9JLvaMEXD3Q
ti8OXKmMbTYz+tbO9c/He5LP38DyKyx74KkvDwWgFNpMLScb95WEbeqLjZSBQAL6DARh/Pcusl7W
3NkZd6AkmQ0k7zqUFosqgFUaDIGMsJyatzABuXR5lPnqygKhK40stYPyLuheSN/6jQ9cl+7roMW1
sBpGp68jk/w/lDbzQeH3T6Yv2GtqT8h6CysYgB53b7y1j7iWn4pPbbowUKgwVWs/xT2Tl5jJ+QS9
0NYtpEMrE9xL9yPbIGQMf1h1FolMzJ4bySLkeS1sna8QxWaaDrpjbzifRSL/IoEEAtGt2kcfrsIR
GilKfbcu5/S0SHODJpbAsBtpuMwiNqizUTHMPBrhiZTmqb/z5u7ocLl9FplkJ0Knux7OLKUEgItj
ksUGypB0y3YiKaVjj/uDA1AXm7UoDltgH31jhENWIKJ7VY4dbfalOPVf/Rgjh5OjVDl6Dszkft8D
xIBZa0w59/TBUuEUPzkKu8xykyczrJwkjRziuaz0OMZkUh5UhF1UR+j6/71qHeDPMKXGv7VG0B0B
Q9o5ABK0O2KcdspmOAoCE+St71HygyU8d51ksem3MNpPw9joHWyx4wLFZH570WNnOl6phtVgTtkh
AMaqZjMWNihOYfIWPGIxQiaE5tXZEokZ01jl2zV+/9rWt4jJZo6CIsA7P3tN+p9J09DxaTCS8REf
wQL6pP1Jl/hSayFBj7at//uaaITkTNHilGqNaAF6P1gR/ONo4vVE/36ZDwzT2pqvjHTjjlBxYyVL
O7GAslJ3Ms5kxyBZUQgiN5n0k/30044rNimwYCW1vasfjpqtMrJpb5lf5H5WG35HEjw3EedpW1sA
T7Jg+jgvkPQCzeBsWeXthNxwmjn7r5Symrac1VobZz/pc6JxJxeB6IRDUQDFvr21jxlcevdUktJW
4j3nnKZCvHEEOVyg/Uzj7GqUtVUHfAMVT/UwN9Oui96SELII0UJ8u3+p9zKXfe2m4cP/aPuCzN6c
mAP0Ql0XXArSb16Ky/iaXOZl1YfjPyRUoTZAL4ZZi8maQRxwqY6x2PyvbYAGO93+s/62jSYS06fm
82cohX74cb8mXD2oWf8u7r6BbiKGxH3KaE/iYBPRUVD4xuo97XQypC6guinV2zfwbbwo30NgEXp3
4nnNrPIZZxiUX9dZPlNRbSKUTFl/IEQeLu8Uc+GpMoZa1b2DyrPDEDA84NNB3TbWJB1JCYBFWDxw
vv6Y6MpDFMaYkv/Fnvdlq/wMmN7pQkpG0VufvYeEBjsEBUKkBEXoHyqhqmzWn06Gy5RhkeQGd+Rj
UA9EciMfwH+x+5XEWVq6oF1kU+Cgo75Pm33GuJv/hnA6PhI14LEiUKXeaW+tE2EJbhGFm/zQZgLv
9dK3Xs8qWItOR4FyhhCVchUEcXUJG+mWYuBQniO+wKviX94yxP/KHiK3w7/+x2FuLQZchyliBYmA
fhB21HWPFuMJaoAbpHHsl+NBU0MwA6CmFODPC11NkqRC5pEIDZAx5qcn2feKRvTZPSOZuKR9eKkW
PM59pfvRqii1beg0YZy0BrW+yyaBfyZIwoNL3RDevHqOU0OJPvxqFj7jkD2wCIUrtwIpUxmTze6E
Np2VUehC054diaRC2UpbL1iOaynz7xJY4kZj9siElfCzj/BS1Uj45bPPoDsdw1rczwNGQanNRnOp
PzElGoXb94GtGOsdwbp3by349x4D7WpHhxHA85MPEmWIkd0cQaE9GU9DVLUZpfgfmHdH7EFMCids
NKYf8plWdoT/7gpUg433y+2DZs54XqJtapDrpcTXAtX93gqV1VFkRVjgdhHqA0zTr3ryYtx/AIXC
/kPU4Z4tlIWw5UIjqCfgSK+eyi5rDfYYWmH+vhLiQvdAsYtXVZlv8doXqEF7vJsVx45SPwN6fkMR
Wlzh7YUKMrmlcoT/QKA97tIkQ1daYJKMIlW82OvbEAQIs73nNBVIKF8agiu08NknzEt9WqBnZ2IY
H1NF40dtfe3E+DOH7fTaZMDIkWeA79/HSePtFWlvEVcV6oexFoy6uvIhMT7eFK9c/dEEIVU/nnjx
iLs1Hdk8vkHsffi+Of1GMGffEmRxGFVFHPseQAklrrfK2P2XCnlcxY7g5WPvqPIO6zbILQycJyUK
bjAE/zMpSFp/AW8ifahZZIUfbnYz8ot0cUCJUk3NBQ7XNI5hypOxl9IcxoG6rLSTwH3N0wir5vfc
/0hSLZX5VNnKCDXvl8UthXjdKhx9tZBrHh6nn8JxiaPtELDOl77soj8CKqd/Ev5MOLpSpw+QwNIv
gOQKqcsJfQYAI97YMTiGhOW3zBbXKxuS6UECBFPKAWFUNoN49o07de9/IZdHt8i49jPEas1KJDtV
BwOUoxdbbT3dK2Yaw4Ohlxgr7yt+TXhklWUl9jFQLvP9bGRkxTgqd6aU2vDzhTYS2Ni0uf3NYOib
8GQ6C1LnQooo00y/MmDqPsP+81lVRCLiTH1f7VQgPgo4rihYStXcdFrnLV60z0of+cDSfjvj844r
zCYVaZMNu7SJWTE5b6EDhWjss53reG3tcOxj0xdkk7TCrSIeE9ByGBLDi4dCyPwy0fL5ngR5dm59
YsfTLwX/64lvwDdnHhroZA9k2fujJnyr2jocH+Oj6vKsw0jvMI+/XEQ5nYdyni2L2awBWHkyBRob
6I8b6BancJ7uKfNntkP8nkeVmucqQ4AVuhrQ6JGXrhqkoQqKD6sTQTJHAHSQnSc2gVTyXnfJMaU+
RrjeRrmGgecFRk/A88qLwbXXTdO+h7QxwAuu4Xl3LuL9DoeApNlc/RoujUuvHzweuveS/V586vxr
zuvtvXJ06KEHAkoIlF3j/TLBNI8DItAzx+NmkxacO2xA38/440UmqHANWxvzLoeU7U0JXeB3WIUj
FYnqwW9i2ofUiOXK9hvO90q0VqydyFu5izybKzViPJRynauKAt627S2srt9PHI3bqUUH0QK2LUh6
9ksHaCopDQbNJp3dTMgK4WQK4XS8amNA/anXYzesQTkfbXgVb4Pj3rdOxmbtsVjeI9w1wmu8ZpoA
z4IiZfhwaql4WT2eoT6dDthGFgcdkAcYMVkOokSxU+b431k9sFN4FhnguJeLyzUmRf41fNLOxNAe
ehE3pGQRF/YWbbdpGzkpjHxn/eV4ONClm5A30DPl6PvlSLA/nSXSAxmMi81taOdz7vfdcp8qJmzT
x8dDHlhHsSGdBS19buoeN5Ec7gXq88Qbar98j1dlkTJrCMJ78GXcWC9hvmBMo3aZkT1SmNP/R7i/
O6Ogd7YJsoHxWWuv3GFolylKIuJzJKCapWnuC4AfG6GGq2J0kL83O+RLYjTYH9wjelVYrkVDU4z3
6ulTOSE6bCXuFtKgYRoPb6+eYaE38imqLy8BeonPTWWBqbMkoNTU3NU7C18PmWNV/dyF+Ff+Knlp
tg2xxiMjwqSjw7/VuiYjHBTn/YJwGWTRPLSw+rUtJDBT1B8c7887EWZ/lSyfo3EdcfOJ8j+t/7Wz
e6VZCWyfA88CE/moIuNmZ++znPROA8QyOWILKMMRAj87yLim/nIv11qzU5TQj8c/X1ipeyn8tLNp
YACfb5brk2pJjzEAk2Jx3ZFR8Ugu/klf11P92lMvcH0Mw0/2B39gCDQ1SJzpRGd0YBmYgkcEwUzs
Xe2OPaT3W6lESMGdVgeLccdJLwXjSWnff74nfde/ckjOfsOC16CTElMJyamobl9w8rO8I/R6VHRA
2AsXWmNVnJVW5h34IgYL1TP74XKgGMKVt0G7cq/GYrDKO1Tlu7GE+rclDDbf49Fac6dFwaRHrDiC
Onv/KtTEVsBUx006avbBUjPyuuMHMWEE3YXi9BjiulVriQI9PXZJu6O7Up/a2PSOhFJqAy5MiQNH
oepoRfnip/W3vmJEPPMTtsVyL6NtubVCfYMuYj2n0s8dSYTpc7x7I4A4oWLszwTOXgZbWeV0SWfG
xQQNVAyZgTT9mzRDnPlg+qPlTQAzg/VqkpVy4fw6P3UeSChKP2+fTxmgYg2RfYn2RAEizmXtXxY3
xVjvonfr9v92jO0nf7t6msJfFJ0pOmv2hEfs/vlO5LY6/9pXju6RhlI8QqCZ/K0DeVIJOGo5/oLg
yMx3ewU34eB6wcLuQkfZ1kSwsJ6OIGVB7CMpiInRfuLDI/+4EgSuH5rKGIbx4bgVIpF/TxPgr3oE
0WCJsViUm6oPdrU24htuznSm45KxkknCmz+XfqvL5YYtMpeGpkf4+5VtmI5Pld0CU7cEtjRd2lAr
RbjfVIlD/KOhApARNk9QE/86aNVhix+XSqTbn18biKqVZEKz+vXwF9AcJlHpjmtkggp+cusihmfT
nufRKa90wNaMUCnfpWxaKs7RRyOunXW+fG3BsB5eWL0+bthEaDAOQaaj9LeAAdKMzN0nemf4BdMN
PuH6exE5lYMMHN7eihnMcPo5vz8oIr8YFKGJkXru1z8NGMuhcRb005WtFcE21eaxi3ls90iUP//O
QsFLbfxQnbKPKAus7L1XLtMbvX0l67Iswj8i1jonou7xaNMpEyTWi7kOnlsGn/jpOv7JBJlaz5xW
DzzwTAF7yMbyBhnXTZuEjrEp+nmwFNqn5P3JTbmIIbWqrBkj058CJ3H6F2d8RjHFzpc/u6gMMkRP
FyYUVaBaBfjYwIbyoQ/DkkzpaZPXyzXRfLU2fp4KLGxJmapzHLB5OUoMNT82a+fbVRtBXvomZ9ta
R+j++H26M0yU43LQrnBtXf4m/KGNFO7rUZN4VJ7ggiyO9xTU43T1kWBrLcujkPj6Mvv/OFcAkapW
teKdJqQNZHrhN85e+CyVE2nzAdvDN5Znks3//L4OAxA8AZNL6YH5QZS2kXl93M5PoO4jtntZ6PUw
pIULl+nK+N5Jp99gLwr4PzPNyrM2gSzpDs3aeJLhDZ8n8doIymeD9aHuEOXzJvLTbx6Hq9ZTEsS1
kg7T6UY2hnwqgLjW0+hktSgu3cy1tegs5O/qG6EIbZ59W7UMq7Clc0UUzpiTkNnRKCJHF2ylqkia
jOnQ0b1PElUNqSpOrcEG6yPj9URZMggfXqRlSjFHaIM+HIW+h9D2F0MIFsKbKMZkOGuHJsWWQJjx
c4dz/WIm2XK40aZJAW7wuasZURrOKkSVZhs1xFcXHAnV3nrbR7mBBiaI5BOKYzyEk7OoNaYrc3ce
CA5ox2iDjB9YFtTnRRkpxj2WRWuFxSaY/YxMmrCV4Y0o4UDXKUQ6J1ikXZjFsu4IMvrrW5hPZtUQ
2GXvbJ3BGt6dL5kX32X3rOv28Jg3syV9gF+MPkDnHzydzkGcPYAvzCm0k6SGHHw1y+DCW4PZnRg0
yg9D5FFlvOZM1rZM00StKL2I0kX/Zw8GElvZWq6MYl/qH0AtFX+rtNuIAO3FrlHojJoaiK3o3arQ
YBa+XvNpPoW6WIXEFlZth3gVvt1nm6Wyh3kPItV9UxlTLnCJMfQhgKWkRybOtmnuzJ9JQLxZm3He
cilNvxyjw6YqCK9MOZucDzb5xXX3JyttN9JRQNx2ox8N9aQQu3onTXwKnWRX6P3EO/FeOJ9R9fHE
M6WvmHCNB1OLFQkoacjBxEi6JXtSgiqFH2dTjCWsXZmnz6B7KLIuncdpipbCielg2KbxSuGK2oiY
dSg/gkC3BS13Cn7E9LQ+q5ENotqK7wVNfkxqYuzj5C7n0EOk2kTGG/+RpB13fxRSt6WeTAUDHm+0
VfI65f9vaU9QEsOXXRuP5YI/WT8AkxPzg65tgA0xLbolNrrroRAsKi3TxHXUOkoaWjRsI3oFtcQx
Vq0J1Iiqli4Nv/JPmnREJsV6eLN2XYoifQfUu5IirWdFjloxyUBEItPl5xic3nkvFakgvhtoes0P
BxlXn7XJmQ0M9g02nuus/2athfuzE4YkMZkhW1BnMSulpKdnZQErapvsvexneGcTDUmbfKDKWsox
SnJ+OK5c7gNkpO7noay4BXQlq4Fp1A1JpLo7OJ0O6JtCZIiIKXwiy/9BJb1Tsg2XVmv2vujF9WPP
eHvZj0mgrO/sBPyvHAVOmEMfYyTrFY/sADDnDiJEXOwjwdeA+uNafu/vza9d41jDKAqQXIoyIBup
fdh2vpwXAT5Id3k5RuGtVsgMcM05viazidZCgYNcl6M8VcLFmFG5NyYr0BZcFKTWMjhindznFlJ3
geez5SKy880FW0RTA9sQr3SUUt9avQtDztE3tYkS+BEeFoYoZvKausIM+I04P+8OywPFOfsnyv0j
TpDmm7b+3m6iPmeXCUMi3bekrqtCBLve0uVq/hkpwOkCvQGUGnOxszfPR7NwK1KM7IM3JYjD1ggn
i92qH6kxK6WgKQM5siFGj0bv94usIRflW5hKVmgIsuYR/sCASWCTFhhHseZLV9Q89ea2FKu7VbFh
HU7cF8zgoNote0vPWeC+eSOjwZW3ufe6QLNYGcnkzciQ78rr1VC2IG0yOS5nb06OvvEP1zxJn5Y9
l54gXGviB90rSPg1wagp0BdUMVYAJlGNxV76dtfYdjJK7hL7+8Muw92Z2XhzG2jONxmAn8DEvb/M
DpB844Ish6we9EExLmSfKQv/Fod/AqSYufiXYj8T7S1McB/hcN9Cfd6iJ0nHTsD0ErenJEbAa4oN
NJwLZqnB4RnjfuYO7vITYZaeWjmyYq8Xk6CKZhClaUN1fRCea45AnTQxgeXTMSL82LcImxpUtk7c
a96XqZHxQgq3Qf43j9GDJmEsMFaGgMPSnmrMqzCDtgEXOfr7WC394X8xvNP/t46z1WeZmbljBAa0
r9uCz3WuAetKZ37W+4rzckJKobLk39kUujub+hmBKSWL2nt/o3MEdfAm28L1azguBQR1mtFGsdm1
Y5cLI9DNNioGeRHm44K/+27D/IFUqjc/TQqq36nxJx8TNYM/QSF6H2Hd7lyWI6MP3AuIoY1nV+RT
FwV2RY6CQVIwSqmsVaNTySfC4KDhk+hnWybkK8VuQgst5J3AUI5YYdkJ0AAueJkn10U8BDpgIYkJ
xq6/X+grqu+hmu9GQOJ3rk7hzUE/ChhQAB8tGXIPf7ZnPkm9APcZVti/YTXdcaACpiZZL1XO17yC
lc7Lz7k019S60L7+fs/mnEHaGi/td7Rdn3GEy1URHolUM65WjpK2WrdfsdAishMN+0mw7lQWz21C
OBGofy26nm7G/Roeo5uLC6LWrI+vMNEezf3nc0u+J4ZOGUYOzDSTlRhpA/tshyI3s463RXU0zukY
d+PCLX2R3mvWsK2YSCFyXjXwzAWC0ku8pEKFTzYnjb8QogAlgo3focKrqsyU0WvH3D7wzIlolMeE
ypOlQfNMlmnjfTWubslj0yKhloqnEq1rQsrqCkVokCKklCgXJPy8cmYWpzKtjn1U1CNXI3qOD2PR
N4qZPj1xVs8aM95rXhoX58e9dFbicMTGFIGgC8pXL5U/krixNJGixo8IOxyTiCfl2hdzw0TyyFXq
MJA0IdON9mWrNg1Ik+8DTltY55v0790KPsZvPv8lFS/+OE0FZu9Wx9CO1oEbLfSh+UguhI2HSLZt
i7R5M5BZvjuvTLr+xjXuuH/4o11ZNtqDzzGIbSxNWekAjYjjUUgPn26/lCYMitRQTxR3ERnOXEei
3U8IKMjdwbvA+/LWG3vKJ1ZwPSErKC10sxwBMQ2BuFO6CAlHbF1WjU9lRvsrO/Esn9HVIqqIN/1L
mvG38bQ8HX+u9v/kCW8zZ3LuUvHlUbJi68tr4lNPJI+cWAC+J5IXC52nBCpm6/rGlC6D7h4XRufC
462vJrYwrtv7Orrb8wqw1wEm8dkHHFyEvTQeUvytyUJ12Pv0cDiWHihQ1RjJwG4P1jZfV++g5Zfj
vwHnVZlrao7AZukzkItrhDook0IPvTjtze3IiVF2seabajhhg0SM5PZF8wj1cKOBRPZDLYIpl6ij
105t7S17pm7GJ8KrcvbhqfZPQwhSRRSar/ANKomtPU53IHuqvxHaHYQ7msXJgTT+LypixUV89whm
lIvk/RxHIgA+N9SAf6hyAI8SgYujTP2va/wFFQR8HAsfE3I3Nrnt5fcpBh3xjRRUeXey5STUEJ0g
nvOOzPXC2ladNlMSZcUQdhK4Cskio5HerH+Th/vBIZ5n0VCDG+LzYJJoh1BuOLSQk3JePTAe9BRX
hSkQNElnEGAK8ABUaXFumuJLuzQ0I/efoShlwpPhrhPDyVH0A/CFlBzbPxbFYJVfYSksZV2vWWnu
Wz3QJG7prsel/U2vJ3x9WMoZBTaj8veAnwXBHG0ZTXV1GuZqjZggFPNaWd+7mnzD1Rw+LB88IXey
FT9PJshYSQncGcOKr8tZBYu3wD/o5e+aWA+Sr4fTCQYjuk6NQL1r+j6b+mqGChvVSqAUx0cFeCNw
tI2EVAuJEYZFsBY3oIavzY9VEXhcyurhQw3qOBirh1YqX0kbaOEUH0zW9fKelecXuomKKCK56gHu
paXG6zQGOqLuYLvfRccSBos6H/y/0rTMCzA2gi20AtBi8cSIrLbRE1u681NsY7QnchNhAyho/EyH
xEpUNKH31eYY6cE2V/Zm9tL53BROo5tkdlOz4LzWmOH8MUH1J2wFiPMrqsIiQlBCt1uVAxjY88R3
IzXtzidNtNVaDe5i00Y531WoggsTSwoL91yAGbatjSQl35MAJVjTzesXUsAGK2l31ucqsHMumfvc
emJhDm8YCjVZG3eOOKsGmAYvCsGqUgX+Ramw0z0SaKBxNFilxjyyYjZZtGTRGKIDFFuGBaFMcD95
6ktozUri6HX8JiyFuKjv54NWR/ToJ8t/W5ZJcbs7m0inIIlRNvxUciw3PriV44qK4QHBwr8zAnVu
q1JcRAazgyvbJLNqnbGnBkbrmjOgyOeOzTgijUyBZv6uB3JMujsoHHr3kE4nmJS0j5vEPpuWocQo
0stxMOQwive4FJmD413NwaQeT6753nNTLtwbHTi7v2mLcU3+sgrihvRmrTlwVzV+k1Zh26P9MHpH
J59VKfzMOuPet8UrTxl38XcQ9kcqe8EpUc7wmHL9MoYwKRIunB/mXu/j/3o+xhXbEPMn01qCSm2W
hQHsf7su1FaXz1DUOJ/n+SpHceDjrf3xxwYmDBU090Jizc/HFxa+UdOO7P990xfw+91TvUYVz+Mj
Gh3y3DMZJkaPDJKBZ2OxNqA3udZRjRWibRaxbZ71Ofv39IGbZqSDiVB62hpGevoIKxM3w0wXJSNK
NZ7yNYh3xAlQ30L0uLw97azBCsui9zXWq6+n9sueCKzrpklmzh1vViaMgmMw84ocdtVp4QlDYDXc
4YpuBBlZoGih56AX+8aEcUL8sbZkjifs9Gd3DeeOB13+vvD+n+/wjA8XHsgZBp0MfWzOniMsdMUE
4Qh8NMwvWWuc+vQtS74TyBynREQwAPYN0tOT86CvfhwlBQ5WI2Uu7I2viiMnNhHq5hnb5BkK9fMb
tdgfKFtFDp2cCvjLmnpuc0zw1LX14H+rW9J0Pfn4KVLhJEKQTBBJusA8kqYDdV3HDXHByEn8mL8i
VEOawAfMCW6E7+IHwSUbXRpmBNxgUvyOnFJ8vbzOrC1baTfpfujnw5K9EAxVvVPn5vpsPfF9sOpK
kKqQPKf7uJEGz9buXetNHwtck2W0oWHhjrYO2Of+tM0whkLxd1Tm3IhzZ/jl9ELij8Lf9JJTx3HW
m9tIssDuonLzjyvUoTLJzV9q1QjydwFaXEbWhp/OGlFR0VtdTRFcihUhoymWvSOcSkDPoPwOTto/
GDa5CW82daeWX+T320cTWspqf/31jpL6jw2R7UsPA4xe/cjpohJMt1e1RprJmptgqz/yV6hh0V6h
DYuY0dNc7GlLXP+KK65xq1EQyu/Ysf/97aXeOJQLhxxg/8PYp9ZR+ynIWh11iJNN+nqYboQytj6z
Nvq6tCwYBWZC2blJMPyoXQKrO5TudDcZA84lKvvZOQrslQqIyweLnj0jYs8flK7OUoFJ5qvGrdDw
V8Uerf17JEQpEu0HNvnVzD8USjOdfLfXkEtwOlmQOsMuQdjgUz1lVtgEMaWWJ46PKbdvY0cX0FJm
iQdFUnwyTEXW9pysD+XRLDn4mMJ7VJYDcPPCL3n6h9a8eyZzuzSE2gs4bUzkxpI1/RG3yFnr41CR
eqQVngO4nIEKhR5nI+QnOKm6/ydJxEtX7qAQ/pfrDKyiRBwfqvldnur8mMMh4CF1NmeHcxK61lhh
637nBFdGiuDvxUJzuDLpqL4NAwzfSNwX5iisiKO5OSYElIzf5cmSE7vtCqkzmF6hrhKz4UYn0PCq
ibvxOsl+hua6WGU6EfBfHBF+g5UCKOHBm5diqDi5BRLFmH1hTbLhUYCUza3llWun1d0Shl3/R6Z/
N5rhvzZBoo1ErCKDL73N2aNj6PuODNaWYKNdSXHG7nEyNVCK50b9YSybH2q0D/B5eodYRYQMMeon
BtJqLJCO/RWwXUK8pUx11JWnbYKCAx+x08djr/k0OL15+ZTPaovy5ITdQZqnVuVnkcwarXeHbYaP
fxBktyGNxeOE/KwZ5lx9nlmC0OTzQ9z01XjTIt2jLek5K9oj9+RCXJxAfq5Hcu1ltcsWdOO/DjQ+
rK+vRNztr2jT+n3wNvH5ITUXA3Ebl/rTowaq+0quSvPK2kC3cN0kLLerBKbARR9GQnaTiKK8wFA/
cHUDj7pzWngeY46epH3FQ82fB10v7ps6DuIkROg07jlRCkK/ZUgKAKZ6j5TnrFjwwYSwu8pAhGpE
IlmwIOGfTqVOkJ2/XWgGufiIn2l4th8zIdTEbq+w34R4+az+xDQrmrUpPsJR9Fblfx+6CjyVf/k+
tda7ZtFzjERrQ05K22RJHcS5GOpXGzbUIgQeOHeFHqeHdbmLDrRwcC2ctvDN72L0UfJDLapaLD9r
0+71GFi56fJ2mFk59YGBR22+9p3EclJBcLZjWqMFerRRwNYYQ8v3wBMt4Mhk0vGh2P3+qud50kUQ
8AGxBDRLrO4xBkmpd5BfGhSToriVQ8mJsJUm0reE/8ied3NqcE8lzmuhTIHPJWeY0vZfh224nLTc
ju+/W7nuSrYjKnvwZi/UwAnlI+vz+Q9/uu+b/+l3HQ0grD1ENACSoKBGfY1reoUGRnURY4pu8lcq
QUfAgDh3YJQy+CVJAcfLRvMWoTDSmZSzjengbKhFTe0z1oHdTyv6toRLSinn17BiU3CCo/3yLrGG
anx+l9pydEbxyx6ts9IBZLEeC2bv0z3wGiruiN9rBv9SQYWpZOHmXZRc2K+2b3ERdlBA7MeL3u1c
Zodes0rrtOCtWL6L48FWL5I9Dkif0FCXs0mPLGCBxl/sbpz0fORcJx/eCaDewvDPRsUvviCPMJER
BYZngLujJWEsxLbuwrJBjiBs4qGRIm7mv4U//p3NGxouGSq1l3VDtGDWgPJeXDvRsERrLgRKVJ5v
B6uI79zSx3P+DcfGd06hq61axLgdjjdyJPml+cMXT0GTPqh6A0z/D8127iu+VWCAn6OC8oxK50Fj
8OcfXT4zqArbzvOdFQ19jdpjs0tUadIQ4IC5QKSiaNomfbH+yDmNRnWQDa4g+ndVLV1Bp+gwatDZ
SPCzFH5GttCNw/yCJ5krspL2mt7ciINjZsibyMUATIq0JTKMAQuOjhQfCRfV0Xs7rbUNc4JgpTf7
tbiapXAeTfDKLq4wAZpDBB/fbAxpAga5LGhUvciPamtDyvaXuBH9w3CCjgPHXVPsDlJsKz0k4KLK
eAwtFnIdkmofOAfsRH2awHXhQ84fCQURID4D7dP01ESRASHeYuaYU3K/WcxdoFmaZh14Q704AeHA
Yf5vUEhM99VBmYSI9YhrK6syDYYMCQPboylJPDKTsTBUgvSusJ0w/AiW3nePxogQ0wIQekkhFjvh
c/KZvi/32osv+a4SvwP1ru2DY/FWwyyZ234O1pOqFJHyTzq1uCGR9rh/jF11CliuG8rybKsf0wjg
Fn8TAnYQv0T+IBoh8fRRhyl4qEvi1GkdQjUz0H+uCn+IyZFu2g1HCdBar690amcde1stWfCPphbd
n3Gb4DGiuyade+KfR+UJEVTWssaZk9wZbq9coTFRhW7uRxf3DCJhhrXl+5cqXllY3mCWffvDkgER
4Qhk74hK4Is/oYfinCz0WCfBfBXTzrpclMPpO3v5daLh9rS2nWyMWyrgP0aUUw1+gmXyLp61uNQN
AduC5+jwfXrUhgJepKkz+VQpxx4Lr+AV0J7q9OSAeOykgQtAsSGwmeE8g3r2aJcaNP3yW3mNrFig
V1XLEfvsG8oiu41pva1QEp9thhWg3jbDs2oxBnesTywEry/oznPL8EUgDeVyhaVzbmD+ek7bWrlg
IlQEy3Lqi5ymsGpB2ZWNiRzpdbHISqZEfUY5CRizdHTVRZ2s6YGP5FMmDdJpWN9tRPzOVfsawNb4
vVc+a+ntXdT2hFbvW1D74MjbcasJeL8J/JljwYNGu4pE2t1TgcdAynJ+r0zwnZ1mCLdHb5xzhfAl
EP4jriAGBgI19lGe61PacDyFHDkR1nwmCkksqrDoMDMOQKP/LYfvH5BluLBA0DmhKHW6ynDiL8jO
tRAkX76yrek6tHOX6XUFZlD7+OVU014rui07v0aUNN9ublOYSc6uW7r/NF9WyWwGwrbdLKERKG9U
hWnmrlXzb4jc9RK4Ycq3D34hKMvHJPsOERK0CHRdlmaOywsL+ThIUJMuY4tiKz/82/bcRB4fbTaL
BO555aararvTysLHO3yUUt3nWSF4Hn1IWAwLxTXLVY4v4ppSFlpdU9Q8B8MKdt6Ett1JzSoinISz
sjplDK94QFO0FIkr7xyB6VOeAVzdaGSK+nAH9ajvbH6VPYpbXc918n4oZpNikM2hlmABprVz7h2s
hGBd7h1uiD5FbwdtUXvGILOVVt3WPvRqWRw7S5/qXZ8xs4RlMncnS3jEFa0cTLtziAQIdx585Ot1
84nNTxFxQI8jFhsUH4AVRFDVoQSR+GJSXqaTHbjriHbz66cA8aumrTRaMLW31Rl2+phSIYC3lR/3
G4Q51Na7RVpzUKx6veyTuf5f5wZ1ocVw8G5+qrOLPciRtiUkZDoRCKKyYj2xNHwxpT1s3moGa+FI
ejkYzRDTI7PiTHOUE5m7uEGAXMqHh4dKfDzQvUG/Y0Z50JFYH6igKn08EntG5n24AyQE82e7e0Lr
oNsYW6Mo8nAqBEyuQkoPqOtppDsbPOTFRuggQkllWsP0wV7oguqSMGs3prlQIg9FZcBnw2RA0ciM
FC3+eHrbWpm9rRvrvSMNb1toqi0Cq3GD2fUY7PrnHRMx6F/nu9du4CRkMt2Du0w7zxPJkfqhS8Vv
+ipCB7ofEH/JQe18cgMxEpmVLeD5aBevogxed6xQDoM7Q1AEn9vyivh2+jOrgzba0jP4IWMlt4MH
qrf2Jnpnxdoua7/53ZvTNCs6tAuTjD5qa+tNgRqKQZ1d6ziHTUwrI7U0e5CAIiPPzQZ1sODh3IrQ
WVWHy1qt9bFBSCSD7CJ3dhiJNt0lQtWCTNDsuXVkgpfwO6Na2EMKwKkTYXYymwlitbDQNnWT7GLM
j7Qq7XmlE9GTMKDUSgRwI2XsMpE/q4CUrZkwYomX6+efISQnGYshrioLp+Sum1gY42GhFSpEA5/8
bMjJSKroS76V/sLGLo0yiDKeY462TONuSU3VdMzJQGVu+jNy3vZYbV7CtIctP3NiTUoOMDydkMnp
X4oXIX1OfHLBEgWEFW6hoD4uwyAtodMmHv7DyjadD88kgB4uTcnSis4mrGPLhhytYsbEs8XKgCwq
JoZvyj8dgzO9gYSncOiRUdYNDLcK6UCAX31RO9R3ZAJSCC/9DEWpNX7GxnjCDycVXZs/FV4TVqdw
trGYMFeCF7b/9iRGQyVwXT5HJDdbSjBmQ+ibReBIZV3IeZzOQJu3oDxwln8VFdSFDeclUP7gG94Y
fHfrG1QSIar50rnjERz8By7+oiv4wReJyTCNF2A+xbOo2Q5SoohEICUoJsc/mL5NdTQu4YMGVLqZ
ti9UhOQ4dF1PL1ovyi+JgnipEel5rzlvdMb1Yp54yhImrSJ3RoqJi9yrakSIEkCZoBHSxHUZ7VPj
ORZ06FG3pauT2bReHOZYwsFS4B1o64KadxX5ir1pjFzHhJlGH+gV8ffV0dsu10X3ysNCjcxC/bzm
GNvWbejR87YXZdg2FTaytTGihZpImQobUHzWP41HBSDPm8sdEMYSTQZUE/KCmQ4AmTnsA+iH9mmb
H0JRb96Ix4oeJeiY6pPjE1URdQtilFAP1rRB+m5a73UtHPoZWuY4LAm3A5GqsFoiC4qdEpixwZy/
VJr5leefIfM+z03huLJA3+ajhHidZwe7tPOenwPGb4ahdPg6bwFG0umRa6cQ8Wxrcvj4Je9H2kvf
6FGRKfCWeHhJY9QCwKhGYomAkbyyh8yRFliTBi/B1P+g34ZZZe/O2cduaRp3w/qfL4O82m2tJd1G
vfFbWcaYN68arG9TsdNNgEoeHTJzYbbnovjjIAAjV/wm6VkzvpnaFcQIhrfGKYYUpnuJrc4P/PsZ
hYhQlO7MXo0ul0QJ34QQ1P8rXzzVytubVD1Qm2ms9y80PKXxB7cIxJhPKy7gXntx3j92WEXQDbGp
j7YcsGErBHFnVUDIKb+iw2ncQfxGuhkZaRpq+f6GXAEUOUtVLh3r1xYUfJd3HxwcnGK8HxojkblA
2FR+WuoQIeJ3+bJfAfz1gO/r+xGuzoD2l9g03PWwEfhtKXASMYFuPSQErvZto5HA3FeUxFvMPFb/
7CX/iBojYJXQChJlETpEHpCsfQIpYd+osCWXIiZAux/iLbVs99y73o+9h6empYjtuBnHufaOjy17
FrbEKBF96vGueRq8EYv6SuYJjGv6sWnPhEr8UJMf3CFpzqWXGFVFopjcivFWuahDVGJSHvJTF0qS
C6i4JSckw0fBfH0AQtEu0E479TH3pjV9bI+BRUQPpYMiil3XVD8O9k0Ilcf8TUu5yoOk8cLa/qSU
yhMpsUUY3hQgoPS1JTtJfjPOJoiomdjU80z+Za6KNYH7+bIprzzIn8DbFVs0w/vBDp3Jmgg0on73
i/vBLbr4zFajN/QjsctNumgtEeGGcW0JM0nTnqCgI6nBeZuK3nmqcci/ijprFYCBDIOTiIITaLVA
LnOetGbiZH3zj3nHU3d0VehweCVLUyH0OYrZgmDzf8WliCwvtNXUR9RLs0xn/QcJVyQHHR6aej3F
cga2RPk5njkkRErITIpGPK85RfpVnETMB++z481q3fQwYFXomawR8RuQ6Jq/knuNdUy4Ecjkm3Mv
MHkuPKgSZqo9Z6ZH9e4Lr0GMFyFH/wSOiRRoAuB9Ea+a/w5G77OAdcnieh5peFsZPR6l5FKCU/C3
hdFVXPDPE40OhzmKCUVeNnzohOl9BGWs/Y/GJyai7qG+A/G5AV6Y64PZYBlmyxLlENa/LsLii7PX
Y1U6pZJfiLG4hHNlqKgIGmoh5fRPxHviCO9jqbjRhGsTuIZ1uKtrNNNDzLsE06L7qD0Ej8YuATyH
hXaO9XNeoNjL6wW1KgCbak1kumytM5oQspDAoNU+CYaQScYtFgaBW7l4m38V0O5EMDq7eqg2UeKH
YPbOsxe8ZpjAawLlo5ynyNdLIwP9KXEJv4XfMXzsWzBYOaOMRNhO5hEazIgPuBaVnBxzc6SQdCyo
BtO69xY6r9U7eYEFnVtfNZf6t76jzUPbMTo6lysw2cDQv7WD3rmbD8kB1Dhb2yxRQKvobh/LWnnl
YBPGPLwthirgyu3K6K1ltybycfCUdsQVSTdMQjf/o2Mbl0QuIFyj/PxCXpN0F6Oiovn1qjjZne4+
BngI/rWxXEgNKYTpHJdzUMKXYnQh9gky4w7iOLtxW/OBQcHiTj8XgLppG1th1KlK8WeF4JOJQ7g/
fVPtx2xiYT46NcYbdmDscZXIOK0VSXdR7Wj3IeqkDhc8WTR0+l3u7S8eKvTRgdfSf3HeVx/I6WTt
85PpHLlGlAoxlnZl5FJzyggSNdTKeedKjQubUNCd+ozYRWU5Z9fjtO3XbbZ4IlTW0b+4qV7soaWc
7oC2af+F7iGGpqzurD7tltEQwZGHMaQEe5mRaoscvLC9W7DGkpINWQ69uKENvQ5pPIpbhz1WPO6T
QdQMN7+oIoMrBREx6VraZrzNGE0WrphY6/5xPK/ZVy+FGygzulnJ7uOk6L/oj1KueRrHOqcIwJL8
dQDRXXIIoaKUq17B+2N3EEppxwcRfXUlE79LYBPh00YMQf5j2dl3jCS0m7sjKEf6mTV9rGc/LESY
yCW3ju7wqDucJdyslKre8hviEegHn7ipSVYtzEkHTpuObEUBaHKF1YV3NdtTLFOMCoeXAYIOqnWG
slp+uBJlkQhUbjFv4EZ1u2gPHboZz/znD90ncGPaY0g8YNxccNCM7UzEqLpKtvfLBFEYyN4pFKBy
BwhwXm6CAUVj5F0wiBDOZW+vs7sSBYlpu2lCcQ+z58ZF4WEtFOldHDs5dVKi2IbMMqIqL+F8IJ1+
JeKL9S7NFftxSS7L9q20KF4UETS1byvfCgDgCpX/KjuWxUFQ1N/tnAY3QPdeQJmQMp3qFYlx+I9d
eHSp51/D17QEISUCMxOBl2U4j6fFIgCD30bh40V3cmkbUDDIurWjifRbtAzJqwHowCLNBnGnYZiz
6lBN+Nviq90IacSxntZ1cj+LUHnI+mS5twuqQ2zek94+BuZSg7En61uGzSQY8b4gvgJLbP7315jz
bFQGtInb3OCf7j39M4znaD2imvNMFjU/QyyBl2bZ7h+T0MDsclm71a+m9eY2koNeOHteo8pGJu5I
xK7QBl0nh9GaX0WCkJYLBlQP+2D1RU8mIO7/vmHCMLQ45PIM4P2UNKVdUYwS89TuxidfvVYUK6wP
5r2dRGu8bFJ+wreK0eBv8DY5ZyaqH8aN2lVNGmXsxv8kHVjnxS3TtuHDCoJ8VqHmiDI0s5QBrbr7
fCtr9xMG0hEEe/84UQ8URWHLBfjeQEe9Rn+88vn0oYPL84wfVhDs2OYV2NeTehevGjURm8gTnDSO
K+fF0G9jLtH7ocBpQ5JjlMI8EpFQV2cugg1nt7y4TVUaLew9lLrWLDLKScTTBdEzbKPWHhRJa13b
iv14A5Yps9MGFPn7Qsts76+n7GaLmolDpJc7tNUdilB3XRrSmsscYQTJUVy83zDVhWv2NemHkOyr
3Y0i4NISmmXPnkX6I5pytK8lREP0N5UMqdkfUh6KeZrp9EZkliKYJZQq+XStgF/Hy0dZxMTGfm3c
+EQQvmvFnRwjdohs1GrIAVQ93b5+FjaZ6Cc4MsjfsS/V5rFb2CfH9tX5CMAPjcKIUn5TSC3aEKYf
w6jYs4fH0ftjh6W3Aed+pfFTfRb6Wrpjvn+LZ4HV8koojEIqxtTDSLhdE8+CMd6yi7UuQSafo6m7
/FTKfCk9i83Je+TIb+RA/S74SqCXllMHkX+ICEnYjXyUJF7F7wiFRegxYskbJfrkJxMda4hhIE03
UFjngh1hPepjdOAY38Ntt1JbIJsWJr+2FsQuI+0dG4oTgG0EqhBLEg+hRh4/rlEjVsahc2cwuS9+
fLD7G60PISRWb2ERE/fCuyQLe98Wi10+frFfnumjAdJd1Dk/WhL66wWEXEqw1xwZe4KOToXyQXiQ
lszVJLzUDDMH/DWKEjV5gKW9EOwnHR8g30z9JTUtnzc+tAeY0vD9zb2jejnRkFWipQvIyxb+12kD
fqwX05JB/RGvLEOpeZIrsZLkHVAlvtOdRZ3+Smy9DYCfGQX/T28a5/eFZwM+BtnPvBq7oJgwbTe/
lTmOsnhhI5lXmufj3ZH3oxs6Ak68n4xvlEFoLQXkdfwMrubFK91BeCHNvwBPTJdslNFNAUg3Z8U8
8VL5xBRqVa9jzdVj2VPVB6R1BDZ51cHSom1oQ9vMBsD8PvKEktQS1CC6b3hCYqJ3IdiFO409dk0V
/wDiXRmCLVApa14VatYN8p5LsmT9YPVO1H7K0LH6jWNNZSCAqaMo5GWZLPJolupFtmXnWv2m5GpS
f6gKi1DQktQCEdtG2Icie1oLNFG3RkqK3nAHSd/B0d+33AFTF5fqIimt2R15iDqDvTTT757DR59q
9OlUKsXJR0S5XaPUdY7XW+RdQGvNj4fZe1eIg7NF/5b2wbzeaGEwUgMIrONFng/OKQ7LrJsT+Tk/
PLyOQrY62AC3aQeDkntkQbmkWVbBjcVMif3Om/JwgJJjjtDvqjHco+khjiMr2NedaUpaCd4byJkS
rEJiLtdMhqWr+CE/oNwVB1/9C0R8CvM9RrtgqgPVLmEEb9eSNlypUd4xXn26lXlEWktqJjFHCLzV
xAazojhQ1J1Li/1SfXpWLMlodLFjzVUV4yv8dHh/kW0Fe1/Lo2cdiZMDwMiO65n+akdD2q4PTwCG
dU2Nfbbm0I4/o2nP9oRnkVZmNg8txm0nKWT421VwSbiZKioBVzLz3tkqz8jE+XlveORy2t1ghI7D
IXHNdTRk/NHcRMBk8w3clRPXNRCKCnRDzMa3cCcGarrOVJmsIWjKGyVWWWiBVfiE7cDsjM5s+h+e
vSriL6i1/lwcZyn/Z3Hzf1R5Rps1RZLMRTOuooin7ocW/gh7cdG70tzLhn1eBJnFbQyOvqsVQi0z
ypQh92lWsRFb0dQ8fBkhrc/Ho/WiuYfkM16tiVFJuOum1os7kOq06K/a5SJAp4Srr5TrfZ0KozWD
kso3S/GNU6WLgKyXV4hnlS7LE4KCoUn1Uc5tLPSfiaj8ApRszkn42pgJmQkGqtKKQN8VXkpjMI7z
t/tySsOd8ou09h27QBSjqGKPydlS+wtTHFT10e6rIOKfwsNzcoAq2mD35MS3zTAJsDtKnBUcmBN9
4evU6Z+jXM/qbXmmg3qzAX4aiqwqsWtKX4//+kSzMEeVNwjoEYeWmPiV0UgQpUufrQmQu/RJysMd
ysN6R/xVw/RqDA9kg7FbCBcYVy919r1E3R5FcS1mDnk8b1j4u2i69d09/nfWiVzkGe/lcQr/+P9t
Ne1bzhBpFAGb7FOcAglnlSdEyqhlhjL3w3zeCR0Z2a1iMNfXmgixHchlqdoNbGo8B4kAPgbrCHBt
5aGbuPNsnEYqMHXtJ+zwpkSBiV6fz7mgyrALNfc9XR076OfDEM412DcM7+2zJyonDGiX2mH0z4Me
Fuxd/WDgxfLHmqLu57cR51t5+o/A32/chGvQyFzwsTyrhZtj5bUQafZpaL1EdVcUBm/thtd4uduH
KAph1g8S6dwte73bONKTBbm/jOz2WazPKXzQ4YCzHi6klbQ+UrMnVyfrvl6kTBJgSthu3c9NV7e4
DdphrKSMaBmn4SDi4F9IFkj/LuucaLHxqtRMlEVtNOmegmzTKYkib1f5G1GA8OtX++vKkUMWYyP0
KuQ5pFWksP+Pe0E8UEwWgm/mewR4JiMjq7iAf2OA7g7qUnjy7WLKnqfilEVlxDkq0AvaDS3beheL
ZsqNXecCrXXbxRLXAd1Lz8gWNTtW1C8Dqn9u0p2sdwlqrs8hU7hTFRK58w5cYx4aaXWnaON2d8+C
1Jygo+d79XZIc9RAjEK6uTxvaXhoZMaQm/ahcyF5B4422ovmW75VYshZGfkmvD3S+ADt7gjXp7gE
76OZ2Y1FW0dr+oFrN7adnUm//BJCxURBOf+LkxwJ1Fu6RPmiccVVCxaf0ewQuRQFZuhVkxYSfqHp
7e9b//jbgAjgk9Wo4sjm/Ud/Lr3HKNIN1XBerRw2M8vaCEJUYVO1zb9iB/qQIzQN9jiy+lUuGUAz
2TPPBYRFK4S5v4CF+jel9wj1Q37iDI7PYJhC7TCbROlV5bEDXfoapC225H2xyzPnkg+st70DZudL
vmBJL8tX+9FzFl7R87zb6kfOBU7dXgAIxAdv0LXLwUQn6hMSvEvB+CT8SkOOT7OGYfLgw3JTg02R
4WJh5DaNMjl1Fu52Hc0XAVWTRmqqRJF+Hj+EvCuMcQj5JGv03UL5xkB5kO09jrQoEwfA/QMdYl67
tIUU9HLThSgkfmrUsZKX0XlzF9NRa61Mk7WQ+buxIy64ljQgBCbENFCrk4dg6jnia5okOTbEYZs4
GaMQvN5ez8VB2aU1fOYYW25xC+7OLMQrfrhBjxvjZQaPX6irGXvlJBvp+HwtfKkYyJKJtYg/WiXP
1L5ISyUxbZja/NkVZTcuQSCUep+FrixvNNfjW8rYMgKthRc2WX/V/NuqYH21uS6bjJUzlQ7T49pF
ur9oCBgfOdEBtiRSLuAFFJOQqGAIbbtUxnbIgyuEUpPYhysE4RoqWjJTJJkFKibZ7WaFLKQyc39A
gJgOiL9W1RP7Q7z4sCy1Z/KEkBe3QAoDGNJ1mtJ+52bk80GTsW2VfSTzbsnuy4GztuWWfBHGlx8J
DCwU81GWg/2EVujouZzt1KoaVU93e+XExzuYQIP/cszEATSquJ50v/eGJDIUmBmOh/uouFo2L4Bw
4Z9gfcFqRWpSKv1HqdcbE96WqWwlJ5DMe4eEdpioXiKIpE5k9biPeDuOR0QcWEP7ACxC+S1yVR77
FPEavvTiakavtaXjMyu4OTnLNK2uFk0zkETRgmVLDAFg8/Iqr23PaQC/6HFT7h5N/JLJ+3PBmM/J
Gm3mIX5/TVsv1bDlsbZ/qa+gh8ugQjMWIw/lssLcuqRxE4wVaBF3yACi0/tjUchDVaq2GbRXGCPB
X/8S2Bs7vXKbw1Fs+cj/fVij7vvXSbU23aW8+p66iNTk4ke4kzpfGEGlICthOWyIZpy0khasCqXK
ojtnhB5Nv3WI5BwgeoTl/oz0ioig2vODsXDOijqmdk9boIUnUbR2jDB8CUdhU125IfBtiEJ8WQWn
gX2gTK+pf4bDIt9Fx/lKBBnMQRCdKKagF67SMMbKUhs7LqXSf40JFHSHuggcr9j7zdZAq6iP2I/Q
sd+ilp5VwL5IDw2WVqOZ7jvmhuknb1JAwbg0skWmDkNjNDZU+BTPyEIhpWwB0N7JdY7cw/p79bDZ
+ZR465eXWeLD7yyQMcrBB5t9S2v2IJIng76NKY6YtC1tkGX9KuYYBzMa9prts5z6OD/8EmtNu8Da
6IFYiSAPMp3NMDuWkuaE3h1I+jU6kfA2gZlRy/y/C36h0bNJM0kUdccp/7oOmm0fZCFz7ZiEM7Z2
wXHym/ejp+BsdnYMp/37ny6av9ZcKvTXV9fbnaoiwiy6J0EI92PJu9gE/MMnDZC7Il89eEcKeKRs
ohUs34k/FZOfsZSxuqqpQLJA9HHuvcbG2ed+uDhPBnf0BvW+zF1FvFi7jojjxQAhPk7TUOOajtFn
TobNOTGDgwCWaie690DDJa4VYfSLpQilcQ2Cyd5OXnktCu1gvI67rmVV5Ag2yTxwoKzAjHUJJrof
gglqP51zrszN2EL5No2VoFe+B8kYuN18zNvLoJLlWzmqe+Ww8P2oTr6B/idyQzPGZCAy/kZ8WngZ
6aPliESa7ePYohQ8zS6cBazj6lWd7PrYSYwsj9Z1NIsYhMa7BPtx6cxTt1eBKl3UyX8aWhIXP4tZ
nG84PkNW+vWgW+rx52CpSohBanXAqoCTjx8xH+ZepQE/th9aHnpBqBv6JOjRpqds5bbOOjeFgPAw
kjNjF9UAlRK9EoitDmCrCi2uauN+eqRWvMwX3moM4FINK91X2IoKXqN0y+EHeK8Hom5CpC6J8o1Z
PgPJIhL2+GsNKmWdGlXU3xpn+biTDVcV6TKet7VDlnoCKJR1TXB7p7n+LNu14b7necgixenRwYDA
9s/4hvhZ+jGqj7wQhKFxy3swCt9WKUUkqWeMPdtnAeRraUnWrILlh+ysK+vlrXJvEowNP4feEwfg
oUdJ1av/DiwA61uCg8icFmn+k1Zn/UyMixtd+7FZU15npeyDqMxxY4ElRC1Xt25kUlB6UWVjZAt4
f/PWolA8TXi3xwi7VTLKmUc1MXVB0SVvs++8RoWU6JZCEVVZUYyTdm9DVmX3ROj5BO+d8Ob2VKVU
OGAf5yTUFfaItzLbN4xQFmKfSOb3dXQOfclVd0PUXFLMnRlg44ALzVV57NRkd9XI6NZswK0go0/R
NaXisMdNVy0UTioO5qUirF9GZAAtRKhFWBWlnuRp1/K8q0hRKZfVfhZyajFGR6TcHMr4xo2VichN
t4zEAhQkymMQ6CJSnjdeFWebIaxwtqdhuA0OuDzN9QbPXMmPxO4MgU9eqlzL2i5IvTwdFdBX/UbS
aY0x4HlhN3e235tcA9UQnAgrtpgL68MfVh8tbsBYGNW/F0n+SQbYD3EcB6GgNQsyZ8BRrDlSa6A0
6SdNBLHEvlrH+T/c7AOJ2GMbSs6lHfG5RviZyYv/FX+ILBl6zSWfNLTgRTKSnqcgvLilL++UfgY9
zspESjupHiZzE9yi3ASYg2wsfSa+JU8WxkVhoaEULJfgOE5hBsRIvJTu/fNUwihqrI2jloamgNxz
9yTk1OYc41x9UXittNOpp+thoGI9u+B4Kunqt2DDNEEXmb5pXsSvSk2gSagXVuKcI2mznLDQZmNl
DsIILi+1YFhLkWeVOTPnsiDuxFV1jA9RRkFF1YoLxhHoOt9SiNkEZmHHsG04cI12iOoNnY/8Mu3P
EBFKRUx0n+l+IsRSeaBSv1GGmgsZjzEEuVTxfgyq0lXqMFexiCe/SmDHwJtGXsBds6e+nutIFMhJ
bJ2vNxjYY5Qx+Hs60Kvnn6C/dTa2CRoSDo0AlpbCPwZOBCJVl1UAeDL/HwnKLf/r4TT+oxbDqqRn
zwp4LB9q1MzD+UuiUEj2Hxm+rMpK0Sbm/9LYvSm0P8SdC4MnAzVcj79obtBAaPGFm2+ZoNrDXIfu
9GLWZeK4yByNb8Bc1oZxDlbl6d56a3cZLrJzx/zJ6QDzvmU81oNzzUhSNUpYHkINdcbXza7mCDvj
xKn8yGBx1TixDUaMC8AX8p3OdiAhON98dNrE4pQC85Fmr1S+uBTVlvfV9d7XTBxnwz0UiQE2fIAx
opP1ABoVVr7aMCcWbnvy9NoKmGl6sr1yg4uM1KNA6XcwT7/TvnrMGPfdHLzcjGKfjbMeP3c8Sk/k
5SMBpFMy4+l1W+/3kA3+X89sfeDu4LE65IEYrIp1l4LRp9u/5X4oNo04iim1yDk7BGmFC7d9fP2u
G7EVMUm2KLqh/aDUyR2YM6sZgIx6+OQJvuYhkY+ImaCXKaf5oIyEY6WBYwUoxVKveCQ5FCRXjUK/
p5mNJS9+kRARttbGG0+JzXydth8yOUxSKXEF4cfvEyP0N8w0PNnUoorheXUwN20V8bUKIVA4poug
UE7pcGM82K2ONpBxow9iyqTKfzqYQogJ6I2dxrN3FkCjCjJkPGtlMgaOu3XdOAf5oV3zlYkHfgJ6
374qnn4WuOA7gP1Pkbl59d2Lvr3RlivSEIaCYgG01v00YCUW8gNhuGGLwQfSNbH0IhtOriS8STrA
qkvk3Lz3BNm3mtTxx0mIxP8lXiTOm2YD874llPWfImf5Tafztct6MJLOlGrcJ3gapMJsj3JtM7b/
NMeAbRgN8FtWy3W3/nh3XmZG/3dqnEMfh5n1bn+hGTIJS3VK7EAt5hWYAapt+8bq8tVMQeJQtqRr
6K5MM4wdelfBYl0KffHHXNIKU4UYux8VCm7VHxbWj1z2H6V4HP9X8bzIkdLy4kOejjAB9VbGQtB6
LGm5TIH7Odv9fQRLaZcf1W5+f2lEe9ECOl496GAASMwAKkXEa9enSj8KEb4T0m+FhZfMkbs1ZWt4
TXACUm0MfD2xQS4kBU/Bz+bEZpzd56R4lEyuWJtEu/RQUDw6K8JiAkT/9C+S62rMlF0IMcacvF7w
GXKuBdSDUdqx5ic3vsfo5nbguWK8s8EUbmltN179RCpiWx42FSB3sbolBtD4Co8c8JMiOla3FaGW
+Ynl9+wOD2Zrhf7GOYHLTtL1WhVKhTTmSFREMJdRErzlFNvkPcGqxm6/TjvsxxagvnDYP3EqJ2V9
WC/x0/ZsMGbaqkP+q1x+k1+PtDqtI+hfUVauHDdzutORN/xYhtdEB88NnDFxq9FMTHpOr+0MDpnx
JSwY1kUivTWI9r6os3oFK1d+Sor/6Eep3hLcbsGyXKAtZkbTsX7DySxLIlKOpuYtuuIGZykZ9SBQ
LpAdoBtjSjPvH5H1/Bel6jIP7BrPMJu5WJnPLTw9f4jvxNU72ZPReO2+fERCYAVcra+YMzrOBXJb
IxtcjNqRQlebckEerbqruTh6xnpVThTTfAagK/mq0QsysXHkuZ+FHiLakUQJcFz+ucDLA1E4uMNv
FJYopPhf/kWkAlj1Uji61/RyhBiVXESKB9WheylHoGYUuLWT+pVvIQ0v98+BD8Fm3BqD3Ken1CDy
8j17qA35yTmNvwzh+iO4yribqwot5ZluuwOfJXhfZQY2g6PWwJzVEjsAaDr6g5FuN919zhqW917G
DanD9UJtdFDU5zmayRsir8D2DRdL+hAxRohICuFOV/mh/qNQJttW8F5/89xFMM+ljSHuHJ3WvTSY
fpoJvWfhet2LKJwRJiN3/DiFKbFIO+dePMA7u66pbQTPdW6rCRpWwiQaXqGC+gDdniWbeHhf41It
s4NDhAPguBeeG7TQwYIPm3YVGIQH8GMbmhQhFOUnPpnjvgbqtDG1Vou+P0DKgLxO0v33QBXZFOUv
gEbxZe/3sASsjCKm6yFqJ+Bm/Bu6Wlj8x0J0wT3NCTfha0nlq1EC+EgJ8DwjDW/rLXjiNvxY9W+I
pE15FkKQ94po/LAZd4SHTie36iZ3sdvTvDV/uf/6nKGEtHYx5gPN7M/UAQqZd7vDZteFiR5cqMQA
3sFSDHhbWF26WjzylgfTuzbsj8NXLib5zy1ZKXhc/yb1nbH0hi1WhcGZAtYC/GHQ3WWUra3R3RCE
fm4PovT+gL7C5WS9+8/YNlnIeAMlaIzWgI4OQawxSRNsfsbtluDicHlLM1ubBmzvjzoD1PVVoweT
nNwh1uO1gxDjLsJZzOLkOYdT0cs6CAmQgFHi4OxevITqW26aehFNLxOtM1AwITPZ+PJski3Kqlf9
cDXvxQgVbTLdof8htvchgg2CES2onw0GWfxv9fxA5qTpyJqwZC+Ra7Wlr8WJV3CoP4g3nx5uqYNo
hCE/1hf026WO17RErTnQmUeUnF4wv0V27TzdYXcE8tUJfQujYHjiNvTiTCT9UoG+LCq1xZg1lXKG
tIIvJIyKmq/ZLiKQezfaonzACHiPoY42YjyUMtYUxgTWYF+PUlAujt9RtbVQ7mxG6kxe3g2Givt7
ItJlzOxA1VFFcLq2N9o3E3Dv398SorPnEYfqMd0xaw6S3VL91kaQhVazSkvOYjdIt7PUxeLWoLFl
bES8VYtParzzhtjt/KszOkBNHG/smqcD+YeoQ3uKlsjvHiL7jrn+Vmp2WO/FfHhZhEU5xp793/CA
PVhNuGV7h4woaGzcYwenySFA5RqZoXbHBp8PWuq3NO9RsNvq7bY3emuRNjQxpXagDY3w/QClm9Qx
X7SCXAIDXMF9Cs9hMumGS/tRd0ZJ0PrDbSsZm2ttSkxNoFQ9i5zR+fQibkjBxAxaMttl2+urUpKq
1bkpRNVnpoB1pVhjhcEkaSz76PVkFHtbQDIwKeVr6noYf4SdSgjQoiiMZ3v/tVZavXDJF5erS3iI
jmvDNevpyCkm6rg/q+QrOIubTJ6NJbKBEi8gdvJaV0AL9aZhFBYv1dmf2xSmXt+7Bcz/NFLeWqpa
7kxcnY/vS8qfW0qU0V31gY2d+5tzwF3oKyIPYUpI5jV4Cr/rRNjwtNXQY4qfU8p+bu9aoKAYlyJP
mwh1CYUom4WT2NL0TbtIswmz8TRcYvPwRAHZOW0rpaRUO6OTuzTAn/K+nsEkfcojr9o43+/PwYYS
FSVsl82UqaKD3xH4pqnG0hiXXSKGwzNeOuhEwH2tuJZcO1NEhuFx4HP0/yMybGmXJs1cnDY3v4R7
ZUkeXug/BBw9QYsmxnpXm9XYXkQ4qduKhHW09qR0Ygm28ycKcBORMmdDmbqiUs9CUN0YI1whLb/J
FEViDINPyN8EzS+WFNHq7mbuI9JQ1ybOqAtWE9MahPurFqiD8u013ZryPianXa0CKTsVvlQmhBsV
rXV+Pk/cX7YH+TamsTYufENjN24HGHVPLVZYw2ciY2ti56/OEKYxCTARFsE3jo6hzXD03Nwhys4h
D1aLaMr7itWhmk1ARdQ5PaB4YzvT6OwysbRr36fZgWn0XV2+7C8uLJGUFjmgfm9WTEGGNNRk2izY
BKfOisd3M7LsT1CC+0kOfqt8DOPrQZRPjRTpYUPJpT3In+TwHIbP4PqMhRRuaXIs4hpAnNWdI3jV
jiEZyBNuG1r6DqvTNNydPC+8FacL3+eW8KbitgvQlsMgwbIci1zGWKkDZall042e4ySJUnJSY8w/
dhsNInjeQWRsctcwcx0WSeZ9YuTEd4UICr+oAx5RntpLfqaWTtPNx5LcVqjCM5dPF6d+kh+53vgd
Gk9kyEVxY6IuEEfhwM9d2x7FqaMEE7FDCQQPOcJGFlEvhhOz1diSQqmXvd6b7n6bSvG576zgmhI2
vE+13yJfHz7+Q+4ABjAgnHmIayEhwfF1TUjFall6xuXZOa6kHA+EYUnqNTfcspBQuE27cIpcaFot
RS8LiEgpCUYYlBVtMWPE2aP2nHaW1NpUG+ySCTcZo/EqDPi5OahDjXQw5ZzWZiFqOwXBWKC7K3BL
oVVtGnViEMflSn66bNuNLQEl4va0EIgL9t4dh7wtC1YcW335k6y2ci7b1Fbnp9/V9Rp4yugiGcgC
socQSdv/98y13CAW6kFVgFAjxG8jJ+LiHmhzkkiHuevS9Bg8kTRVeIwYfm2x3yFmd0CfAqVJTEVI
Qn86Ie86/QF5Tr63cf6q5LcxFRjFVxuOlf9HEfKZhCBE0pl0T0DietvVcL/Wcho/yNoiXCADOzBd
lil6F5cXs3dfmbRLLW/jO7ITUHYnTC3/44KSxozdWNR0L1hbTOWfN3hlZZzcZQeunkwZRKO7wOdz
cKtaDrvZqD/4sb76NRkbecd5D2XXn/xw2eAhF/kirn/bT80x5qSlGCr4g0idUNTRBDlqq9uaaOCo
lsO163kwJb4RVEQeE4EtPBm/GudGLJ8izs7Wb5JJkPPqMUAUIxda2iUaOB4lKOKieNI3ZLIWblcT
NSbtF8HnOrRXfkSzEveP65RZJCpryOBdwiE+78Ddt2UhDw77R2f9RY9fSm9AwKygUPxYzUCCNuAb
KXP+S4Qh08lh/hwE+TILhrZBREN2dblp2bjYYBlv94/AO0YUmXtuzDE/5A/6zBdmb2Efs3277hq+
p6ohK+Qj4qZ+En/SuDvByPg7/Qp1FdXgW9VtBYXwu4HIFlmzXD0or9Ks75lNk31cveQ7sYgSEAll
bAikz3VaIg8EFZ0EVOSoD7qyRv3eNkGJEB9JyEEvbNEf7MfoJwmSGIwauyG9aUqnZU61WJBlK0V1
nVjP/+3GUtb/oIWkuX5YVs5kR96GhthVMg7aAdGb5kjyGc2BXB1aNuqQphzsq/b3DQzvTnbBTQsZ
bvUk0MWM4Coq5hRzyvA4oN/uoGOyi8kfd0pcjZaALtZdLfqVYinJ03pY5Xh1afIk+B1IxjjoTTu7
RiAOUy/pEfNudxh0OSEECS7EfxnJMa1Lvn4kK+w8cliOp3an3zhabJs6eves0XxWu8+6kGVTCl6C
Mewx43ni1AnNRcRG6i2DstEHk+4j/gMsQ6jRDjvf3OFYqmGOSn3K1if5soC4O4nahuJK74hLD9yr
SWRHaND35FLMreZDOPYIpEk018ad3dVMBVdERk4Zzwr63oRameVTthwUbdEVhKG2SaGb89e9xlPo
LI3j0SoqSa7jLd5WvDGJhDNcDfR9xU7RMwdAYIslQtV1kMXNF464GajOb2H5JxzcW5XmMbz1DmJD
i2c6PHxLM9GQSG4uTsfbSNSC8DkuW4EBfgtlN44LZMEKP8olE52GP17WLsDp3OrXe4y+5EMGgPSY
NpUrg9JlGyAO88i6l544inJPwkpE21UepN0O7weYTlsWbknjysxzsMHrQ5okQ6JXZoPp9XMOetjd
ejQ38giTLoq4hIm1kVc72LfPhS+7kI5WVqm6/Kvs8ryT5rGHmMJZ/uzzr67O4BDSSAI+GhzVgmYw
2Dw+KRP5Y9VkipPH1lcKATqHmKp3urjI06mCUIZ7mxHJOkABJh1DA83DuK2vmTZsfCMzIGPVX0i6
eCxVCNOzQpCJPJpnwiWUTdgSpGf5J0OlznYKzo6j2jvG+pgXkN8fD1Aidz/9ktvtH5D5hK5hqDXI
H9kyqQ5lpQgIWLU67GHvYww2AAX5IvVbrnbXYXQGvHP9LnLVzF9N3KE4BkgCnGpmN/1emG0xwhUx
LM6PmfzTudS6KKJz5JXPYm4SL7ZQ18w0iQ599ijUPqlDFwKZG4sLkWQ3PTw9D/9CHY1gKD2Fu+c3
zK/R/AjZSBlXWOAtB4Rh+luRsYx5Fl7IdnPRu745+HYjuv0rY3EcMM6yh1XIhf6iu/qHyMUhYfjj
m0PKBYWlvsJfALIvwLjYy2t/dWl0OF9Nz9Vj8sQcnXKlmmzbdziIKtrxIPsrEX6QuLpMwUjE/t5r
hvus4HxPdXQARIfcs9d4kVHlzThXB6ZgZojBhCaUjnjTK2DvyzvRQVhCtoLnPp4C5xlyiHOY2iqq
pMY9gcXceHiHOMVNoOvD4GuQa+VzwVk9SivwF7hb6jUBbEBLlvLmXDFypChtMv444O9bVgkMGW8K
HZ0AzFlSEQQDdLF6wdS4JIpI+zaVjOvERT93fy97udC2cAJAL0zgSjgH9BZCQKMlOppJQBNeL7Sc
Smpi63ALSB5I/R9MmAJXCwrEF9BSVD0doabmz1uY+wCzK2jgmceN+90Sza3AZLXYqlypT2J5+q3R
CZ7fZnWeH4pqEcIRoy3z3XE2iNzJeC2XYhJ1odjjUr0tre6qKSRuvbMPcUmIplBX29gvt77egiO5
95ZEpduTieBYbDkyqXKPqLN4yHfadT5ETjYqx/5BSztp7dPsw+R+q0qy2ZS1uiOozbUj5iDdx4aD
QTy0xArrhsZ52BmK6Q7POFNEstH/Um0nCtyEDUFKj/TdzWdWTPMnfi1F2KCI5wS2AHJESPf312ep
kHETjUU6OFjPrHX47+2Jc18jBKZxs8ataa8OTpdh4JWwAHO7BkW4hWCizsCeumCa+6l7GSbMUlDu
yf6ydhkETkwlOgGiiMqu+7gTHIZrFftY1nruq+wWuO0VEzq0Z4jSaSNyqFC5OiPjaRhXsVinltIV
Pz24V9S8q3yxV5t4O+GESp8JxMo5sbQ7oWJFS4jDgcPV7t8Z9fXNpsC349xSZfPsWb/jpJTtDpGV
AanoLK3d5aMZjv3QwEfXtldmB2YMo7+u6j+DNjUumBVT1AQEM16jhMpnVOTaW8EdhQW7BTLvjqtV
dKqAuQxnOV3FY8LlazsmZj9n88R7sHO9/VF5L9Hd6q3/FWqJv10RAN7F/IIT6q5IN9udKEKNW9i+
tCuEITdp4eHUz2Z/l6rLTY3M7CJT82YCAWStPuIIK6cGr79vNa/8iG4QGZJpz/0uI2B6uYYkdhUz
o/zNMQn/283rI/L4EW+/Fz6oVf7/Mbnk6Nb2F27D7QYm0lxTWVzqEPIkimaANSI/Laf44Vzgx498
Z3nwQQ6bc94XWXg0cM6Ov8/tLZg2vPoxo64E0jfFFc76Lm57T516VlQAbKR1KXHQlropE1g2X2YI
QCNVhLBtEurfDKrq83ILOZjaY14TA3nb2Wn28UC2hjVC1VB8Xy7sL1AT81+glvGHHm1oc3Y9mD4p
v1DnWBYehJeDHN/ZAtmi9Gs8Kz5yiRCnVOTcg+5sRkUk6VJ5zDb1morbOb43wLhQpcYeET+bBDS2
o4aipI+NngSMfQqWDA71kYJe8olswDdcREBTeAyOHADFu7qhyR+pRZzeJQIoCKw5iOapL/m7zHHU
0Un7sEFGiy5VvyRlZ/gOBEOa7PnuR2OV0iv8NO3FbzGkoPlPfQ6Vz+Oq5CbFznb1CAzDtDZhmxnF
Tunjcs6NGCuVAC1kcE6K0Jwy5P3MnEyXsdsi9NOMyLDI/XD+LYOus31XImed0g1apyRPXOfyMzg3
IGZZdlv551tmt9qFB/2vd2CENX1oa0q0dh6//aYV7YcmudLHXfiq6tf65DSsEm09GzvrRVKRigkL
nr8qtvTNvdIpfhlIg7VZmxhrBIaZUr7B8xB1UIfWcULBe80rvycTsBi/0JZovQQx2bpZdfrdToE/
kodhXCsSLfp+W0Ml6c3vd6hnNH+jOgOp7iVVA97VCgin4wRWoEZ66QmG3ynl8x1yROt2ZQMpzAJq
yhTAQyIbRMcabLDvVZXlztvrUUT9evysM0hRYXSFKtuIqBjkqarI07i00nSIHY4CPqB9hEy3NZVK
ADFe+vud+NzeP/sFydnfxKB+vyxEW5WT405L6o1XsyvyxFoEPFW+XPEfm8SGtxEagHvhT9cGnbBl
Vx+ryxM4DK5bCBHMvc43aN9vRzjZLTJkdgsd7TcYc6BYDSSYrqN9WgxcL0Ivuvu6VCr5hXeuDVfw
JDQ4sfCTRvxWYjzfoh9OcvRw4cW5l3dC/5mqYsnJVfWNoJRc2nRpLWbOVp1VdbIS80m7JQryTHbn
WJ7isC1p8SyPEcidHIIlSpd0/BQCojslH0zEDOkCnWNqzPdJxe/b6WaBEw0uPYhntrkcLyrZuliq
S/b6rbUyWoCN7wu/LMsr2KfJw8xo5a4h9HKHXhoo6u1BrKzaA7Ot/haZncFWWlCKqppTO13Lwa9t
ZWhIQnugkuwAczoMCh5BUP2cGKs4fKPhjl0QUfyC3hnegSHunUTn29CXio5gkC47oVkSAxtZjZIH
sT8tMcLu0kZSZWX8XXTRVWzDOtiwqRwIxUSfbL32P6zQ2DspFlKTy/RankSaiW+hCp2wqy+PYk7C
6PrbBuNkwopUTNGE+9CsASWPti9JxyELFyDz1Q0VWVRSnRavGF2NXR2VeqavxeZpWJtzsvuykYwI
UihA9PxBYndtWE3SGdEJjSh6M/EaKZTXbLwTTJR3rSvK8kOi7cW9TsQXzbGFVaw/+4U4rlf6xNtb
vf/fxRIX5tZqC30xy6jydvjIHnN514jDZym1Rh30+emhrZrwWTQJXw7eSUtWhPp7t3rUEmnsWgN1
G1DqhmTh8Lscnc5fZSci5n9z9m/WAwkRAmO30sxZRpxm2a8EfqFv44NBnVrI/1y62JobU+71zXzS
o9rQyymqpgUxnIHA+MUxrRVgD/v/Z19pH1FijEc6c7NYqo56XHofbKuoBNbZe59zSheVdqnIFBWR
1Fbs2d6WkOC+DMnPoKw4NMJipF/E3dv1TRd973BrKFDYj4NL6sJ53cclT4EHFlmFrG1JOHhxi9H3
+U2c/U87hOBjYbwi29585TFmc2Sw3NKg6o1q8gAaxfvoEjwHptyw+KCqFu5k4yr1YBnwMR2pqRr/
Kj8WA35x5foRhiWP+UhELQmGqrwuFidhrmcj82E/FHBr3oyNJTpyI9bnKyVPYKWiv9ilYD2+6p6J
OI/xmN9p007U6fA/2OrOxU6YbAlcjQVOR9Zj1IUkd5fubKqy/mR1S/UxfMibl7pZogypjC+PA3yl
0gfcKNTsYOHqcJPOcPQj33g4wFpXztyxliKY3+Hwb7hmRKLjaLGafydYu3jiXnZ8BO+oViCh03/x
lJ53kHoDnBmQIJ2NJjzvJH8s2V69lGKrS40VnR3BC21Sw6oXei9ciniVlVneonMQtyaV6pA7Dgc6
sidx6AnXDIx9I998mMHIhBZuC6fTkSRokFKaPB7ad6U0xcwyC4AF9sD7bYWlUc8+C4kVvZpcjhDo
rqdS6Uwi36eRWI4m+dbtqPj9NG0KYvAg2v9MGkcT/ZNlUJkphgBWegz2ou7F85LmDWmFkBDpUtyv
RLz4/QvS9UOsPGEA08vMzn5+lh6GZACwS7NY2W5f/vw0KhQfHebL7m3u/DgPFf/BuCBoEraINnb+
/6Qo2pXiVdUtG89MgTWSEyQAG7bbLOQoqKYIzCFVWGR4h2303+KbwgDBzRLuav0V0AsIcgKQ4KbK
1zU0pL7jVvOvEcn2qtnNbTOhSSSgJz+uKRQle2SyRqX85INeAXgmTJ/IVHwb5HDCZe/115tXbVFl
cEyDxIuz0Cio38DPgkg2fkHs9Bjjn3JMGJSdptBEMI+adb6886kBtqNciSeND94pipBgMKGUP+Sb
AddUkkUtkut47kVbxC6RdJ0sxFEJ/jXPxeDVpxAUttuAiCB6vLryen1uhFt+VT2With6aGm1dPgO
hOiyBbudKopOFcBZ//oxV4C76VmmjsSPz3gm8pxalHeIl5G66YNiUyEmOrIALUQfOehwDlqF8owM
gN/Evmkt4xom0S2FV2gminLCiOdaXpfzIWlYlMVWNMrJTyEhRSFYSl4G8Sa/hxkKg+MRrOdkibA1
wW5UjuYDPNE4rpvhliFCdUPEP2t0pZ6XzTAwDuaQszGATJVeKhPpz8p668YGoxvwXLgDxFC5XvBd
bs6MEfCkoP+8aSckzqYgC4Zg4qqCljcx2cKMxjMRBl9mWHVZ9G8uUbcTB9QoI1C+FPvTkFBVwiCX
OPzpNag9RsyF3qFIggVygTwRn+ev7j/48agVawvCemuuCKF3Cqdb33t3WalcmU3L4ceUwygrPcyX
uIU43turqw7v51qsC96CMrXhrsOZq3l87qgbEaDWpxk6GB+pFHPoRZOAoquD7idoO+RzzYRfF2qY
PbLJ05TOMmAgW0OO8pHNg6mwju5Vc6+pHWBrNlPE5zyuSUjwPrGdTdUW8wJABm7KC6Jh7TZWfQ1S
zl1s2nsPIDMHuZy7LBr4i919I4EGDeXUkp1A7lybLLBKPoGYYZKjjeFXthK3pplh8+a5H2djWy/r
4VBXej3/k9j12JfCb3z4OIlVRk9u1Ieu+UQAPWrAyvVI1B+yuFv2eqfUD2QIbFg7Sugt2hJNqm7O
SNm7+GUhr4zTvCam7vjZHD0gUYOxSnUiirJQrA2B+cbFUMjZObY7hAL45jGnnjbKi/fhkEg5Jz/d
UU4ZSL4++903lkgrhuFk1ONfoodd9RJqvl2BcQXlLt1EtCFxZiQK9rp3n57n4DCe+YMdi8zEe/9z
l4QpzmkZCvOLIXPMSWgRqKWqClMQan/S6f98cp2P1ex29UkNzULqKRLGutZEhcIOO3nfrkVgoXKd
5oAWGPITd3LB/jC5ZnSDx5e1PtxXYI7Yt+sxhzRj8OxFKOFWNQ+CWa9xvpgYdYK1WToWQL7Xhk5m
Ozp9ZgdTwb+sm2WN/t32ZLRUwoBoj8oLzsEGoG2O94XDJWeonqVUSC6YKkVeZC11Tjfq0omFD3ZE
IlGZccCJOBLQ+waLwMmk1iJbSry9My8evfrNLZUhsA+SB6NMHrjscxckZxTE2LV0dK/EyORvTQ5P
jrw2ydqKfkkLHVut5xzSp+QQLylVjMAL2Vu4tFtjV3q6YBE9ugWcC8EPpycR84xdCM4wXJsDMo9M
KS1Xrgax7sKlU4yOMa+Hy7P3a+7oDKHcaOdL3sKTIep+vnG6aLPI4CajQfww0d9UnlGCLuo0dPXB
EYGUqEDUqvby3VtOsIjSQC/GjZpQYIRcTGCBzTzN68my/HTFWYElacduvsuOMANkFd1dbk4hBUD/
h5/WDMApT0p0mjptuZN7LPabQlwRY0uwlDD15oajfAEIxjL8joMYv80WLZ6+/8y7a69vQ08y4G+j
4oU0VVyumSKKUdyKeVZeyIQ2ikWNOZ27+L58iYgzplGZLT7g4Rfe9S0295uZM5g7PF2dj5OGOiE0
V8n5JPuoD+ryqL+sRFLfrOEozbjEt2K17gqhKiSNjB4SbfnhWrDLIIfWaP4E9SZ1eFOcw0H0c46a
kP1Vt499KjVuHYWmg5I3GGnP1UZAZ8ft3we2xBI7wIquYVXMwcI/nqXIu6e9ThaB0QSP9/7yjkwT
iF8FD9VcfdPhR+K7jCKtrdr8p8wF9S4t6RpZco/AVr8k0D+MhaRWmCmFj6/nwTd8+ROFuyULsT6Z
dpRbIWibfso3bQjh2c5pPFf50zeWySIL0sovcdD7ONo2AYD92snhLKlKwVh3WOIs61YY2GF/pv5r
moo8WVzZlra5loY0pX6pI/91XCfPFQxTLTx1aJvR8PEZ+b5omsU2ye4IOhhGBhi5LCPA1wwx0sGA
pXvrqDH7hqPj7ETFJ5wqJ8rGUK4Sd5TCcBGUaJSa+LJ93F4h92M1Ycel+sCEb/cchCfet+1JraGN
NnyXmz4visOD/fka66GEmUtEq+RYD7a3zCLKxANM7OsVa2wMBGGir3+okuB1hi5XGbL8wOWbFVz9
ZxFVX9JQamxJ7qiVYis+CE1/orIbgPgYRHZwNyiGRkUpGKQf76Gf3iAlGLhnoP1st2RybGU1aVk0
FwcO/Rq8wTc5kZyAhRprufMJPr9dJ5SC6yUI22VHFUY6S6zL5oJvgbffcjc6peofguGnwzKk2NFA
Ka1nKKHUvFrkbnt7fo+g/oTYDKWkptU9LSKsheEGz4pC1Zuun5EpXVXWVG+A6JeYFfveFZdeBJOw
CXf/Ndn0US+lrwP5J1vv2VZg/H0mxxbLRFC2QwFg9K5IesEpB4kQU5wt9GJ8p7Q8ZwdIHURnSw9q
uPN/u6/yQGswAYMiVWQB5MjyQWaGwTiTUpBNIKFRXHk+MrMHq6nHEuOxU5ILTqnpySc+RFR0B3FV
qoI0kgb1s+4GNapUx7RHJjrHl7sDE0XWfn6nrbdqqe/dt1b3iObYfzwFbnAy7f6c6yh/ZQ6B84Yw
sF3qbTrPaxt/dEfo6biBE8twZwP9KBPXb10RU5ekwp80ZU+aaxMNl/ScIcxjfSVp3vDJkBvr3dgC
QwvR/REVefWA7evbRvhvpgmasVLq1MXSxZg3F27wJlzL1MzcwLs9aTkSPuezEJenlOr1c6vQ7MXw
W7lhkP8BTexv63BeomB+WvWS++Tp94AAE5F45Ut9lJ5eDk7FXIBKz5csJkEGNukzYlNgWyMOMKDF
MmfBU5Iq9PmYH7NTPf87g1iagz5ulPQyPw8dmsofM+SSIXZOAYj7GnwR4SlhH+ybKB8034oJ+rD6
oLFTlVdtW8l/ySa0Ej0Bd2YMYG4k3yTDD3c5wgBMlxaOLWokSWrC/yPG0RiCvwXxX4dLeHSznCPe
t39Bj0vXeMAXI5YMFJh9lJOJ5MjF3hgHA4MpvggWldtkj+2G7rzzQ1u7s0QWOUBMiPN5U9sKjxHj
UXE5xU5U/HB/nmvafuWCVvlirO2N6x1+ISQ3aPcd8LYjVXp3HxR3Qii6I5Ac8nFrRucwn3grLFwf
VvviqYiIEqx47j8aEMcWhSnXXGmA47EAIPQuFFJeLvyWoN3mFl25dH5hnWywMrA4ndZ02SJbZUJy
BZCoMg54ye6U08TQuvFUwDxdvVKKwgwsXrecMJUv3/VgccPGKJKa2YQT9RuSPFW5iQccbMQmthHY
OJrnC2HUL4psfWkMHiNmf764Bc8T75zzDe5Us3hEnjj91jrNVA2gVb29/HrhLll+hXselhcOjEdD
bmIahyGDEd97HbuvVDPs2lCknIpKzh4lnPlfcgprM9A/p4QvaHXn4JqeUu8iBigZ7q/RrHpDTaIm
d5UTosXhMKRvciW1wiEd8r2uagEY2ul/1kXhxwQxC5yZls9mkAKpf7UNVsCZZl9WnCQJs68Xv3PP
8uYg3XGoxIMDMyif35JGSIrmA7IjzbRxbR3d/7Rle7+qAahO+1IzujfTx0nBW5C1ZrncvcK63cvB
LyVZWkeB9guWl2uh/MscKsruzjYWm2wu7qQelzp0UY80gMgyUX7qgoLH+rXz/NuZrR4+a83XO/QH
vlIEW6cmo6PznteMc9LOi4JZkM+1kaBh1zfi+y/VEm/V3dG4xms3v3C4yueFJCQSG4CPke6W7QFA
AFlABmKMi+F+5xsCc1wBApK1P93pfwwZ6zoIcjo0Q+7a9f2wM44/pEE5Saz6qxGfT/co5Qxzd+XT
BPt8e214rSgAspmwQAGJ4jdkgl+XWNvOKa2tgniTixMfmMoJv/EEJbPKfmQWAYSCdZKMISNmVzQo
zaYtjWZOBPaan+6s+/gLa7Uhfxqg/R1L1B7MgOBBdGN/A+lj44Jt1Okb9u1TqQwea/3IgkBEAla6
30dzxPL9WcoG/JUloCeeOkA5cGCqzhgZTOp/l3F0WSOhEqIXnh3q08Nw5+KaC5aEbNR2A+isJYgt
nRXT0tDfbl60FV/v4kXz8Z7jQGhDHl/b1Z7EeI5xIvP3i+Bf6RRUFP9CPVqid5NBnAVDa3GfhmdO
deG8SmQuZexXRDlAOTuKybbFhoFVIcJ/xm9JOf71cy+jIxo1gRwlj+OlS39r8WndjF3kOrUqpxsN
Ck9gLLdDg33JSO6h7qHMXt/wV4QSNka0yig7YLxivSfKCfO3r9x4u3y7R/tHTTpx4MoNlADPE4Gw
jVHkGEnNSEiFxMHqZLKxOXWJJwPCeCbRHqpHJRorPznxA7CpmsxGCKYqChpNXFg10oM1qDJChyYo
DklyIy8Si1ooLMd4gnoYPHh+H5Z1bCMC1+m6G5Rn1TjKo+HJMJ9FYaPvPTCqc7RONPIz6TGpgDt/
A3ilZTu6oo/k7g6DwX05UxE/aqtcxZqv/Di5xznA1cKtM/IquOm4798C7wRJkzTGb/HzuyrPn9y/
R9sX0BEO5XTe5isrNLTK/RZugaX8U6kGGOUt4UjGRVedldO+q+5A56CxUPcTgJFxnTtir/D3BDqS
jFpHem8RyB9pDz/Nf2G2t93xucCLqlczzA0unwHZbZmEwJdoL+kHFleeQB5bsDY2+P4rcDlcqhce
ozpDbStty5pHPseAyP6/sIbGAQSiOOZ17ojLis5M9frj+5/FrFBOYHCkrd4ith31E9QzYTqo2yLy
RzA5MlffWfHtqc9lQg6TBDmiwrmaP0swljwwccUCGl5Hsyz6OU9+07fcVRnoaHpcHbF5feb8NZxP
3oYPRqjGW765IkZyjuXVUeyyvadmQEXGZOW5t7JUSilMIu8aWuLyeTvRzUvEJdrzinrqIj0cQaCo
rSKW95dL+kRgZY+bSebykNL+L/vLKNaJUK7YyQHY8wH5j6Qz7Zih14D4LrJqCTdaaYU1YSgT76r9
Vtt2N+ScWrTHw2qxTZtaPwn5b4QTeT6jikMRkDiSbtOipTrdanRMAeNmCMlj5j7VfjJehv4hBFmK
7XS8+DdBZUsSyD3bDria8OCYiAn5UXOZ+1jeqWypMw2IY0nbeV0ZJh6RgXb88Ua3Om3N1Amw1CJA
ciTyPHSiVFf81xlJpZtHrB2OyNv8odO1AihRTbiy0Gn+4H6BIasGzCicl57NXGFysuvdypJmt/SL
89PgbGi0ODC6Fz4+2+OGnqGKe5A2rDsrKJAFeyYTLR7Xv6Q3+uWbYnjhqw9modunsAP1X1SYCtK0
3aLeRSHppoU8Bxo1cHLJmYhnGQM8muP9oQQl2gJRMzYxc0xYjqW+WUqbwMUdCfZfx6LRxeZkjHbv
VL0WRxfnInZDGL+42LnGSF5wqRbTbqfyZwG03+UM0Y3FHl1y2oIK9mcIn7aFd6K1/MyBKZ7Iy1Qp
Ni4kDBk0OF5Hofu0Od1qAYtEgahxW7e9CdP5iVhAmX76yB3iOFH60qOzzWHUeeqGOvAT6asR4hgY
7P4W4aKCzRoLnk8pmLF5xa2c4A9VA0hASp4iJMNhEmRmC4SB5nmS7bZLCQL1NSGq/LFkgAYtwy/R
+pVvTmdobq1QZyMEEdtxTcJzBryQ2SYfsXLdRdNmsyo1yfnH9cdV5eHK6fBt8b5aM3e5xkDcMvQd
NLbed876JF+yTmlAGz7GSj87dsnxG7DVwSdPy2SFjLY74nAne8BPGxckivJfq5BOEJ9LDOqZmbjg
mORvKMSLRei7SOOmHRsMQ0yXG76ghk4kndouMRY7UFg6aox2YPy1AbzrdZoGV4lwnJCmCo161Dq9
j0Cv2yN0/Yz4IhRe+ggqlzKNBNjlv1HWE2SGpkhL/f9jUghp4rwg0nxe0LyUbL/flFY4Ns6I+Bwi
CoFRv1Qw46LDLkrR91aTZyLrMiR+EAm6vs/xIE3cQGAsVwC7Y54fkfTKlzjbGpt8qvlKwaJQuNUn
/JOxcBqwxnZotlzW8EYy+4RTeNL1H3ONWUkUGHE75mJb8o8mcFwMNk3Es1tVkVwqmrKhhcfJQUyo
pQJ8jILPR5W7ea6NSd9QDp56aoiq3J2krOuFKyiC438ciCfV+gbP2OQmuMJokhoIt5Rpvm+FYMPN
PyjkJ5L9g/WtqCnFCdLKl8T1cVJKpBY7nlFNllgoD1qcyY31uqzGgqJGUCQYQnjlp0hDE/YN2+2q
5aq49VfZWXcsYlw5yewoM7cbtiwXpnkumz2eFqp2yyvCcolGog2lWGh/BQrN1DfPikjLxtGOzrhE
+mT13a9hiXesCpRV5ukLzA41UgK9HQorG3PNN28XNY+ngaSP6cvNYgkJdd58ogwy/0V3lR/9Hmly
+f4ek2bG6LwL+24CXYLkEiTTzMUIm1Gn4ZbSRpVsKa91YAH13a9go88aRycA3KOUiTIDmCVBt+OU
wYVVr+ByNOJLdY51wSJKmHA8lB1J5xAIVsIUkfip/3Ii/olw4HhkJYZNJRQhYO8VnejnMQEX6RoD
dwa22PdlIwaUQjhVfldDxK95kprzT3elxuiOzNviyCjXVDP7yI8CMRJ5ezltGONLp0tKAAA2jh9O
gSisiwdza9CBPPSHiP/Hq13NPhtdTL8pfuN4NObb32D4bhNHtORe7+eBIQ+13fVqCq8asAKCmZwg
2EBw59M7O9pqqOxrGmyNG0P9P8O27bZFZgvKo8723eaTro8RK98mVu8TV+JqNwcfeh2cgAwBZr9y
qNhz5ZtFPmS8YEsYWJSjDSwK53IvFPfXFlP9su/wmaaqRZHseIvaW6FwsVZZRU5/fjE9AHdKDWKJ
1ObHYco3Zf6VAkgQH2NkV93B8/NB2q2AWFJ/T/HJycemtKecrisKVRpXbo2vrMm0/5nIYt0c7eYJ
sSd+3asEyd5CCDXrdWrg0aRxOz35CPS/Z3SLcI0qtpvCBpimGZd7/wB5+J6vpRbLMFfRD/XroNDJ
WJ29e2Cq/kc2G3uWCfS3NKfFhjPC2tHw4Xp2mGWOEsUhxC6Co6QHoL9K6N5b/jZNE/bY06xZeYM+
nzD4kOIe42qXvEZ27zR9uMNAhQhYR5H6Xdm8HQXA+vkmv0Afwhav7q+a1Ev54a5AdYJlBO6f/vX0
dkKzcL0dQjDPY1mG548mP6cX4jx/CZ+s28K0aDG0CjEa8vXI9TS+734pUXh2EZh7B8b3NLSaot1N
gepagR8F7FPpgqVzSV2ZtHG56m77W1IGIKzt8WbPvYNegE4Z3Tr8/06U+7f2TtAEmhr8DVLzPWE8
+GLg16O0Ot7Op3ZU/z9B5Jh/MVRS1zc/20H8/cDJeYxhYuMC1b0rA4rkWQcCvQcSFgkOOk2DXiEd
M7FNdmhNW6efrcchLSFjpKY+XFOZdedHbrHdKJrUC9YgIHDM96THizCA0NiodGl7na6JQYaAgW+H
PR5FsLlbpqvec+mU3rCLFi1ZqA+txkakOm7L6tax3nHnbJyFcnKN3UBaFqm1EZKrOCFvlTnf1Qx4
NjivM7uFv73XM7PbVLYdM2Kud8yMJEIXQ/qCAwjGAFb/N5GsdIXaQgY5UAVGtPXu7jJyicy9Jotq
JEwdlAPy9sWy7SuvaBIBxo34/P0M6IObD1pQNb4/HzEpEaFgsm3rpdQWKeSGFZnWf3P+yDldOzqZ
YeoHKZHU3VKHNqZGmWK/GrhvvuAneeRowooPeN+EVt6VklX80wTqEoUKt4xBNBW6JBoLmOP1bUak
TdQTxkBoiBikjdiQA9U4UYF6/VB0TU2hCaktn+8nt91xK2KsEdMNcVutb8PwuNUEWXMiAlX8Vlik
g+jOingrzfK5jAHuRdWDUQbl0mkbOjcgVVzlGo0f8GgGTfmcV2NknPMKHl+/FZYQsJipqdrRoouc
UN5YhJFanTSxn3d/MNeAC87N7HDPFcn3lWRjwXGQ1p1LhIBTmzr3XDNCrqm22d3Dp2Q3G/NB0nFp
a54wMBb74AOfg3sUiKDwUa8fiGX9T4ff1qRnG/e1y0/AM7KBGvAilabwJdwOkARMi3WN23S4Rso9
Zp8H6ecAq/eEotH9Doo4CpVpQwfgZdz8ogQngLRUaSjFufbJmPTKFZ/GNwG2ktAvDYJS2k//bYeP
Gh13EXBccP/949prprNZjhZQXTuyIE6osiywL5jhDx8JuMmB9xKYE6EYkn0PW1esO0pkbOCmrSHx
nan4HV4ha88cjUxCpUYSfvYM1l1cdnZHNHg+VeKg4EAbukzkzfSoEQ46rFv1UEqtUe75NIKiaBgY
1182VRPnXtKFHyu1D5Evkq2U1QYGamnFDvPY3eTkfHaIMrMDw4a0vsGNTJxmzMs9PuqvzX1vK5bO
Tl0LcTyOTamNZ8HJJvcd0y7v5vd/oJciaJ2FHlPprp9WVE3RyrfdGMoCRzwAYtZvzX2+z8hzmluQ
5ca+WJ3/zDRm+f0hHUbUZa+7pP4b2mSL/a6epzkmwO09hFYoVkF3QmfyuOwYdbN/4f+S1LndIQ99
F4y3eJ4pW+/C8CQq1n3yp3UTgST7+zG2i1z+mZNj11z0U+D21sUTpGGMPenwrC018gIoWpNQ4GSP
wJTvJp/cOM+eBFR/23SA5+f/Gv/P69Fo0fjsgTywO4XSG2fJIdsydIvf+al+mngndtcog3QLxZ6Q
cCqrv89hRltlQprs1U2cRYjLXmTLxR87NvQVRrOf4ZwtpTE2dNHMm9WtjPKnJVnQI5CDTkLgiyfW
IdEWuADYUy5uNSsKQNJ8tc2gS9FKjef+QbP8Y2czlCuHtUBrCy7iM1opIrzTDS8RUoz2wMUPX5X0
LoUmnjRn+rOITVwayeoFriZGSxCT4arwQv0oxzJneOfQvM4s7+bGM3YxbAsgH6YfeERNW0dApmVd
3Nm073qUCWFieidXVEQYmYz6RsJyCxiSCV3Lcs5mhp2h7dp2LlDDVqc168p0Jj5l9SA/HYjW+lJj
Wr4JWWrhxGYv+XzMhh8uo0mQIUV3MqGix4kZfvOUfXO1oeMSqRVr3t7/I1Kggoq1ab5r62JNFeiA
8Bu3vobotXUnJOXo30KFB5TZEe+A9X91k4xAxnGqEUsE+F4BlM/j/SAswMmSoCNquX5WNMODMgwv
wfS5yvsdHN2k00KJ7z8R54sztTrSzXPQgOv8lTmE9LrSKTSzOU75JAqjjFfcKjkdjnncr5OPLHHz
V/n/PGO1WRodRCH4KuHvT0uKQp7Jlh/WLFOXCCx7MYNohuZwygFqoZmuOEH8ILV61BoP6YJ1rWX8
DRjbQ9xKtXk592fyifnyaidxCdDcw1yLtQBvZdls3qJ2yb4oPqiVengBjHQ9JPUOpkTDYETL0jlL
6980aVUuwV3lgKbQCamN6WEMh8ANAT980QmA0N+um7dUWsemzRpIzDeuIQxtX9aRUx/6z4Y9C+eT
uR3yr7ntEoyClREebJHw5RSv52oXDCDqjASQgHKkVarVa3HePOru7HIThJuzLJmvas7izRzSoDBk
q7pC7fUsAk7/U164Dis4hSu2mrYWdAK756YffsiHBVryx2szdrzQg0qGIjC/xDuj1uzX/CpVp63s
p4+u9ZH5x6hmcI2KIrsgCdCQJaQjHbEoagCdvrVLB1WYuqp4jKVnZ4kaqld8rmhMYEa+UzX7CF0y
dupjdv33F9tlF2smTY8Gs+pfhedGv2QD5zRQPAHa2RAfaL9xb6TWvXGfYd/5P2M2kJ1FlBQiV2Lq
fWk40QOPYK9z19goU3HImVesaLINDvlTcoWTRrwdZ97hojhFVEzVXg8VvDxUHcUnGCHp4w3xWuWz
k8XRk+dH1WYpzXUuvkDlsIoYt0t7NaOuAlDgVgjflqrfH7C4DkXLkSn9VS2nryGqifp+lkf+GK0j
m+U8UtzedkXevW6biuNtS9e1/mHbeGhfeFC7f/b7+IN1ZBZYaz/YY8HyUSTpcjm9AvCFMTLsojrg
duUXaIMuotPV3SUVCKdcEHFdTYXZgu6RG1pRihhVlfBH6QrS2vrYb2SRvlCqzMna6NAMmSE8INYW
tykVoqPRcp827hDX7q2zVAuGrt7G5WmzVThoykqULaIIK5U0C3p4YsoBMRCFX6qSSI7o1IT1LoHd
aEVaspZLy9ekQ+0P88VyvE8RTj8MM9XM7vD7YNDS3QJHwdZapYgi5t1dyLW/lzMw2uyYgiZdwER2
rkAJQcc43ytmtJRvBXMGGMkf3C7AJBgQLZSWGtun9508BzWimrVK4Il7akIY2GfFZtoDCM+++Rn1
d/6rOAf6dl/MsqmIU+lKcnMwmBh9C2zVzoGy9/Ce5VSL8gSnfc6FiEeBYnr8izcqHu0/eP/ScVcL
/NqRRHSdfQmCcec49M1SwlA7mJKVNLYI3MeiEZLGuS1cUh28NN/9sABIywclXRgLvXUv773cWWXG
RuoqsAA2dHOselvsIF3HIPsQFtvTV0BD8mQVfAaAc8M0r9O7SwYnAn+k8U/cEvIhkmJIveSsAa4B
+sVxD9WJhqB1dCdHZssU/e9zexpmiNvtFw+aRBxAIfCEmsV41dudgvoMWLNqSzD+/7GQWPgLp/+v
n2/Q30FRI86IRaQifE813OPGeUpI9Bu6LVKcR0/gDLpdwqldwmgd/gQz71UabO1utwA/n/yEtzg9
mY+LGQt+/Sj/jt/BYlUPHREkDk3yilhVVuDJEV3hWpTGIbiZCo4oyIAtGD5k6/OnZyYE7lEmM79l
TN7cWpT5Qh9L/jsMkDIsqCPn7aZA7IXBtv1TAaLhipBmj+Hdaefclpns2FpaEviDJ+SjRiRrVmu/
SUHlvjFiXT0yeVdubAprrLM8DLjmHdzLuGcAARmDfrI+d42kPvJtEOheD8I2bganLi0mJVvNXHBY
BfEybMWvjPsF9yRwfJGmm0COwS+Go92DIlX9C/UhHyMQzXlKythLMgw0DBpNWUpfWWSow6foWRqB
7MntU7O5crr4X5ygPgnNdMDl3kr3IUEwEZNlGS7kGjMQRck7c39PwfOHwepQvGsML8dSmx3Z7Rik
6GA7bu9RnzUPIFhxR8NsOPp6Pf2raKz+gitx7ub5MQrbQS313SH9qwobdr0uDx6cK5ENFNy8QihN
v2ZWIsQK+PdbcHVjHyuPJS5AfdnS+NL/7XXUv5UIzB039Gc9sAO9xCmRMRrP+7aVoTj3bNz+/VHu
VZ08jELL8egtbpCXti6/LhpvKZP8PYVISTHVxgnMfyqyqYn0E7ZG1bl+FizYZZnMMKu5WX629LD5
oR+9aEqCTvOL4Zgkz6Q5+ldXFh/Bh4fMxb82BjS1SEtiw80WXG1BL6wsSri3TorXTnjPcrM4Qi4W
6qpbkFA7yVO55lpvbqABcbWxIv48W33H6lUG8PxCosKcVaQ2Bsr9qASZjsZGbhS6yCb6DiyVts/h
3LQErW52HTarHtOOuYm324iZSd3/sh0GZEB7ULql6tdJpkEMfSO5ly1ShzS6bVjOeb2It80Xpud6
SK9S2s76cKgW3FQKi/dJLWWBPZcfIusll1R5KQEy9JRyi72sZE6XrKNkG3v/HB+h+mZivh2pp8Bq
hJQ6A8YyrcyLIPhXI3+cvtzubpnwvGOIvkrMHjYJwTvNytwBaJ1bb6ornpOOB2ZZ/RGq6PKAly6G
RrtwGUKuaBFsTson49o07nAjDLaoaiak+EEQmA56s0bt9D6b+y6AUFKxOIkl9LrQ5/WEz0TSHpau
Cpyxue8DTq7xjhqo2FQ267X2Xo5NOIPZeL2GkJXyHLhCHHVnTT9jFAwTcsUNHpemY8N8QTa6eoDd
UDbPPIktL7iEjz9jnV7i/oAkwm05saD2OVqdpGiCx8n8tJKNwYi7iklXZke+VO/fO8bxZ06S/Hhx
Qw2EQY83jFWw08h9P7s12asZ0Qyn0elaNd+7UnyDLzhvinX8UVs2Y7DX8QdV72w6lPnQJTR5CZJC
zKTMbIA3iX5qkoIq/Wdgxs1f4UIuXngSetzWS//CLalCnFXMw0RKTbXqykSlu3sCdklY1rBt7Mfn
pHaLa/LWw62tvoUuOxHlF9Oi+CaVF90/NqXVqG6wjwhdG5AsjPyMNMEzbdO6YFBwOmfsvmb79QZ1
bXeVUZtEIL/r0poWUHMcTVNJgfw5d7PInxcrkPuO8n79JU4WVLbcRoN8DgKnDksCg60V91htSli+
/RLFAqwmrBO7gJpUCdcmum59UAqbxubjXRvVreZAYV02+v+q1E1ojgaoV8TzqFDwYL2ypxAv0HbK
r+ztbBMuCfpxwJTrYglkviz/4BNQq8FqE+oke3KUrdiKhfcpu0SH9D3MN7Xefw9CWTlrIQ7wV80K
Oos6Cj8FkwFaTKfyGeVCP651e74rNStjuKnUPbPkDNfWziPGVm3/1onOuqMcgtRPoJtfA+Y7vxs4
XBvH15yL8IQn8kDZi+sIIrxpzn/t5CMFUn9+cws/M8mq3Zy63e5SR5eOZTxO/ge2inBD+bNqLY+C
zbj/W9TSSx9OKFpuMmuq0UyZ4Gd4bqW6w4UtB5j564Q4/M6JwLxowPQezhFqc3/bXkyB8UBLMn6s
JimdYIohmcv7FhnLqIyyv+Dp4WBAz8OPyAYY6IXRGf4RF/csUPanMAGzL/q/Rcq5HmUOAlgumwdU
RWEyRCXR0m7lwrpCq0EjCV00mI2mrYIvlNOX5IinCwsVT90DyHHneGLa+aWu+h5PYSjoCSG/PKMJ
i0pu+kihw1/+P/XYAdewL9M8aQKs14f4PcTWSGuFtgOEIHPzak34pd56ayQ8yb8qSfw1yA104LPB
VcGsTm+VNds68+R1Pz2BYS+bj5D8VOfbqN7SXXM9eMgPbP6PA2eP4MwWb1SU9+II3NsJJiUSmdB8
l/0pwvSqcZpFd3nK+9pg+NJ9TTA7Fl002+wUD4oKDrbOLyoKkezMjcekpoXv2XfinCpNvgYVAIdz
aqTjISjpTSJ6g6H/yeKRZqaajeLhalVte5AtXivWlTs3XLn9S0YmbLw0S6pH+Mb3shCXH+aBDCAr
u9JRpxRTUjXnWQ3rAZiz/0UrBBrssWf6XETdlmPfjnN5Q9oXchr3UiuqIKUC7uya8WkuprBtcNSV
hbieITcuL4wK+v1+GQSYCvanQoyTwPrIDdIP5ewUORSjRewAN+Kq9qu9XjMo+SkAJvw6hM2TQbfu
OiKiOLG05EiuRbYqJC3/kfsmPJ+7bvo3zfYJ2a70y/HpjceVJ/ngeTUy3Y1TV9+8h5WSRk+bBx4e
0eRzomIx23mF/47m7HKPE9i/afG030EPQzjsLSfDovZLceTGfGTJ16rAGadAZzfL5W+GoB5sjI3X
K+qwwYO50tW6xAHh0YswQp8qbAdppT2fItxPITV341VnbjA4xeZbPe1Be61if6oUnI/wZwNXm9XY
Ckmw0cVII2VqCdTb+awu57Hd41Pt++k7rsw4pohT4H1BSKos08LKgAFELP0QrJiT/b1HFGHbIEaI
x+37NInIUbGSFc3QrW0bL5P8/273sAfSEdHV4eWT1QwqmxixYX2p8zFzrUy3Ak0k5b4uQrBffP+x
AiG7SM81HteTzUKlGyh9yCCEYUCdoZEpaVUd0VdLj6AVfpHpvNpjgSnJt4Eqs6Wi5DxlX61/2OUh
5O0vmSzo74G3U+5umPkIU6Oe8fETODdfJf/JJPHmu3WMDtOc/20Nkr7gT4lmzgONvgSBsjIVFAJj
whRGIlEZztbWbpBHdDgR7u8zLPAJI+f+MjOfvu7+kXHKhxme4DkhLpyioRcYrzeufdXN3/OAbOI4
+lTnReKMz9uZ+zauyS+cg7buSF9Mmaxap14I2c3mWDSxWoggqF1vi232fT14g49hTNR687jY1W8i
oln2Q8OIgNbeaxxxmq9R4NKmGXAOO87lH4GTxn4Uu4A7E41uSwdB4J0MbFkVm1sd8F80SbYjU2YK
lJD67hlW50hHZcQOvq8Y5JiIJ33P39se7rJ1uJ/733AD8PGZ59flLGuG9rbpVPBPKTZeTodqj9+o
7vvyKunucJiE1VbM6gnYTIH3dnGpwQ8MqwavNO8kFgLab9G6bq2lNTKqpxb39/Ss6JD7HBg8PxQD
aq9cn3epWAYHafFUCFI1xb6CX5EQuaitLg5cJ993L4VikKIWQkmJn3MZDjzQLOUJRRY3WhAhoRDU
AzugEfzX3zSHpIpcbsa2a04J2lIPP5SoMMV6TwrzEmBRQto847YfDIea6tPaZvm+L7wqUqdhqIis
dn4v8APgel/phqF9fM7dDE15Vh66Wa/DvMvQPAcHKtyi8I63L/ZjhKUT11gYAWVOAHa/HZIEslx+
u4IvPxFZDZUNlrP1r7AuHW71xaSKaaEOvAr7ycLxG4YdZ0JGp2cO9884QUoptzS1/HmoC1VJuTOj
/WZUPn2q//1CCegdRIjblLhLrxQ8gGUZGeYc5slT1OJw4ozpAPvoM6fEONr7RHPTUhv5k19DOQ8O
tUHHhsjn6I8Qo0dZr/BxmjyCGJOqpjnfPoguD+GZu9MQwVI0qmX4Ns8m57pMlpSEG3IYcg64dqE4
fB64Nk0GqxMwlZF3XyQyZ9pKifI+EPmfVtHzCPLLvLzfwXCAKmpubt4O+dkMYOEi0aE8MoGJB6wP
OB6IJMLaUk8kv0sFwzDtlkmYynNitrPjxdXGgnbTIYA5yTzYUZ0S1NvWMaZCiuTZOsOwLn+oMt8y
tbciR1ZzWhEuwyC/ZOlW92uXH42rLyu8t/UOsXK0Hh6544TLFkq4Q6pzmPuOew1Fh+LtpDTeBqQj
px/g25lwt48WyPRJ3CaQXcPrnHD5bzV77apr0cJI20eX+xt/DiPNg7BRFHBTwplmeJY6asIpksOw
CqJpkU3n+qcioVes/3INb4rgFtpFpGZAjJCTHeY2mde6s8doD2SDFCJk3UPpdzI0gKBud2PQpKER
MjwR84bOqK5+S/8CbwJYF7n4++rgbREpJ7yYD4/uh7u8/N5NwULaKb/TSQDlOwncx0diHjL+L9OV
GlUQoQ1kbDcvFD1CO9/h2iAZOH937/oq2sQtPmdfuYjmgtA7YQeydQhgnfKU+cVpCwMVT3FJVxwD
tNXjadAa4p9f1vFNfaephclUPol0Mo5qD3XpGvc8lYeqh4M1TYqEcBQuE7uyF7bZxkCLO/3in/JT
lfQCIupRnF0B/aSxsaaVy3u+Ww4OQtWpVfzdAB+RJz/W+Af/5sbOQTUfWVg1sL3f4CazzJm9wVhG
fYcmBzhrEethg0OxhFSvw2p7BEUBGPjffV8H9rcZkewuk7DqHetsJNAO9+mPe1o2VidgrFwo6Qge
TkuQGpJqBckvFYpKfPgBama1rULqBczYpFVPHuLh0nBCByPEKAVGygx4ec4KhawVl0YSOnI/EQiU
EQoamkS3hyYBGfwoBTasA3P0YNlNY15ELDxNwB+GW3uLMc7OvRyoI5pHlLQbwRc7wmiJCP68ptcI
8EnsbfjebeYw/msaK22Vavqc3onNr1tXLe7WFfxKAC9nZP7gpxI1EcyumWGddQ3uLW52o07By1qi
G4ZouAOFLMylLjQ0WkFR0t3OewNfrLISfP4Wt+9IDt+/WB8Exb1NKWmrU7tanRxDuqdS3DMeWf79
WDlb27dT23Dsb+XwHI5Ah5oqUf7ZUbdob77dYjJwL0+IKDrml97mKjxrD1tGQs8O5aBNnNoMzfZ4
Z7x/A5hxo3TjlqmN1Hc/xbc8Li7oDyHOJ0gJWLjZ04U1XFKzpa010OXvyrnIliA/kgXLsFKr7KuN
4mlwuOFqpbx+tabTE6TvOGKI93vgNr42J4tnOIDaTbsTstb0rrKsf+7dm8kXHRkWgjPyS4TzCs4C
G7vU43ROqdIaY3YIhX/IoyeBJUGpVHRwDVyIElqtyEnxxHfIf3pJbuAcDQ1GIObHPOfopnyevibV
6LgZJbWWMbzDXM09y7i4HALvaQHctvzSv+uaXdIO/Wmx/zjXNhCISNOoLMwFu5t4NeqOllP7zn0s
kcRCxziwGV3H4nf3d1RIhr+iKvGlKSzraYCW/AnaspgKA5Ijr5ZCh0S14AvlQU4ZnmsqMOgxjDjl
jjj+oDOf6NxicGXBcyuyTrKAx4uTbHMPIjiY6RKYP4lbdp4SmmM2iIXHfOt+4y/BPxby1kcbmGg6
EwuFNq+tpdgB/NYfHer39jsK/n2xXfwgATBUkkFVmvnC5iyE/qrb5S91108CnjZbUXkiERQq+BTk
AGuEWddQv7obt3LCU31a1zrMmwnRu6PXe30LnD8GoGiZ4exMbufzv+81L5EwaNdzqOxWMlvK3uCS
OYzGA4m0Q0DKDKn5HvABl5MxlVDNKC31jOhU5IjUS35PH8tiiX1Ng/GlpSylUnw0Bs7WmzHDH2MH
j1q2EvRNdT6XV3gzOiQFIZgf0KZfboTXWJnwkHiwqg0MLAFHh/wTmDqQdZKJX9kd0fd9cjkGNSgp
93Cc2zR4J+LQIg5AwfHgD71p1oHjps2qQXC1y8JUeXR+lVXuNBPu3DFttd5idgkc5S+Y45D4H2XZ
dmMBUWh/JKt/sPXGzFx4oyLV9ozldZShPwxeS33pvZh+BtHd794MhzADHhdxL42YzpB+eqbeT1sE
SdEI61WcPvXhoBBdNARoC3Rzl1xF++DBA+5yG8jiNIZFPLKDScBZ6lpZpv3w293sRgqLn3NLN/Xw
Zz4bwsbJuJrBhhEb5nyz/xkX3jh3eq6lSH8QWOuXYV91MdxYFRUk0hvaxIvF7853+yWRgpXc7UTz
aKqVKciuZGxJAk1E4FV3nBBLUWLJLjNFgampmpGc/xz7THD+22nZNpo6iMUY9FoE1FB1U0LBQD0Y
PU3lp4um+HGpwzRhgZsBqKQia6LP6nlLrwTYR3O6ECz252UxXUlgYpTyiSU3D9+2lhMKmj5XzYQl
TPlTp0GhDLA8AfqwGaUPrSJm+5jHcerupDvbS4XwlkLkZghm5Q/dYVUJrkua6iKuzbAiXk4Z+ziH
OEmWKuLMSQmm3w7yoABF+S6VlrocAAL7dDWMZthgDzny7QlVQFYnDrO/NoGGFNtha6kFwA3t6+v8
T/zT7FW+4eWYycl13+pi7/ztR6xFwrSLwOS+SgPYt0qvf2KRTz9v8ylJecJ5UUyPuVL38VkRRNs8
J3qDy1xGDjh73fZhdnmCdYUezZRXwJnd/k0w9fmpSoxjnZN6OL6+dO7hUXGCbVfJtQLMuj99wCdq
KtIpWX7LXXpW6R9139ewWbzwrKSFdSaBJGqfzX6+MPjwoiymiploLDYt2jQmjKQC696BhHs+VXIu
XCbK9jh2Qo7ZJHf1pAkQ/vJ1VByPd0o28PKvkxSovEUl8TbwZh4O1ZIyJhoJu2OTkKASzrJrCMbX
KFsrFsaubUZG3aJRWygDGlKuAXSm0U4BJZ4agaEO7foPZRgCuuvgEx2ImcZAX7Uy45OBGjgVyHPM
6ma7fAmatCVSfCTyBKRtkFEbHEtFwocSd3D1r4jbatLwDJ1Ovxkre6BRqjR8xwNTAHEpNcIrOENF
u7XkNHKJkIJ5Z5KtkDFf94J/n5jaZEXzsV7KHF3gbJEL6mVaVyupCatuKC/dTrUWkXSitER61oDA
tYmsRyXIsAMrOujY/Gb46hOdTq3C0Gp4jx7Kglb1Co41Y9mqn95RQWuVNfeNiCRkAF314YAKWJnF
SQi2Ln7pfrl8y0J1ZfGkIqaW1pBr1szea4eVjvLjnm//aByxyh98BcLLbXFLwdPNIYck1fjSGidr
2pzilX3V15g84NjYwCSfAkyKDgAp+x7STIP1e5wy9ZwQbllABUuViUy8+LwdcVnA//9yCmcrXHf4
LDUBzzm7A6kdRavJxUJ5dvPRYObVsn7JHKveKWXFXVIhqvOUB4oNUZ5t3vdSmkqb32FAwHjf9MD+
CdHR2x16uj/ruf0HV+JoZ7hD2WypUKmysuPuJ3O2wyB5nOmh+JI9FDOqibx5spYu+pUsOkb4ooT0
74eFZoE5Clr1O6bb5zZMKw0XUdh/DK8VGtOxS2omSUqxAGV9l5Hnv3I0Zp5vId1NPiuNS/kskojx
gzrXlIx7F0i9dXMUaYcMVhEmwoDlS3KkGMSPA/aXHMP2E7Z177kYEfCC4jHcJxlzDDCqPxoMbpOQ
+ek61mZLa53gRlseZS6lR0PWY+xECD3ml6cj2rqy4ipc66/6bTj/8ipKRD0fb5oT7xjJ6N4RpAuV
Wc3r69S3UliJETmwFbYsjDHSYr5wbgcwQWTNWjG2c2rnyiOQ6tD5e/9OT1UiXeQBjdV1cXAFhfDi
B5f+lqEvfvJagvWYwIeZUne+Yx38h/hDEx2kiWBpszdecyiO+CftJa/LSDpHSxeEsCBnwUfAp4ng
gMhuITX9g0qWbnhn6puBHRVnAoy70WI0z7VbbncT1nZW0r6grR3wTbqTu7Vfm8goMr84/EZDSbPF
lS/1UoDN3HsjEXLVyCRPWaBsPzYnB26TqV7JcI50BSujvvvYkl9KGg8FzEjvDhKDvdHUeRtXDPX7
ISa0w9kiXl6+cUf4l33JF+jhH2YaG5B1Xvm/DGR5eThToW/O15R4M3lufCeloTnZHsY/SfmGmy6o
SSKpwZmvyUQeS/fgSuc3/4zQYwzK3xU84ZLXFGrZl9wVvijLP1bPbFxiQFeqnSHOVeTD6z5BDcxr
GIMPZxF2k2kvzBuCS60LOWTGnfa0+rvikd2F84Je5xUtqAK+8o88KoXgeInqPJoQ+AYtpqFZUhJG
yGED9VjQUYbN/hXcymnsLjGnsEtnnLCm3PvKf6S6EV/cFpsQKlyfaf5qB0tgIJOOG2OGN7XPgs/a
KuZSmR+QgmRwGc18qZUS4+b/AZHYFnjjUHmvgxI7+bsgLg6ZAFR/bVf3F6P/mYKz1DgIf/dF+w2V
1N0jVhiM26ODpHX1+558vJQk4++83FV9EnFYk1FXhwON9pqIOJ5kJyQix8H9FngC2jy+H7XwINw4
yvFIGzeTJGCmjrqOfJjbST2D9PRsohBlTcmjn+vw9hrZkdFnPRwC1+F2yF74QAd1PvrshUz2hy0D
lRkzi4+qn25d5h9IygstB0ELIFWX36+yV9BEBcaqu0zbRm/trs3whF+itwfDHbZ4Mb9tWY1bP6Fc
vyCJ0pWPLpz5HGNFC441ZRm2BzWNhtP9/BTO2Dss3X6K8uPre8uzd1K9TZ7K1sE/BuZw+h63MWnx
xJANbS4xSi4iVIPvIql5jGuxKHR83hUyKucYuS6FOcvwN4naPAb+fZVgBcWvh9rKr9g6SMtRwR18
P/Il6uJBe4lIGspsM4M76/RAJcgyhHKJ1B+Vdzr7KIL5fjhAsY9x9ac0yaKDLfZaM90zrJOjHVKV
BjVnlxPHUu5Mm/NEsZVZGK8N6ea0w1vZ8c2uTX53JEXEcuw4kYJCJpMZFIS6tN1cF7ucyfHIhhJF
Qf43oXOssNrOoOyuOJxnc4KAD3SSZovkpq3QW7e3WFyX8YTgC7k4Fzn0gZm4ldLheVyQF6tZ+8zP
7RHIoUdoXnXsO20ACUddIQm4bDU/QeFcUHLvFEgCJeQUKj56JKdFRDPie8xAP1NYKEGJWPyqGk3w
sZ1/eEs7S89wjQXOeed3Kov7hxVGi6kXPUWpPJ/Pls4UvWBGxlCIzdG8tZHsZljCkZyEPLLdmfJV
mOMC7rOivpOz2/XGEFGkTYnTVJc9FpG7J92dOdlJeGy5CrEFbzLM8/x3SClYbOH6Qz3452qCW6Je
qTWAw3D1kcyZjGeh5E2NVTxuJSHYAwIey3rZfryKrAR871K6p5s44EKU1fvrw2ribUSosPVtCiXF
sG0i7Z8gcCs9nM1UBt2pntWTMjChwXbrUSrZZYOJIo7JBUPgDvdpgLwGGCrLTfL9pAVYv4zZiK2E
pgKbZtMjcEQ5mforWQa51BtoQBvTd22vU9E/d4vVDMasvPihxHcv0MrvyaykX3yBfE1YFEN7Pp40
CbR4dX+DxKhUPKfBFjYPfkVi1xooNUy3ECZ+0pBfzqCot3kZ23Fe0suDawKIW91dqzJl5AqlColk
zbpc4t3JwAdqaqzDzJnGoPqq2VqoHbiT84fVPxJT06/z/xJF4dvnHdfdGwdG7essnRvUQ8tQ8Gec
JZwUxJR/G3ZFbXofTVuUboas9n2ut0O+AQyUWVAT5YueEOHn+BEb6DsDHLh0MTTW/g7kgGCJKkwh
RjqViCpALARZEok/2p75Pb079jJjypK+PkdgwX1kWm3KCbiAFwgOtu72oThmfLNy99Kgp5fm3Jcv
PckWUCYUVKIdYsfd+bSPErYRwRRwptGgGqz7eoQnTkgsCg+k7CM9tRP35uPgyO8cuYzM5BVdPwqa
skjwSnWvuUTm05+TsWxtzHmkaCUfDHdCVtqbFqzG5/qZcNNyyohgLDPmrsXejCRAnfzVALmcbb0A
cE00Qp2h4s7vqPfAMZVKhMGLASMjEiiXHJddr8Mt9+cX9rTIjb/+FgEa5wQAXwcXi1qgKlbA28ED
JdJTUBY/Nf3LXCmTKrg3UShu7wJqX/ZtHZ1U1WG1mtp2krc2VhM5RNsX/R9G9l53lTV29nHkJKOn
AbhPo1tmJoLmE/+Nf0QikvbbN45oliQ74tFe6j90b236TQ2hXkgELOCxbD/rJR/mn01LKUxHMU6P
SeHfC9nrtQW0SslDNCf87eDYEPwbTYrNqfADKx8nMMcezfjMC4CSLyGD1CnOf4KUeHR1dDxIusYa
JyWbyQdmtDYykul6JbVDwkvgnuavZnpxz4Tw62/PB8sAV3kN/8UMruTVpqbht4n5NgZLQu5m+uio
/ZgcjXE2sUtTV2MvGYdmjCyf6PQVKEpEtF++zQ3vXHRUofctvOeR1FIuu0YpCUEjwYOh4w291E3M
LV29wtDnzSH30roTZxossTWpo77G1KN0+RZ6XuK5GqZ8M7VdJSiLWXZUzM/RwYwFKk5QIwvZXKDK
XMt6QLF7ir5cJPs+yt/aVnyDuDKnJEv72mkQGhSLVxPF9NqMslemQgf/EFzUDq3xiYHGnUiWnEiS
mYyYNbEiFZAPXuyf31YdbqDuRN3gzmw7yYudtuVLO9YBAs6EUOXaPi1Kzmr+MTQF3MoleQfYsqxf
6ondrM8DvJsU5K3Jpl8K1PrY5LAT/lB2/K0gSNUEhaVIA0eTw0P4/sAhGGFKMmyr27Od5wE6nLRt
8Kxm+8+3HosfNEcoS7M3vlUU3hIuYXBt6smoPeQm3q/HV0f14Li0zfQVQEX24XkYJYiiJ0u+QNe9
pjXquq0enrWm8iGv5a0eZGfpT8h67wVim3NWXXjj+wt4fQ9cbyPA/somaK8e/B4aEYIpxs0dQigV
y6BdScjg9xeNm+5Asuq8zcdpETvA6NFgiIu1ZymTghnbFUIsJT1V5NhXecViA/ENIBFaLbVB0cig
U9sQSqsmfhoUQYPSdDv/eMSyglipaJAn5Qi2a+/tbK/gZLil3l/Fe1qrGLvdreqKvq7TNGe/6T3w
0yzf+gE75ejXTr2m0vxTKsHTSYHQvDf8ZSNw4wMPshTKNzBpBdokB4/3Mu/EPeH8jF4fqjTpLHq/
ZmgZnTunAI1GJBfrlIm+54etGu1i2pUKAGyJnPMKxqqxp0Cm+MkB/Fh0xnN4/hfxF/1f2afrQfaT
XmAhauuDeeamR5HEV1+9jLgkQ/5H/486uSzJYvsDMV+akVmNty2UifVAFS1xL8GKyiijLOWf9Pqe
IBqtACe4kVZo5/VoKT67eU72TxXl86aRgkF35lKmueJ7EryC6hroNj75Fuxr7f6SQSmHuZ0VOP9b
8vRi0DXjrxMekYm31SelvPYK6ySJJjI0gyD9mxxmwkYmm6x4FCkIlgmqbNuADN0T0HH+Heaz+iu3
YWJH6DsHlxfE4gUl4EuyDW2jHrJN0b+PUPi5XekthZFAL2vlVd5F3QwKPDZgCpMCHnErGEBwrBIC
LwHCoRxbujf6zWeSxPsmJXHNPC+Aik3ampT1wfOeX0YTWbpLkNc2gUZWxACzWnx8I3NOWdOhFQNL
divgrmuKQ+6DDTzikEVMAHYgivoebWpm51AYNmD1z16VAl8zxjTDw8KWMvKwjuDLw8X9w8SUng1F
bvOdQKJv11AkcOIcglHnWRTxVeSRvrFEWilackAxbWdZykFimHKjJbN6o/9nPrk3zdM9IQpjYLy1
9HWEgEvCE0KshCq4sm37JbNpcpwcPjXIK7nFeuVK9Yh0IojjjXfIz+BLG4dXbs/3S3FNUukYZk1C
i6i7fRDobMxgey5JOEvoGQoHBcKFyrd8w6hnC3Tqvek/HGZN+0C6Nq3tH79qba/1YCx25opxkzO5
amcxSuybdGF/NbUF2+ykvb1Ld+clpLC5RH6MkIF8EDN1rgZOLzQMZvWb2IDmJ/ER0JEj7CYrqDzQ
ZWcQPPg5Ljy+ryilOT/qyoYWw3hLWYwylhKtv7WfJT0hcaOJaKfakx6yhuQZr4pHSZpjgCWg4YN0
DVVkUdmE5umxbxqWVs7/XRC3FY9lxktiTp5c7NoZOntFhzSO6CUorUgMXkgaZidO7JJInhZEVdyx
bzWeg+RG6AXxrbZMvhzsj4FOJHADoQCTGImPkmkRxxlsmhaXhjHBEH2Q7CN8CsEcYBinVORve7jF
iCvt2wXCgGglCEqwtGcxiC2ULqrFs9gaWMqJNbmHawlGGwlndAJBqPAenxJPAEHrGGWWe1J2t4M9
feMcPJN3NpdA+tBYkb+ptuIN9XdntdddtSqJcOWLOocTt32QbSJN+R/le4XGwQpsiKtYvEQXzKRn
WdQrg477tuRCKQ4LWHsttALlUtu1NHR0hJ/Q7FPn/TNZva0pERPLc6UVDHnc8ClU8XMXJZx4jXRn
oG9+W1BLwCpbXUUbDbF7V34SIapYKNJQMNHVuXiIjUoJl2QlzQoFke9/3iCaCQt6+7ZaaO9EYs64
B8kENYe+Xns/hyWOIt/deBhIjqBF6yZFDiwaz5NYGNfVfJx1/Dm+Gtj934hwfljLOpenRHJK3mhs
DHlfr4EHtS+JjVx/chtpc6L6jAASSWvo9ZOw7kDmmdjuF4gSuCgLxqeEfCmG6ZZLUBX8uBYxX1rU
5+6l5ea/QETnt+Hvv1e6j+f6eUDeVyrFrj7zBd0Cms+fm+bPhSiP4KiVI+0PMNVHDh7kAhpGXm0D
4nqYiDAoNEyE46dua2IYyilZdx3Yd1RloCuLdWTAiSFoB6smQUwTexy2+yuZgKsbonK46p31lb9G
B8vHix5AzqdRaXZxrw5ZujUWmRGJ+Zf9WA/2zAVNUOxBDETM66f1eACSSYI0P1SeaaCI0WUKG/Nc
gpNhidwVctz3r8lllJYtGWFoyag5YeRQcstDK1sVEqMHrcDBxmcfqri/+0evd7QSxvMzolVBh6ye
HvM66NpJmkXtPlCWsCmpHpU6Z0BBUHsHHpPApZsAq6WVZijxWcMsvzOT0eoyQ1k3cqH2UN+6ulKq
TwZAuS7J57TC2yV/oNxTY1B+2eX9ntzAhPUYNe4imlVQlKUil6imI5i/ZtXx8sjKJUOSpSdB9cLc
Y3yk+mmGoJTIn7s7wkt+TQT1Wgk+bdaqfSt1BVmuQ2ak4BJZa4sZO6DwqrizkOQ+glPWYCAKT8Z0
QUVNsK4nI14zMPGvyWPohXHXM4vbM68M+mA475tdgcAjTuflS/Tjsf0uTfGyttrNQK+K+27Yvjql
yOqsAZzmOPgYaITHh3HE2Z4VZbudug3ri0ZO0omQNQIgUwIGAaoGMvsGybotRU+yQLFUVkF/jtja
1avrtCy3tICNawqDplIqtl3do2GsYFIbtTXISbEz0Wm3T2MilpgOPNJxn+6a0hTd1REz6lliDZ6Z
id/3ndI9DjwJQ23Vba2fAnpwG+WYlqqnwvIW2E1Xy4Kfe9+x1HrYZbN/RtjEMWCmxXMrtUto9lpi
vCXZiAWTBxvjFHbHN+qUvPHCcts8bejhJcf5GqM/yurVliGhtpLYgLP7WDro9UHh1w33tFZ6T6TD
EVI+yfL9CFeQRXCsDPUmubOflL1pKlI17avy06ZC4MqJuws74cuizx1pWTvHcDRpbzkgzbmlYCLF
98YIgxj8GSLl6bNXolvsikfxWZY4vLiwDDqXbhzQ4u9STtSslXbtse0oww0xksPDAPd7xRLDG3Y2
N+yfUb5hTELasDpByPx51DqlSNPYKRlGQHUmTO1IfbmkpahTEqjKYMdrsV3dw+pBccivJ6Jyhy+i
DcdvzJeqy7Tkcd4puorkStugXUvH7Wu/S+EykHG0sty6Tva8/m3zadlk5iIEABGGHvhjZgCAnRXt
NgUn7W+ec7aEqHsfLBo7NMWBiiB5JZdheUEEp11T9ABPvdkYAE65RF2l70x2Vx1ogV0iRp0YTLT9
tkpp2JeMnt/5cZyAMF8lf/YZXOL65PdI9ob0/QUEThmGqNq587AcD7K7Xm4C/UOLYH4aZ7yPKF0i
kMKBuzWLC/Hz705/AvHd4j+95ROzNyWKSxF+GC1ZtZy8sWGh3ksriEMXJVdj7LIKY0/Njm+ik2JG
9SJMj3ZDNo6eHiZ1tZFQD8NDtaWHlar3jnv3KpQCClzTOm1YNStUpXzBln1p+km2XfxEY7BWrUxH
NjYVqu3QZz9GK/ICL1SlKiz7BpNhV5E7uzzAkySMa8whR+zoZOd1VYFNH4kA2crIa6CdoUZU3X5e
0AJXCIiQBWbettSR/eArgV7X17Eex3a4f9bD3Gxr/ZmfXlkGOftoarULPG1tcPsoT+xRnQ2iHE30
9Sl4ASpt+2hFrjC4pDaCe20lCwkeZgxyeKSmtivDo254hHGlwYd1XlX7A5cmF1d2t9xB1KXicixP
fZKbV8usoadpdIBCDrLCoCCrSbD9iQsh+Rf2NxCIPSgCISKCS7qWkg7xMSyLV7cYiUFYRqw7F5zc
7reGhGCsIHBNH+ju07gQ4pwzfe1Bz3pva2p3g1DjKOuVEMK0bxNqg52Jc8uVhUZ6dhlLuDhJMnaV
vKiY1u2tHTlWHGiNIBVfWRT8g2zlcW7Fa1A/+A7SsIZOK0C2f8XXH3I5AlhD/b0Zc5vD/6+pdZC9
4gmyj9c1BYgKsStfK8OA9nmtsgmHedGAQYO34GxuQdTUsS8e2Boj6gyX6B6yixaa+jNw6xvKaeTy
KplRQ3Pj6J41Xi44Tg79MldMRyeUDq3Wft+Olhwu83YAPInmySm0bbWyqF6JKPRBRj8CiJpe5gD+
icO36QiHD5VLG/N3AKlnMQ0rvoQ6yFh8ffYv0Pm517MZV7Kc595pjeXMJKPqxJwOW5VTGGw/CdY4
kFU9/OY3Q8qXarWwRmUgCFhhjQEX8nJDB0twRS1qP6Es8M86b0SqReUwWTtwXq6VehASaXpiHp+X
9Nb6TYBYPzEqAUh71Ud4P0vLntWYtQLd3o6dHle/1V51MNdcvQ9uQz1O/MsP2LiOk+ACtMVcWz2j
y9P9AHiYkUgua6nHWKYujk0PJFIn5hlPFAXrJuF0MKNLpqR9mEkqX7bgmjWR9nXt2QWgkB0VXLNc
A9sQ7AXvCO9S/khu5R7zza3dUMPoupdD1STdPgOeJ6CzDbyblR17+H8eYh9VEFFgq8sXdKUdv8/m
9uZEvfMazxNTC7xvhusGo5Q4fq8E4cMiHdEsD0TqG0baW4NFC8fqMtHT4EU1QxGCtVe6/AIxhNxo
w0TfbNFd87DmIf7EAVI4R54cockvChTIi7TuSKbr/m1VDreUxfzA0uOw2/7KuPz8eZUnCNS6y7Fs
qSYDnjU26RvKEUBdMZhB6dqhH9evJCNvpVZvC5oyNuQ+VOyIhe3HERg02/bkGYDuwimaxRUeZmMt
iWwimVGJgl1cPFsTRmdB7sKdGeDp3sagHxqIQquSA8Ny56rKkYLrNYZ/O1mXaT+1LJ13Le2bzeN1
vHpdtKjb7vl+LNIAQzAzEoKHWLlhb/Bw75BW228r+icOgGOoezknPgXHoEmpFWwURA0rMLVEFCE8
COdxKE5/V5mgQPljaNJPO7ZJ+ixQxqe2kBJBZXQQkD5y8VjEQtnKfsOBe5QxDNlzAvvOecC1vE1y
xgNIW6d8YEnFuwudXYigAT+eIMaXxV97HoYm3vl1WjNys/NqOfQ+hg+DYeaVfQlEwmNg3hsi7hBs
Z9N21ZIyZWEstPqx2KZ1N46cL2h3ccJc9AZduh6vSELAm035AK5q1jv+V9R7qCcBmAG0UkKjX7lL
kCScc2nKYkm6C2AodNdCSW8HVz0smPDMquQnzK1lZxaIyUKC3DsFqvrAbCQCHrTpjO5QtUHMb8Xu
h5yXVF6Tbpv6wVF4TOSgnuaDogsI8vjt2rG1ZP+jDfHw7rDPcsQ2aGgE8LkGol+tJk2JESSJc3dv
m4UPcJvrDA5FYzQTi1gVF3wFCyHS8+Wv2PUUzcbZtJiJbBpDNBFpW7vkW9uSXwDb1tG7H693v6kU
YzCP5QctHFIhRfFyuqMNw8Q7+EAdurPmL/UbviIImnc/5tX644gbUdkORtsUWRrIvMyrquLhgS5K
5o4ff0Vop0UHEJYMe8kibhsGP1585xGVP0Nsz/iUWQodDEaR0KDefwX9l0Elo8rjW+Aj8rRceFTn
pqQL96y0FkRwZLjY7U0+Yxxvz4Bl9QApJsqvKdakIBQYlsjNE7NkYBUaxgoAr3yhuEpcI/WiLNQt
G+S4JyoXYOt1srk1SeBtW+VJzhn2/MGamctTgwOodyHFX+Ih96p0dxfqfAUbZ2ZxFf471xJlN8Yw
eNxcrPkfTZ5Y4DGaa9UyRWC2nlGrOm3400yr+ear0R1dwoOra2RglZfNw97nfEY/xraIvIunwR0J
AdcmezMzMbsaiKOGBUhCTQg8A9a+vJAYMqO9voV2cYW/YfSJeFFrva1yr1KjDQkPCdcN553OpqWC
SJ2ednnJfoprfQ/xeDi2q8mpMWy/bCjh3ERUoP7R0/M+tLxPrLCqOz8uuO4PWN/sfJWNMMpN94sh
b8MgGqNHNYd6NfR8wxuO9wlgg+5C6BXC3VnV3Atqn/CWHL3X27e1JB/LwhTaw8s2vs/ps5MPvqbx
PNm6MBsMHnER4ab+HuAlEM0T/tn8KcqVApizuhwDHB2AKJk0YEh+oo95wzus7Slobn+XQ7JSQiKk
TD5A/7PGYJ/YQ0w9yTeX9zGavHGuQwG55uF3y0Xu2hmGxw3lJF48PI3rhSXXSkVmdd54puNxrn92
2eUOalEFHxkQ0NU6AX8FdusoOFJ0VlLChB7AwK4/NTZADSay++/dwRoT/aKpiBC4B1o05XsiGCSc
EDk+ddUOyAbXjWkxlI2BxzkL8ObBD1WNw8H5SchrntRzXUsoobVna3lss3s4HJrn/tXGR4bSAKLk
0kJm4OzP5t6EsT4NhYLOZj7mMut6s67dRwTrWz6bRWMZqCRL9rmcLX76Q96PHlJI8rzl+ay7XzK9
lLoc9WPtBZI5/Db3mUftBwqLq6gsE5b8QKErAj88ibqu2tLAXyYxQE2gIyvsi0tartsSSatkYpra
KNYqzJg8V/E4eWqnlbiC/YiAtSExUaijnBIgooZB6GESA4ZEyKqkdjc6kdTbvLTpXZWDKWyMXZRv
nabESt2j79vgIEyp9lDTkTodeO9YREwSVZfbbsiVJdVDR1zX4ZDl+PFvab7Y5xNvPkeLl21SM+1a
XNXEGyS4T+YdoUQeQIqyQbU1rPC1PV0E3rnJtVGbnCav7dowBdp6XNWNIYkasAw4Iq21Pn9oqJlH
Jgug+WaH7EiO3GjXCB9adJsP7RhWzor7m8QAPSPrpXzRQ63S7C8f79Xxg8MgheuGG41UBIRLViaH
X45C4G0GDgQciz9kn7JxEl8snEFav9FrbcO56TP79e6xHiHw+DLuqFWMNSNB+0nBl38h/p7S4du8
IAKWm0iBUsyAr9OFaGoJpJhsqERXgmXiItT6fPmNbraKg73S4S3sEIwkeCrUxQrSeboWAN00ui/8
MTGlRznsNK9PDSwHSxMfnFMLatBPYk1T7Z8yKS+M099quU7UKwkITNl+LK+JHe23ryDLuQ+MwNiu
qMYlRoQEwrgZbVV/31jPiwiI5QW3oXjItDHKtt5/yMbXtk5dfKaxpoyp6fXHhkAEwMxD8KlPu/Ww
Z/8zQIl+BBpTYkYXzce2JrHFzDdAA19McRh4cVxhIdFq9/OCwWseIeyQoYafzjWXJGGoUNUIZ+A5
Hz9ZSH7noV6tFHAZtJ77RlYBKbDEbEhwHa+sA/6cPH4yyPp6A3PzpvIA/VlOixJNDBbmifyiN3Xr
zYUn9FsHo1M/kc/7atSYNne/k853tvKnYh3MwW9dnaSZoZAOu/gs2hG59G5NFlpE/68ykySGf2dh
QJHCkrjOg9QFAHLEM2oi9iMyv0r1etzdhj4wBuWXxw/dK93ws4sUfAjmFgrI+dukVDnT8OxRuTAn
oTj2i7SJEZGqHt6GUeDGxI89G6fIAAu+Y3I1iczzgKcDAnoxGOzddXx2joD24I1+hbpgE6axhNn8
n/E1d47ZEV+hrGDTZnBPXrBCugWu4lL5TIM8KOsd0UG9Sdv6Qp+gz/2QVbJk61my7kMVjbrFIBMl
MLFaSycRMqYPRFHoig0ZPDJi6CVQqlFvlF7UCV3XTQ1jqcJ/FBIun4FxZqLCiVm0762MkKp3ktW0
59JOlKdSD8KErMFbl86299G68IsXszjuFv0YNS1xz5BnTN/8nPxs3/kC2XGiWiPh/vtBlFtvrmJW
wdZjRtMdEOZJg1vsH0Wa8l7P7Qi5LTBe5aNPSJhTJL3rXcmspozkgGsNW4r5UIPJpzzK8mIShK7S
qnKeBMkJtror8+1DdKprE3zGO/mbY9KmYSt9eiZtj2L//4FXQT3OXPyUGKNlvtZrA3Bu52syWJgp
dV/YuLyK6VGni+Aa18Oj7Bay7IA8ZpUmboO7M3nfm3sQRjfrgPRqeU87nMAWDzYhhzncQwOhxofv
Z/LW4u28MJsrH8A7Q9CuzroKXfMVLrLhnsf5Unnmy8fUd1dEDX91fAJEjGmPKCsbVzedfZtFyTrG
u5U4G0OhwvnUKEj60mP8wWBwYumyplli+NCyAl3MbGIzMcUTOTqBanKHTMWeCPDacfBnnBIXsY/1
5M3lk0HXOQssJfG4eP/AoesISiBaF+TPQduG1lry+R8stM2BbGERxTGs49KrYAhLSpYju26vGQmQ
Iuo8cf2dh9tn+Ej6JQJ8JNk9mPpoOhXvltV0mZhNnWrshgRkGZguxBw8iHSVFF2zwn7QqRhJWxWT
fbX+kAp2H99/dlOhC/Xk44on0gV1v8sMeT37QAqEIFlmbQkNW+Wxsrm7z0U7U1PjinweWAmVRftO
YmousLmFrfgiN8HYs8NV11uGZQWETae3zAbOLZ8AqEUT2aqpCxVkWDO1+41WkXKmSbKJLSbBf4El
QKfl+J08K5jP7yFPIMXBoe2K6TlvuWmADkjI/bCH66UcYdrpbpia2Ef0rh5zKUCzTrPHESlSm6OX
9fbw0K6+XgoWQolczd3VHehqIPbopNWgipu+VyQvd031WnN+4OTAEkHVt6hdt85Awl4t+hoOmas+
p56Y0Yb+N69kOJ64yH6TZ8CSQryeP715vQ0HWq186AVKAP9AuBOuyrn9sjKrbisAwJKw7Bo4Njnl
6xx7g9c/hrkGHdVs+Mxuw32WuJyCgGNviuQhAkjMaVWrHjM5OXWowLCHD2yXPQBw021P1/8n7LJP
XL3equGc6js9dULabawyCbIjrxTh5i7nPc9YNyFQrcCHfhFvuA6PmrJ0VbEmEL03SRKh0Op6EFCe
vn8qt0R22PN7BE8K7bPbTzakDdBiRWZtK5FldeXDyfFbMOm2+huYxx7+v4Ajcx/Z8oH6TtIwmkZj
McSOIylQ+WufDiMkL0XH9EmgxnoGozwuRjJZgyRUDuFTOQciot9FPh+wpwu7eA+KVxmYe0AOqzS1
zoNRxdND2JN/yj9e5Rho+0QuQRjRmkHRBDZmufosvKs6mzTcvh1OYzu5exu0cEbtrvRIFvon/+iY
Pz7u4cza9+j9GA5zJafxTw7S1wcqP3zYB6KG8tyb9xKMb/yHsH5WevhoMDJENSxIQfFlSb71GdOJ
oiJAzP7A+oVDRHIFjob61EHTIPLs5E1l7mbJxiQgB4mFl912xbO6kvB2vVoql8P9EVp1pmD7Q7YB
zds5xPrf3wd6YRfN6SNrrbgkKZVb0kbFHv9HXODKhs8/xte+ZWmOrFSC0UsRwZYZbqfeAaYJoFZU
3qZo8Lhuzb+aXT3IPUrx+BZYZSzPXNLiOqo2a7jSrRvPN67S92li+FpqCNK6Gufs24fRk2OSGp65
OybC2Lvs4gKg4KWAtTmOlTSCXBv6QVtMWBI8DRofs0splpKIg9xE+ZCG7MN2XxhxMAoPdbViZ6wp
00MxYcBhuRoSSS/+kEtYyaacxnSFP58lsF4jxWKQ0qs0cWMV7fURdXSJwmOsjkrHS9dmPO0rV7l7
AlBLI8tEHyYtHPLEtzJjBcUZYG9fZ52AfUwB200IOSn/1zm34J9qP4D5RwYrJR6iqVD6/0ePbK79
0Zps0EldefgWa0k/bK4h7p2+ep9O8ZseNbsblmy51OS1pZ/32aAczvMwraH9SFrQFnkKIcHYgAEU
NfoBQV1/yQFx75GbEtlrbyxYPlbJk3u3AclIt7M94n/quyWm8z70IYTticcn6mb7BUkzlahE1q3C
ZZO1DsIdqvneTxurmJLKjh1Xvl0mgb91/4H/QIKC0pX1qEaqpqzxH18/m/qD79S1uZ4yBDXr1s3m
9HSQ0Li6f9PvirQ9ZHEPtEaeHaDaKdQWeYjHtZF57YrpcoQE0bVdidvycC3CLh47H/64HLVC0dN9
hSDKT3Qh0pctc9UD6Vvr1NEtoL/8x+lv3hZUBjsPVoqk0LmhtbwncQcwOcNlx/C3s6gOAJ3jdVlp
wZ9zMLEzsHI2Wmo+YkXozef74/pFdnqoT5qHxEguX1/t7a+6AcsXI9LlMLq1/6B0tcQivUHtmyFq
5GkdVO3ocmHAWfTABpfA77qAWSGJmj0e4JMpzooo4LwNj7pr0K40qCKZnrTFCknBB0MKPc62ltMG
QqFUyxSy2Ac0nknHnka58MoZejFxJ7MNqTNaUXqHxCcPbjTjlfakjW87GELILnnmfDtpC/CB1dgV
BOLbluXGcn8LQZ2qZrwVHrC8fEre6+JH5deDn9OpgNU4GRFzVhAbPinQLpKvp26Hl7wQ1t1V8ZDw
z92dMT3dZBxl9O6G+YffdgFgCn+rDD5pA/tWP1Kk6wDYMYPjqi3RulzIW02FVR4eO6cYCMZNe+ae
K9FuiwKVYtyUO5Rn9ybo9yUYZSAxZ5dN1i4V9lDNWbdtyebne8m4V/hIaHBkIY22J4U+Paa+7ivA
9fxaUYeOLhKs/sLmd8/egBoWbDscPW1JjNBnfKELOlObtwbKQlOz6gIOi6pr58+tphZbndrdezeo
nCrK9wyXXkxeQPHRgLdDdeH59ifI52fLWkDyVdD6FCJ3L5lRN1RhYs3eKR9rbat6AKG2EKmVmmd3
J3+qXH0d0t+PyopXAJGTupK93Q9Y8AzMry8jC6Lbn2W0PAvk5fykloogj97PavaDUNLbQ+f4MB+/
c45NM7shPjIgafFgvIn7zU/lz+w5ChMdJSCzzyQxOVWVuDzkLuctGpUoVlN9Bdcgpj+3uu3zTQaU
BJYuNfpKdfMHhYy95yLYE6ygJ7Noqitb4IYKOGHPR/juPP4F+waaM/dVU/mDip/FrvCUii5PqtcF
bCDsq/zWuddx34OFZ4Ai+yGA6VeTOZOiCA23rCI888QQ2RfXsyG8XVU2TUYVnGrwpfkt35sF/1it
pQXfrwNzGYT8bM5gzJSZeSi1Na8ScyijgO3X8+/DYUt1sv1IzkZj5Y9Zop6hGLBT+fMFAVwD385C
C5SZBAOOT1QU8OgYOjj5A9ys1HKeS4MJyerjje/t1K8N01wP/uNORNHYDG6HGwNDxUzA5c0gn5OT
b/RKOxswM4Lk0NyfJ0eyAEyKIE+8ZGpvEFZqB2AINWvhkRIc9c/tWhgJxmRio6y58TrClXGC9F3o
iXCCv7cGsJHb5RNlUsqhN2KBzr9h4Dps/C0uJJCMI281uyMPY4E927lwHvXuzTvbYZkeogSa6eZh
zil3FqTj31ZjgZ63OfXnEwJtA6sRKVSyM7q6HNrQk86r7p08koGx0CayOJtPz97z5y5vsBXTEnsH
9yZo+SIwdWsZhOvjQOac1LdlAshj+rV3c/1OqKog/+TcRbJOS06Bbk0c/Mf0e38UuYNU2jPsc3N0
hEv4Nzx2C4PbTsY99O0atU8RipYohDuTp2aQZ39Olr8SDX+IuZa+KjRX9osun4a0LPbMmjroyshA
we4mR8HNRY6krwb3pCg+MjEpZfw5gSybfZdVPKfO3944wm1B2KLBI0aWPTEIL3aWaD1FoJHgg9vy
SgZJSe61H72Sfj7A3JUuR6ayS7iZM3DxCHiA9RdpvS7008jciJ80f3iXhOlEef/gJD4aDxrC/Qwb
VoH2y+gCKD7/0L1sX9MxAHpFQR0t+XOMAIEp0/geCQQvizJ32ZaiJPTZwI9VXEvX0eqw5GtQZ6rs
4QuTgysGNAM66mvBflDnQOI6SipZWI1xvFOJHaAiMMqC+gN9cgZ27f1zpu8jP9f2kCKBZdWO7WRZ
6K3d9gsXyi21myFovGcTlJYS4wjVH4G6uk7imbVOCbTO5+awfvsWrqfOm0BnuW8xBiYsRj4V0heH
4pI8gHfk36EaBR2u+rj44RqDcs0extsr+0ZluWaAky5okU/dcVxuR3IlNvHntPQvBbfhvS2lqm+F
PIau93P18wrj4SfaG7Ls3T0u8gLvz8tKGeUDD3VtdDbvi6+2edKBuGr2ovTkGBRPCKEPjhrzpKic
2cz5WvPiGj9P+Pgcbm4xVZni7jo+9YWd+IgiE6rLPB42t4ZfoAD3y61UUbMwqsczkWUGJUpY63lU
L7JE187+kwNN5CrUALHGIXX3kHK8ykpyw+sbuIbM7/Fn8GxfljryNe+V/1xsUd08SMPbJ4hEPquB
4UL+PGDFVQMnW/f+C/xeIWlX2P6ahVyHHkE+KolHMQAyreiO3wuTAJLqxOpEs8iNA33jYTLli2iu
ImMeHGq8q29wfbTZdLVI85aDHTajGKr6+bx7cwiqNis0Elq8JAY78hYYR0Zi6IypeD+dEj177sXs
R+9vCpisaz6T3KD6X5+mbwGTktJ2afhaDJSnVhgblfcDKvz5HVoSIlDU0kYk64xX/brzd/chdWhO
u+YmO2hxGzmdphUfX8DO6vQw9uTQ1RF4NcmyYwiSRaJqXcBQqaMLQRsxFUj+mIk9Xv1pnd+lE3sD
wCOVEea9YtP2PnGu7S1DmvlwTKTY2RDjinKI8IutdxF1nahFVWb1v1xv6dAFuTir5bKSl3rCRTun
v+J3BgnSHJwt2th9KQyT83VGuEQnOjtRTh3zWC1uKb/YpBH4yX8EFJ5OSFnxVwRDighSFrD9bkq7
DKw0bqg/JLEu2c63ivGRSGjMhAU0xuvVFELwX3Jqg3DTr4xdpgM8BSVzsYRS/DKxTT0mgwYKE6tH
hcndRgwIfwXTyh+7dcelEfiPp74OZhL+U0npckpd1ZvgpQzjraJqW1XBpSIDNXhGE9k4mnONCmXB
RW7Db26up8a1SwtKCXj/Sejmc4rvNltgwvexML+gDRkWiiLOJy+ykGpRJ/WWmcWU/jMOaRVnKs7I
hxv4ss9Yq+/1FKUawBPmFJMjREcvZisuTaDDOhOEDrrKPgbZUecSouq2eNQpD/UYpMR49mEnOEUx
W0gRtTgpB9ot87cj2MiGsI0yqC+TdWykaq0joU/oM7t77WId9AKbG1wOxgZGgyf+Lg7iSAHCyAsE
VEjnO+Pys52hFK6Ly+pi+JdTIYZaRoxKSI9zceUlhlk9l4hKWJC/mHsbt+AgibEYia0cHSpmG9rs
PXcVUHuMRfSxRP2zC5fyLAKeuDylKJ2Ls2KwQ+jQVv6tB8vakUMjWyVuBX5/OKwH36ZxrRKCdpch
8AopTz0V9AhUBAyisQ++aqxWVAC3DT1y0Jw1KLba8Lg0F+1kOwidVCMia1ET1sSrMvsdX3N5SkiI
1yX3YzKOxHQY20GHZQdibReIhaJ6LtNKJyROSZcqMQgKsGvZmS/WQlDo3ZW9vH527X6TMYLLsvIu
KGc9VmnaXFy4o1mUGcfyGVUC0TPJefm16PF56udF8XJt9f8M6hzHIFMgl87vOipWqEosFg+6kHPx
QKUzbmQbAQMpVjJ5LNrKg9Ys3HD29Dmfxg1kkrtkmq8hE2T7XfWQCUChOAwZtejya1xKC2lxwiuY
Pq2GH+QTkeEpFl8A1QKAsG8MVa0WVLYTXRY5Exp+3f+B7Wqrc3hronGwrO8C3DgzgDtY4cibNBNc
Tdo0bf5cwGApnRf8VFdPbflR009F/++q+g18OOOuo8G67LMFVAXJ4qwMXr9NTT+124pW62V8yvgW
lJZ1o3uDY8N7s0MU2bWqFgf8IgfjqXURD7/A73Gx7wEwIE+VTBE8gTU0wnxFj+/7iswsX08vJ6Ux
tx8VeLh2RExTQv7BgZ/xuheiSNu8GNwTx+bWfSMiqBEeSHFTOcstYdxY8GCjU+XdMDa3FEncBuhy
zFUTGWpqWWcrdjo/hrS4lpND36rRHZ4h4dHzhvcQQMs41qGA0f0JXNouByqDS28ZXb2SA1DkQx22
TGT8rQCe0vEscj2LyF37V4LRvwyeo9X0W9nSRLBQ7mYQx9nuBPGE4+TeEM+Y8S9dRLUbBvq9Yet9
60ul8mF8Bf3dy7R7FEGjY6KZ+KsrDkHYRvxhDF9dt57lcZAUpNuKJu8vQ2ZX7Hkku+KS8XwDxqq5
9Zdm/5bUO0i3FU09KptaK7RAMBdhVXOEu8DtNHW85fvfqmpPeCtuM+WNNpjjn3X0ws1OEdTy9zfL
BSnGYA7QMilwlSnw5bzu15HXfmQOqrBk8/fnjRK5JDpCTi38zDXy3QSXwV5chdKPIluU5kdtTXH0
hnmO+olMvZzlEkVDKCTRUGmnK+ffP1aoEBSRpxTgV7boPXTrqGFjFPqMRIMo0aje/1Etl8hZAfDu
bJc/2HqlzTWHpBqZe7EGvKv2qgONjQzCsd0dsOgs9t7Pgz1UaFzlfKyddB8rOWm40XE7RyHE+srH
CdIwKeAuN5OjCO8HnAoPyR/1S+wB0YdKgYphEp+IQExtYppwCeEmCheLLHesV7Agrl47mDLlbqrR
GDU588XGArdcWswUbRmVUcRLBYypiEv8GF/5nfpPSEGGC447qVBvRajOsV6wXxtNaV5Rsywz6YnB
8MtjC1fcDiw+WUOEiz6nBi/luT8h4wjfq5bgQHGo0AA8Tq+yxom7pN0IU69qBL3eAlz8oib3o2KU
5dfdkMtUn6P3QklOYdOCJjb0M5XMvtIBSnBLkQm/7Ydzqz0m9ub1RysdYza4I1/acd1OwJqd2hWQ
5gDxKR0smfW5b8j2XZFwDIkgS5N0UFLmgM/0oWkqyrWluvRDCv5BPcVuA8tofKDz9ddU4WO569VU
aI2YU9XuhOIDE5JS8FuN3DrD+Q/AGdD+0k0VKzs2jIX3l7mjDuOEMJ0Xj7dB/hoCE72+TQl01YFb
86Ug/Ps71HLBC15EwvJk6UZGcYhIaOR7ROw+5/CcnI7UhFEJzUV5rMyRKxWkDIBeIr/RRCHcerR+
CTwKDVReexBInMzP1PFPdY2bhSi8gXTuEv3rrATkDNlKmj7K2l08l9iyJEhS1hK6sLlJX9LyXmVq
tX8iV0txXZhLN4zIpRdbU08vZ0K2l+IoZ8+u7SBuV3xdqoTTrB7i+PJLldT2Lv+euQr0IZ6lZQJv
pG1mNuoviJNWSWB3PPhGMwA8PZSj+31dRRsX5oUt8+bT2n1JbeaidzLKWLqzaJ8BTZrNetPq1261
sWVUFWFwVNEVGF3V7PVPAgOpwTI2nOzqnj92WaiLgPoGsHxfXyy16gUM/LBaBRzcwZaumOFcGBOS
90snYOtmOFMBrqFpZnPnXMNoz9QJ5tAGsdN9SPThnyOVDZ0IkPN9O/OWuiNVpN85I2Iyn8cLdmZ8
l/XYtjZ4/fkNJGkWCkAL38K1ynms68WZqTox2zBcC/CzhbIxZNYdH7JnyGh2Od1qTA5yn87iRDz3
SPkJJAI4gpoRlw6wzTmw0vDkqxcKc8vBR+yuvlys+bWz1+4/2oPR45yyS2pmDVp8O8NHSX2ojKix
piBQsS13UcXUD1RajrK89B2ncdO48gcefdkTG5aWws80OWUNGJgT0UD6ykm05KcBCNVDoqBivQqn
iAj0fviVPKY2RIYpTcpc66A7DEuKVSNLNaauJBhgONVZFO2kHNJ8sxfAQCih+K6Ln1In0Gk3l8YG
f6lNO854ujt6YID/VfOehpqjL7pAiweetSyr7/f18LiRs/aumnE5yXY6FZ4jXCkXmbJRb9qtqKmk
6JEp8J0desBER8na4pdCa3lfBDs6XxZAT0VvEtxbPQ7VkRLH+P+FtRbNSZcoADNvUv+gErPdgqrW
Vr55Bwvog1zLzu91vHYwY7ZmMzUDZpXQ/Y6oOF/PyA3It3UPxRjzS8vTD1GCcArrcPyfJH2usZfb
zq2wVxj5SubGEROePR63IvJlZgyGy0KJsZaQfCh+2ENUj3JWzhE0fcngqUMNgy8cG6HRnWyswYiL
CQGWwTD4oTCe3C6LQb7m3UjZWQnkpEzOOuwslX79SD6V8zhtYcGEv59L77KuNcL6l6kqoeH0O48g
exbkwQH2pgRqqUjciSABSZLLokaX+62znMz2q4KG6HFL7/oyb/adZvAIYurskb3DevNNK8zCx4lD
m7sXAmQp3Rv1VWRHlTH6bZtoXjgkH7yaT+8suYIGGnHA58CQgIHw05bheohNbSMR4g/j2pTOx3as
MBWxuA959g3LRXpgicfNV0ebc4pyVXt0e1u7qEMfGvzVdw93XOKyeNdkegtyWeEqhewaIPZq7uPT
XoT8AY3YKUyHzq5g4pmW2tnNbU6UzqxMvg/VdZy47W7XbGnJzL+0XDZEZQ7rifa2TgVZTv6zv92c
4hqEIhYRv8THlur9ZRCwl8j81rDwDboCvJQec9tmRxaHmfrk+LbGEwK+zHu8RSO+Rd4nizAtOeE+
ikU24NsGB0SLutgamaJ/UTiCufN+GVfO0hlnX7Nkju5cVfbWsD0DfrKj06GzfoVEb+0Pf/zf5HSh
Vd73xzvbscqQxa+hTN3CoLaHht8o+RTOCzU4u0M1eO30l0yNDiu3DW03FUaVWbdBmuh6gy0AzRZc
dZdf/9WlAOWMO+pth7I5CSn0ff5poRfqlKQJOVLQQ5qSl0tKmXQPiZKbQsP7TSMKgMWo6NwQroMd
x5rwwDitxhg/xbHxRyx0aG4JDqLyS/IRXxH12vO06G6/ruRSOiBzOIreO60XZYVeMLFTYTH9YfoA
WRPSZVOILaV1pDlVT/H1xQKrdkN7P6L9fJt9cXrfLkmRyd/m/jndtPnHxQj5VhQPcnzvCBnM3VIp
MA7xdV7EW8SUgnn3t7YCuvVNRLEJxyQwmU9vDFDv+fFtYIMHa9wP1MzK+n6nBXv4D2DonPXlYUg1
YxVwJKmXPAmxN00zlSXUzNpfGFGs8JMbbsAZZ+URrfOMcLHgiQXN+TVqrFJLLXQi11NCrbdxZ5yg
u/RQoJKXmekcQ+YLOBFQAA5pEUNV/qGDUuWO9fldiXWFjMB/AeRQG6Rq4E54IZgYHp36oysaKEfY
HchWzfA8kr06SIzvis7wxeLm4kgQC42/cYn8qieZIHgtMEW+kmLb8wHZvG5O3TcpIWmfvp1MI00F
GQEmFOmB+Fa27d5maqc5E+76X9P5gJNEhWpC2k++3AwiuiE+lmONoVePuN1g6KAs4NIcR/J6C64s
h10vZHu8yexur0F9RNh/bd/AasGcaVArQtSj1QRnRI9nZe7gzF0c+rK+KYpJqN80QpMvyTtrWsmh
pvkSuClzfQq3MWJSyIhRRTO9GkwjckPUNAui8+P3O72XdGXWCuRKN0f5fmM59jpmXnftYZzskcdd
D1bSHD/eF2MbpbqUOAa1iA/Z/gYhVMb2Ds5XNkYE3g7e2ofIL41yU3yrrqqkjFxozHZF15l2zKx3
hhtu2hGubEN+Vty04GbqUBeGWhZVix2YyoG9n7fOpC8A+KJllXtpaQ8dtTuQ/IQPL7r4WTwUGgQ+
YVFXOSyLQtKTY26jZy19YkH9p5DAGyE3AvVIQTo3jPNxkaDiOwKJuLjF0CYe2ef2K2+yfQHU92uI
fNoWNhBd5ORpnFslL+i2kyAHW4q8cnI9pBtqIxcgmEhr4+jtG9ZxTF5D4I0SCSpv3FlPt81cw4hH
jvAyT58g8XHu9qlDUkbizLzby7fBLqgEiALU28eII0sDV3i6u2oBdfm01qM+eMNq13AYGN3ec1o1
VYsab5qYF1MUFjghds98+6lv6CwJmJXh/ZHlRAbUoSBFwpH6xmAtAUcFq4djedi7wPsYXZd71hzw
hvQyWHYqegXtzMcOSn3zY+ZR6gsCqXSjj++MxB/8ATC8P2XKy/SNzOVPZXso24aXI0IXAmT5b/V2
8v9UmUcLK2HCS2PnPkdvMZaV3LQtpvPCbO7qXo8Zkv4RzfHx7RTV0Rv/9r89AOxbdofNUq9r7iKt
cf2/5a2z0DDkNAh0n/JYGFedBxYcwCM4AAs02fSq68dJx1mYzdwFGKsvTzc31Z+ZrWfyDv2QFZs4
TRwfQSON2z/99u6BriJYy0c0EXYs1FnJykfMaEp/TwRil9ajo/TBQaNMN0UsB23Taoa22egYo0d2
SVREi3MZ6m0VSEWJ5muwVYagh7KclPUrJImSa2ribxp+YjPfRUU2ez99nX3tF3cNnaj0EZIdfsDD
BNPErzoXEeN2JKyV2Z6HDe92kZQcTrupcYv9WMRp8/VnBzAHuAXkxPBQMf3k34v/gwfpBKVHTJsS
nxvQmISnbXmvU2lFAFpxzQS+mMDNGOf2WQKMHmtUIHfy5H9kudVWU6sL1Vmy8ipRFgetQ5wMAa6+
82PjWecONf7/ojVHqX6SawHD9xORL1iI7wydQS4tWIAL+7ZhHkhFXnWqVMHcA2pIG5NQ7pA3Vfii
XthIP8ENI/qw/fKtsnb1DEksDQjMcHnXFjsi9MxZo2a7fJvevxzB71nzcmLmUib2LDPY+iP1DJXF
9aMpX45uuyu/QASPJhIPEgKz+vAfmUUTA8rt75ya3/KN8NcsTvCK+BFJB2IcImOZnxQVcTVCLsbJ
8DRSOwZY8W9htiUMI3bdLRpYZUGv1N1lBNkuWf5AlDGPkNmAQQclR0U+S6xp2SbxldINh50v/aPU
iV18ChwITEVemdS0ypNkLthe/AGf4mo/WLJGA0qv961JTZNoNvXC5arRFBKQcuPjARbGeohHC6WN
E6yhfNDDj2i9nicha3UgQDSQ1kzzsdLPVed+5RnnxtL3d9wjg5OyUteuefi2eKA9UxD8zk3LQmqa
U+wQYeRlEq/WFlp5PA6YDBFbd7bhu37C6VRo1rQFx5If/B75HWVi3IAXo2Z2Cko2JQd0ZiEbEPvj
LuorYPrcSr/9FKVZJraVd0d91gcCTKN6SHyNYxCeMlgxnkFBK6IBiMLXGlz94eEGWTwu0de/8aWb
ZGycqwEJt+VRwd/LNJz7y0YfLmYcgUqYvsPEI+3nQEHfda+iRudYR9no7k/EJOdNpvxOxoI7x3mz
WVMgI1tyrOKuQyW1gWCwssoBDG6Si1cawFb1TNuBzMf4mhBjimnk+Qss57j8CEHhV+Pd6I+hZmLm
nOqS4zMfMD/0Gl7I4+wUc0+LUjPMZs5qlIsHCX9BGbF1lUBYSbB1joM+r0jEurwd7KylhlvqCKRI
sP50WUuZ5vUhNN9qwNsscvM7vQ9kFiJk0N854EbBnRhiIHDw/IB5VoeQrgj5Z6rGr+p/6LRlYhGZ
XBrRL4hjtBBrdth8fohnVl2xRjBIxfGoQq05ajVMGWiMnIdASoJ6/0oF81U+5kwKAeQGBjiTLIfa
Rpo3C/4aNDL/oy49c0UHyTTnKQkTC5PwlOW6j/3pOGUHfU3gTBjWe5l0BqDLGZPwCYt09i26FEnq
e8ehb4Cf4pXmSQt1gZzo72vsSmt9sld+UJ45nEpkyYM9DW+LUy8mWqSat8DHdCz17u6OmVXB0pIE
/+zt2nkMN26JTbAtwBtCjQ39207POC2DYgC6ajQggrEB2r1++fceQVIHKSNsax310obrAHMjEZLm
jKiktDpxbrhAH5WORzDaxBhaxuuOON2JjDCBcaXy5WwGadESYU8xxeweCcihy9byOK7SlHQea/t5
dBbcbQbj/kccZEkxaftRMYFdRi0JVfdxZV7Ged1Zj6EYcYP6Tpj6kf5O/EcmiFRqhU8pETYLtHjc
t4sSUNHnl7O8yz6G81+Pjgxhbegh6YTqs+u7UuezdhxSqURWVxDfGd70+L2sOU4WdyekbA755JC5
ow125XlSGwAHsjUnlOeYTLQkPVzGOxnlotmog7MQ6k4CLnxTaNEOWSHNhd37BDAkNqPa2gX32bok
iJTFuFeKqvThv83i6JiLT4FAr9baqQafwv6zQqsThQmeLFXirW3ySsoDKQjvQV4t25PyBMjGeyyd
H97OKQOKSOq4RH2O00M3r7c+f72Lioqcyk7w1pkt0Ho6FoLVOeW9TKod8ys6et5m0NT41/PZZ379
kCN8uWP3YIGtTee3gboPIYQaXfUk8UnLpp55FsSjmTilxH83gYsoa/KE/dt3wTWSNwGJI6SXZMK/
AKCUARyWO3HyeQ81njgmNciEVDYcWOTnYhGiMwk5PO8yoVo0Hnrk1FLwpoehlvb9lQvvw+sWJQjl
YmL0+Utyz7td6Fg5m7aEFQ2LsDnFcYm0kDpH1rjM4dXBniiMOBDCjrD2RLr8YJV5CvTMbTmLengH
lt97vOmxkiB7iTrlWZDqmfiTCOLEquVU45/bCmI2IZq3+wHh4PdR1XPzTgsJ/tij08zHEfjC1Z+8
KbR5kO0cjuGC+14J3UQSVKIAA6Nn7aKB443AIyxcg6a9WRTKZ8QFvnJsgB+cb12B5WKE4msAUMAB
0IZKVwoSfbZhsAhBS+WBRriFelAtK1LoP19ENSMZAsWGw4rcWs3UTwqCpZy/R0hiqUBknSjx0Ke/
StNXI4gfAgPnByCg4l5TAFjxDKxQAUh4BqtcAZg02MUUBomML1ieD6EYPtHJJ2345coU5cIYB/rx
NoLTqnOur90F4TuYCeHAsaC+PE3XgoaSGirYXOeJrTgHntA0V9m0h+tJBkgK7OsNqqYgSwF7jGFv
GYlivKhSypQn5o88p0J2FRSGBjbnPG7591Eif5QUx4NWN4IUY6u/oTlTcU3paf06gG4qdnRkquts
Px6fMY0u3SzE1XTktufzsYkt5zRX1YxeYuQNSJuDs+2FuzjeEGvySKTSP7isQvHh+/TPZu1S97Rs
gWd7k+OY9tseB1qiUpHTGRnZFrJSU+l6kJ7CqfO+yTNzy0HnzFYQ3UBbtyqEv6c2wHTGi+DwKThZ
nRIUY8JM+MbxJe+KjTCzrMerHjaBEqHPH3EL0CpZrGxeuYWaDQUbDp8LwCmsogB/8+QlVGQrpFNh
fsbxS5P7tfTvlsM38lnboa7lfOwVZTdTYYiJA7rABraIAMo0b0hUWSp55p+0BYDLUzfAq37Cg4fX
2tpG/X1teVcZ8sz9Y2VqZRLaMXyVzFbx1WhPxfqgdYQqcFdBBaQwSW+F7YjKjPt1tosUJ3xQCNsJ
YvjJwwbWeX0uHP5rwEWya04pNCrn27pGEg/c0L5hDzAD5nrqEsG8y0Sh9P1oHoCPpX66aDc+HNon
OLXKoq/1SB0UdWfQJVC/lZkShInTm7qM9gQxKxXWuTeQihMYjcMDpMDRJvtb/VabVfeB3Tq7rKha
hJ826xQmG0n9tM2rMYVRJY+6phlWsq1KTaeGwnBhpx4fBarGPeS6qo4DSto2STGw74wOsSw9nHRV
cvwj+dQhZOYCcJWoeTUSQdW3ilch3F4Mo8hgI3gJyUnpkQjMFmt2JlQ0yjYyZLongVPkxIFZ51tH
3+M32/HlfKOArze9t+HEJMJPKNHj+OdTLkV7p/O+7TVb7NqOAoIiBQDL0DxE3i8u1kUr6nAFy852
PJE5WSldSdGIxlAmgyye0IQKf3x4IvbKi0PcdhPJBtSpHosB1T6VeD/d5ByAp8c/3Ygquq5jR1VE
Eo+4AQlfOEVf/+nckW51EO/zfQGosAcNKA0lgzRSlWQKQKOsQcV5tJc+bwrsLhKkM17/Eqn6bjtj
oFxvI5u0ZtmK6y1mkNvQvfyE6G6QtJ/Rd6fI6dWu3ftwo39tr/4kIX40Xsn9HMObF3QPniHoNIiB
U0SW91heK3pCLWkZhwV1yoB7n4XROLcnTyLpS2WcOpfQjw56DZRxqoAdT9L0RqY0uuoPTRItNUkY
tJmot/U6XpsmtOA+TJMFLgmXjUteZLJ4S74NHgyuu4MnTguf3w6t/XnMZgRvY0Vn6kgs0vVovkj+
JjSYMAoJQaKpJw4fl1FyvcoxCEpDcgf04pgIu2GD+C1RmouIZPVh9d7rTMWIARxoN9BZ3Kevurjm
P7Z4o+0QRAFBcjbObi7q7oTfU2FYnW3DO9o03cbMdwa2yBFHxJzvj8bWB3ItVEHeP2kadcwjqawk
pBhQjJlTZRf5JzkwiDR8M4frl0/VFvM0mvCDTPTMlODOEzx3H4re3ysNwzX6+zWL0CjwUe4hlz7j
fIJ/FTLl6bzlDFmLo7+KUM4nSNQhPdfLEBvEYnOfc80vHLKjtJRgrsxq3IO1yO/uIIcIRg88o2h4
Q9zCOd9EVZc8NgWMM+EZuLgJtzjDUAOjD97YhaIJncevUzFxOQ56xnsQBXc0wayFNIdpJPdQXPDS
cYvoBuV+9VbghPwBJXwEyvlLvLiqDLF7lDs9qtIHUJ5tiJfvJsl0mAoUK+aeZwr/mYn1rU9N8uwj
x3hyKB+dPP/7vj2OGytjfcEE4JNN4AbkKEOhIkj7GL2itykGBhG/jc9EC/JwN8mhfxhfQkySiArQ
cDZ+x5T/1zyAdBZvqiJKGcJjiB5AADc1vQ/vaw0Szubd5bBp5SdJcb0S27UTjFb9V5er1Mj6S0U/
hbkOgUkYAp8psEuO+BAomFatD5zLwyMcqxg1JU0sMuErFILJF5ulgW6kX74ZVWXhyWUZ4r8/wiYX
x6qXjbegZrXVyj2wXealBngoaKlqX4MRrwRaKXUv1XmQYXk7UD8wfG7CQwT00jPEQ7d49hyj3XEf
UJOVjDx8kSzAu9MQ8WuK4VLkHlzL46tKRact6xll0XuscHBjaLUNQ4l9ZVE+Y/RdcxjRzxwEBkqT
EmDGaWTwMyZRxqWFThVHe2c/gU3ppCanrGsZ8SH1DyHGW7M5W+SFJflAFIZHzB3mOvNen9sZ7RHm
9+or/x+lpPEQLjx5g8UDuuigPL6Y/bNtmUr+iZT0gJVYuIBFPsQgJU0vEECKhzohWPcl5AK3kjgc
gQynF2b6dOSvKbHjVU/6l/v3TbfqcMmw/lWAt0c8yKCQFwX8kCrTpyqp3Q3URfzFvwZaqU23hWG3
E4kEvm3s0fVp9la1ybVxtk5DauM9Bqevv0TPbQ7KMwydLW6DcdwoZdNs6ZDSqSMBTEbDuW4izpgh
GGuGgdRilshG2wNvg9TFNg2xC3Egq5cU9SIv777he2NkQYEYkW1C43V2oG4dkPII2dSRTyv+xQtQ
vfW0m6+T6LmWhN5UaKtoVrWGh33TOa3qfQ+2nSdbDq7yWor9je7QS3iD85e+636WLhd6PgTiAiwa
gQo70/HeQdbACks9AU93d0gx6IPmTDVzB0e2uhL8gZAQKcs2xr4u/rfRpKzDRm/RxtfYH/oVVV2x
FvUb/HOy4amrfQCpUm1jkA9zrO12EjkHmxs4KW98Wd8cJy7BWcUkJJcn6pxG+GCCqAa2uL1ZYIyj
y4JpjsQmHsPDiiVmqptnUSS7ItqYCTT+j2MzhazJL8FCNEUhAXZztSNPRWUcZG5VbDZUgUDD+tb4
G8MLVsKV70EFzs4+/+aw7IBvIoJXaFH1qyw3jwse2m0OORTsl+k1JxVEY310IgBkriN/cofX035H
k24iRw4VQYaYNQLKDqCeYed0G9sqH+WNd8gTo0mhU7QGq8EYzo8HwgrJseXzRgPPReg6a8qg2iKg
aCvxUk/SjDdT2VgdY/nNBVEZCbV9CCD/wuVqdwzZHP2/XVBSLvM1fOE0WlLDf0ixaSkKi8Q27NVB
2ehbcIgRGcoJDsRUG/n3srbJBP9f1LP+Lwuo8Q/IUsByY5jMvviDh4d9JiB4Z1mpd5jSLYhyT0Ja
uKvwFRumVao9slIK8xx/8zdQ6/mbvr/uVMXsqcdJLDQHLvt+FOvgvxiXqrvWq92kFWpnwwvlGwfZ
XjEY+t3KOwojZXp2mMMzC21ZgVAzgZdipJ0XDaXq3jlsWqIoZz0Mq7D0b55H5LyWMAWGsjQux8Zc
KmwpWDZI2BThCPw8iVIZ5KOpaFCDWc+MVNjqiVkrx1h7FHYmY4TweGnPHlzBQu1GDWocHOqBVqq/
Ftd9q+J0360GdjNieQykkAT+Tb0uNrgtx7GOL9QCr/KiJFFy/FoWJ4dXSuutd75FfNUe9iIBhl3C
RGKnlrgUyR5aq34t3jMWKLyPs5eX85vXj+fQG+GFavnuDtRWVLDnmCowX4cNx3uBLgGJEnf4in38
7rwikWOfdDacN/Z1ynJ0wtx4vvgXk3Sx+CBMBYBuDPQxWF3CIltuY3JeJuCwUKd1Z56ueObtSN1O
g+2JyAxn4r+NV2p95jzi7TaEnWrZY3kQqnkaZlsKBF51nb28LAp6G9w57jHWRiGz83ZiV9kyolol
cusMrjD/lJr5GcK+AfTxieTBsLFhu9PSV0NLhB12KFj47meg5ooKa5lAAcb2Kaab9MuDrgukn6fl
6dHyv2ZrfTaaOjAAj6B1WTIisLKdLvCko2Z8/5qAY9v7CNwQBssJQlovISkS9vqOBQW5ZqjmX6dF
IxMAIqc9ca6je1Gx0mai46oOPQ7hFFdB5+/Zlvm+/OTB8oLV8QRfOvKEIrwnzUaPzDcPsx5tYcBF
4OPmDEimPab/uRRW8AO31xCFwJ5PiESJpm/7gqBRKPXNMLgKXFBgz0I1PxKRIc5ST/EQIl7D4cuQ
BEbpjUHMyisFbIV+55Lz5iTrwF2SMb3qtc4Bam1nbncB16JAB1peWWt0Yhf5BPYIxrADUjBIKg8O
Wdla9d56o/f9QgQ0HoM0L2RW8LE3ZlSiAM1ACYn5sPDSs/VIgK59Ma0P1pb+F2t8QI5AhBjJbUFR
poxhvIfhbGeXuzNxCMPENMLXr53N5gRHKmgoK1EupsH+N+6mWMQU+bbJ9Jl0asxrq5EGbg9AMf0A
T789wM8uyUsTkcbxVLTI5HqCjDWmTrmfxbMy9T1cuaz1MkHwPZByQ+D1d9/5/B0PxedDheWtAkU9
0Uh5jT7JI+q0nfzpTbOoQRENUceo/nBbXGs6uA/gkvVybPDRxgZ8GNkah33QqjTUTsLJnIGbfcds
bKHsgW9MJLfaap2y8Mi/n4dcBeYeO0ZTXRXsXH1Fd5NjJ+laHiwMF2GC3YME3/FVskPpYZzmw0Gh
ihu4E0e3RqeT7AwukCtnIAit/GnfIDSTLWP52VpCtl6SlLb5U4aa6f9cC6g0h8oMKTBpU5Ieovar
UTiJ2mejr26FMytFCm3ordSDWMuGZzGLC3i0lTN2PYi9fWaKZRLwrcPQf/EmE9HEzPjDw0r6jGoc
GfAFaYz7xkkY7SNJLvtO04EnMIxSYh+BlIAp2+4mvg1EBMomYsSWBZQNDrBpV+sIvgg9QvOK8AjM
7TlkMo4tYOsu9ecRU+ycJtS7KpFdyR0uq3RP1WewESz2XN3cBShpcXKDBN9h9ylydZeIZuLlIytu
mteWXxq7pN0IIxTHP5E5Uotcjb6EsvYNrZqodylerG89zvuhYh5oC0G8sdBAXP3Z+Le62FOXFdu0
Cg9EYByUO4pB2k7TcCRtRsO5CDuBwvKVB/CKadLXjZr/+P2MVRhhYdI6UGURAGswQW8/aYi5V08v
3Vs0THJQjTZHcOAX4qq8FWxbDR/otMm4XSyESlMFYyGr260y86GfsH62c/acPP7vQK/4J7nZ8RtF
rkrXqaoMJ0+1TeOAfCj7PDygGoRN98y7TuSmBm6SP+e4Xxzp+hoU8piQ5HbE5ZpqXunsBYtGljcV
WFj+mJM7xTBxuoJUedU0rRodfQuDMRmmKkaSEbcuXI14Ngl7NW3t85GJGZjKc3Jsrjn9OYQXTdcC
IDiRkdN5vhuKL5o42mbJl0Scp3Y4gkQbfXpaSTwwymiOgA602hVEOouwdD+EdctTeFBBfZsEdX/U
XNce59T/RzmBj1BB6qVQZsonnqVn+w1XFvWzJkZjYiBtDEEZcIwJSKtJbA0fZKhA7XbAIY6Y4Dll
EnXOAGvLcx4gW8BlIW03KWBF5KlWqyu515LHE0XF5TCqvnF9wM2tA7gtiPI4t7Teus983YN6hotd
7fXGf7GxmHXE5Zw3Nkso1toQgz2Q0gYPc+irpEMlM81IoSAT51sop/C0cUhRNsRztIzZOWXRkrjU
IOF+XGNWznSYHc25YQTlqwNhu+UjF+5xy88NXC41LvXJXZ/V3kNU3j6wwlCxsRVw4GK6U3dqDIE7
bVR85xV1C8EL20ZmfgmxxzUtrWoyW6jfALpRRyH4fmI1kFBHsBnbJFpuzqNAu+hpm3qCOb7x9+4C
vlNbNAw+RKf2TUU+abJo6WaxbhU3olWFBvb3Om0TKuVY9AYlZhkW+Ign+AwsiCHWU/e30BV/N2m5
yi21AmjwyXSiGICvWudrVauSNgt7kWAxzIx6FxOZ6puZ8pV9luxlIYkIXEry5uaD4ZcBjgo92mXd
IEhIS5r1YGUFq1H2Wg5JIJM8UcPxh75OgOeF1gHTXXhb7VlF0ab1pMJ1W6g7gQ1iHrlh0HU7GBBV
7vlBFEXtW/FCP71kcCWN5Ykff1ibLwv/KaQFhdMoKf7Rh4ipWf2ZGObMnrZDcgDgybmOkkGfsq2k
VFdajczw2lxji+dnALI2hNxBq236mpnvY96Um4I+fY4pHmON4YUzqBJOc+zLOTCqvf8xy5AgHq6D
NtIqsF23a5yvfQJ2IW6La7v1/FL4lI1+O5uDUO11SJTLhbqkuXWRt8sQP3ikVjXQMxiarfAOJ3QB
Mn2eZoIHzyBfeLkVVwBXOq/BSfrGYnB5p50moYe+TZonED6AjR+bIwytc7o6uTVIuh0MLCw9ypfb
6ephFk7LOntIW1dFcMbwZZT5PvuWuZUvAsCIz5fMEHnLDKrsehzuesi+u9N76trOnmq+/j+jQFij
kq0ZUl3hxm4wnTctLVPV4jlA3Rff+OBrYHGcL401DHfoc7/ajXFAXf8y0B27PTp8r4RSfvzZTcE9
k7MnylR0ZVdadSgvLEl7PCpgqxUWi2ZA+Bva5zLm0r7v/NEAF+DLifuCTghx/5IiSm9SekwZSXCx
BhujQFu++5r5gMTes5kvTtMQGBv6cIh74ow+Q5/YiUfnoR01RYFcuCupimcuw8OMLYaBquI2+x1O
oEmzKevrAgLlaAmNJLeU6VQhOeIIC9MMouhQ7B080AlHL/jyo02dmMdjdGszp1Exhlj8pJdvDryS
jiN4+P99F76klsmuK2NS1ip0T815oV2wr+0TBoeUBzlxygHQDRTMCxh0kunyM8X99jpyq72xqiMt
s9iMxWt6PQC5oQ3ZMI9HzyIz3nGZMyDgyZnLrfrfnk8+LQjX3PYfQsM6on5oIiulNqXPx/+Cpo/y
RL2p40LH9cfiH6/4c4LwCOfgaBGAbMnji7wEJ2d9b01cB2O0c6p4ngygi2IKB0S11NQPh9QPGbdg
3bfF52+lRLwPni66cU7nMO5tvnZbpHlBdE9/MXSNete1xmBmSidD02WwjqECmG+B9ryC5gnN1mdJ
Yqxmf7/ASOyqte3lc07oyeYo80ZAXw1dLnFvRVnQ+cSlirBKs/dcOTj0ovn0yW/OGrNiCa/T7K28
FyVK/l+G1pS5EzgJfrFoYMEpXppdLgfczew4uVB4LE0t9sLHxOjLB5vEvoJ/u81lvtm8memftKVd
mXuOmjZhsxScFLAjUWXmdfNtH2vRKbshPlaXMtu0X3JLPz4skS8D1cKy9cMgrXYbYZuysDwAg/NG
7txi1xXwQU1QsrpJtGHicC3h6+nxKB+2CaoSr5jQJbZr/KatQatAvwKAY8glD+yAMs4LeY88lH5H
RQW4JCFkflUgP9EN8AT47wCKm0dQnzm18tGa/9Afcy4srF1oHY8FKId/F3UKszJzxbJ0oQt4HcHH
vqr4wEbXWuLGVhFAlqviJ1GcuINpQBcbJ3OYQPvSzuV3wixk9N1j+TkdbvrdoO2adCxVP7A7giWs
nRvE1P2yWseP+Nxwf7fYvFS6P4LzSSIEgHlbUSvV+5Wl/+E7Kxm/3R1fJTd4qw79Py0IUcO+egqi
tC9h/22zP5GFX5RCy8lgI2PPlNFp8aMN6wjXxPw6I+4zSSI4xzBMC2Yd9mSBAyyjcVpOrndOQ+XQ
gSyE2kdLw2DmCe8Lqcdq3JdQRGhfwuKNmqvEvTn9YRioyzyygvgCF+U4XLYhPjwfDPwjTueWqPoE
bgB5wZvycfDzbxmV6lToV8pfuKHHcFeM36Bz803mojAD3aC5wl3Z3NjMM/rDF7ceub4uTUlTRC/e
UrqPkb32tET5njvcVhAPjDrY1j8WS7HeKBG3iQsZi13cZjfDOd+FnK71/N1iao28nR29LFKJ/ZBB
27QzDr0hf2OcdrIM9OBDRrFvcgOwNsJ86BkMk1p1ka/sABXrZ2y/tvTZd42jcOm/zGKkeXvx65JQ
eaN2ah0iK0rMFEf0KE0hGpKPloE1Ib8yeSdgR36LGkFSinTaoYAtVcW0MUmTDW2QJxarspLKBqD+
0XzGh2iRqrQFR2CoeNv3hPV6vmxqe0gf1JamnEY8bJKNTBVRF9Gb486autz0KKx4+0f6jsnsCgj3
jpYS3gQsQnprkmHbsf1TzD7feRobiZLQdU/RJih4eMhamsaIKxJkGt017oi3aq+A9iMGH4nM/BLj
n/a/Ys9BIBm0m6SlvygSe+tPufaY+MUKvtXfT4ouCs3zO8Ek9v6JOS93fYkQ9OjhMULWRwOiqH4k
GyuMlUvJzAV9TTHcwZLNDBQyxvpjTeKmSOHyK6MMoCH07LDejAhjg5S9paF0tm3SDtzIiV12kuZc
r3A85wGyhq8pu9alblzWxNug2YZHN9+Ecm4kM9NzR2pEPNx24dIFGrN2zt0RmcMDXqULUzxcaumB
8nEOzP26OMrvuVgsqysNXDb/c+ZzNg+YWv24XJidro49uYLWxhhbEuE3hpDf2bl4czVIU12yO+vx
I0Yp99s7HU6GvNQruhrIRNR2TOj/RqHHdPsL6iCKNSlIpRXmyg++//caEJr6wtkh466SL+FxLEs9
7gbD2zrQH6AAJ2cqk0IbHgMiUOmilNQF1ItvFzBa8vG99F7Guib5+cXPla9r2s9yMz0C4b7+o4un
KYM+bgt463+zduN306Y2ABt4IXCbs91CRrwVqCQuMZzneuFZPhfLRDz36MTbRNx2McPMSPzeP34m
AwausewdfTUN07N4+HLheQo+r3ei1Q4eFUAbyiTzKUiEZmYULOIq0UeOMVZWYemxqdx1wKvrLyW8
92XT9zrY9RYmjIoAKbLSUCk8tBaorYEceRc5G0sNsLeMmReQ8swKT9tz1FOFTYkce7kfxDyoVieB
hPqy6yuFa5a/qMY66ne7BfpowijFrkURcTAAdLH2iErnn8n5JyZMty65tEgMMvlVoXcyB7y1iuKe
+2qxo6fyalKgQRN40kp+lLhigFnJIu7q9mYDLclaRgqBlXaEnhuONRUguqriAlAUcG9wnwFSh1Bf
IATxhsmaJM3ePZkONbCDh7lhP9/X8BZbP6yMgptuiBFMPoRD5pVkLoQUYtVHAca04MfD+A4+CpUx
PyKnlbY9aYZfRB9xy1uAn4nMz8Aks7a8l3E/BKmgpgcifTOGY/j+DxYoWtMV62/oD8UOCx+0S4IV
Aj3I7WtuCvmCKJqHkbc6DF+Udixt9tYjFptXZxQX5oGH9nKHJ9+NUW9fFJuVLyRiwIgcKQqXlbq8
+sWGmBNOrL/uHFs065Pk8F53SqpRXtqSuveni82rw2ZVd+jGTBQWogJlx+TBm39cI7vyA40p/+En
bFLR+IF+n/tmILgjdZnyGH49zUGj2B0fTD+tR0Go+UXOKJ+I70WcNUtbU/n06j5LUxs0bNcoRbNo
TFHTe8JMwyWvob7T+nCJr1lwNB8Ht9Dc6URY4rxVmxo/FJuRo0bm4sBrn32C7KCWK2narLPpGa5N
PWnQt6WLsLFEDltrbyMRqDK2f8NZJrw70I11HyV35YO5PLjA28E0hvD4MzEGKY+EMeTp97kAndBG
T/uSAuFphn/3MUHhzXbAmMWizxTcGkFYCKUaNvcxc9pABQhVgK9XsEohEc0+RKv2YHG0L48NpdkL
u4EwLd2pfLRMuSgkhFOQQQvT8GvotBCOkJJ7pNKw1D7M+9cMk4cli6Jra5os+CztVYvJ3E1hpP68
qVSIxDI37WQ3MAOIbJGY4mkovhPip/fH0UOIN1e54KvJC+EmGu4D1g/eoTmQ3jEUk/zNhYORNt2+
4LxDdqjKgWPu+wtMaGfhLkjrL8XyiiHBuDFMNWUbxFcQO0gMM39zjEGEOW5s8zGzaWS7KeSca+ky
YXTOnsbzW5AadXjwSwgEU3TrM7rp0VQNxii5UzYoPDRqU8cb37O0A7hE2/o39whzNMmdV0yVMOeN
HnvRmayB8nIqpJzTSywdlcccBpkUojDK+03vXVEPw/Qz0HK45mqCh1ZGJ2/sjRMLMJuFDKMQiQC8
ACZUDpduBiDvhyDZFvS+VkQxCii56NBRv7GATnb0o07qWy1upEsHuf5Qea2AA2Kmr8RYkGCpbU+L
Kgv1rmkXB87A2CcFcVm4g86u+VdiaI4669dGLG0s4bmH93dkk8FgdcjGpeGz81teU2VRGxJx+7GY
ky3TCLqfjCwODvYbO/0gIpnctgRpv7mCquAQqJ9+gzisRgp/bw7vkSkwbNRxh8hPj20OyHYzGs1V
7SVHH6yUZe384ejdJ9XgX5gJek8SP/DrVqe9CyiiYyjFd+iw/OuZvcBL1ujLKUfknGC6q2dvzNKT
MSeeW+38xuUo9i02pIANOdw+W1T0EpzpuroWOOCfGvShOeXcApy973szuJsav7TTN1sJHkQap5I+
MD7IRoU/HQDzEnd5AhFIAzOwxe1PRgmcAFD5Rg0q4Irjxsz7jxZoL3aStV+3wlvNwk8SsWHkP4Sj
/LmHB+koT1lvaF+z/bT2BmAFe3PB5Qvb02ljH+0XSTcBWxNbVSBWXpH/rrUqNj6kTkqT0BF8/hcv
8NKKYBG+9J6Spvrs8zJKzdv8cy1RrRd1aFuU+83HHnKXr9C1dn890VClQUQHLYyk5V3vtsmCrrBG
nVJjuj9utC1/+3p1A0bcrTxdyzU0j3qfACTcsq03bjA5zbrJejCJ7Yo8yyP0xApGWlfHa23npsDY
L5e5OqPUa899Y6pTWFzrdE04hNRoongkfqnQM6epmzN54oqPa2H9ORpAOyXw3mSF8QT+wH8iEVto
Mkgp80oKqAeB/98cKPyMVS5lKdtTal8RxHlW6TQ6sYUKMPzwsjoq6a1NfKUAxiroB1oFKT1mbfPh
ebTB2LjPi6bpujLtszk5sSvfXuo75/cU6OOcmG5t/0RHFYmroMG3TvvvoHxV4/7qTxKu7Nhwfmvo
T8pc9LZF/qaZFlQzcHcpMLb6F4qIvPgLvd7DM1MJdDxH5J0y4u61q4vpoUZEN8JZNZE6rOTChV1W
EbPuPQcF7By6SUEZX5LCYTSSF96yPQfzhQMAB/adw3i58UqFsOqK5QguEJmsyjjBk6T4Dz20dU/8
N2XII9TU1gxPOspkJUfzkA5jHvzsHf4BrkvPahk5AnfLsLMNHLXg4JV0JF8abdN85ItrKxZyZd4r
O1+WkeBEAqMOicQTDWDmYHOMZHLIiYVGazjXd2xNIUc/iT4orrkFaRmtmeLOIXWpc2ufrB04JZB9
ZlMuCJ8oweSxOF8TIFAvLlRdOpFpWo4EKuZS19wUoMG+gdaTvVrW6KP/Sp1SZs0iky/2JW1/IGid
AcAlODwg3Bs1YUpjqZRz5zUOHFyzwL6iOqTBZEL5KkbLX/Ofg5uSSvGjYV0YaG2hMIeAY+MinAsQ
gc23j+h7v8WLM3gzafVcv+5KW51KTxcd2HAbPkzJ48xck1V4vfGb7L0KKSf9r/DyOamXhfokahbo
WwmEFsYouwklJIdvNR/ig8NfOCv+uv9VL5h83/2jF/IwpjQoDAdcBKtg/hE1eW3vgca+oR8j1fDE
+zUF+5UzFpDTH2MgPpDtUEYhtwNOdxllQoQMk7kKSOnrxytK5tIR8pJ43jQ/t5Bnw6Q8Hk0OhT+6
2/OvkqLgDQ2K4fbkTvNKIx0odTYHMqM32eWU4/EoDnrHO/J1sGrHcxoS9yM5cFHYragFvdpA2RG4
R7ykcpL7Vwtv9XO/jqUrjftgalvZbYdS7NFC0UVpOCBHV6QtJGW3Q5RiGnnyU42PjFsSzZsyT11J
i+Ftf1zo20gDOMH+5S0G3NtVUwKVJ/jBGmK9Y+Ox5xRY0FGFpN28H3Oi5e3sUNIjhEjbkj0Krmzf
bnyIIT2nsKTAaHhmothCISj0eQ/4UgPQvJcIbOLIL/qxvmKk8lA85lU5OQI9hmsxqkZRqquqj/Af
T6nhYb1lRk+V41DIwPPPLrOfy+sCXDBx6BQtH5iqJy2uhqVxMKmjZZoQjnC0MHCeZmLvZHa2nERJ
p/0yJMiFFKtDaNdsBVfu0tRl/U/H1uyavz49yNOwpqpd709YwcN1yOZE7k9AVih6x+Z/SYN0QAHC
2ovJ95JXI1MyCADocb/8x1QzzxZAw0B2gp7dEC+Z3S/nXGlvVSZsoPWrX28C+WDGtH8+vFO/ToA2
snaw2ukK62NiiV1SrhAxCnyzdDocmTxBJxRdNij5AxRrH6AhuRlCACENK9HMkeps0JHCFgSXWnd1
GKA/sHjQkj6GbUcxnDFxaZ5YX93rwcWmxrpXNwRF78p4MaDyjgtJ4ymkrOMHBZ0VwNZ36oaFVKAI
Y21MQK9UKInf4wBFMvt2AExkFpmtB8BISydAvjkZvLbod6qgbGwpe0NtgXgDVWIDdgJbt1sCem1W
L3U/1+6/SwtWxtru0UrT1WZg/cDVANf9BjYItUaHer/ongvsiCuxBMa8Oz5pw/L/y3TH7gj1BmxA
bi34Wwp1eiMUf68HtBRALWRg6/ID2xGUge4I199SoQXcTlQP/sK3PdeBFPxbRMzRwIn0OEpEaVDY
nz8G3y0KIMpemYYFv/Ca1FwYSKd2YLk2hLoixZFIpzXQ128Dn4hmt90gKLSKkEbDtjY4HXj9O6Z/
ZD9kLFsqdyFaceSbYMWS46RqDMMzJTWb2uXz62OBE6B752S16O6AHosTnM4+H9A/A+6SZZU46Fgo
sWZR+IDhG9TX7mLy5lzUzIHb1qLbPOKlnjQrTRjlYmhcCkBoU2xNTbzbN8FunE0FKXLGDecO4wOy
WzocO9S7n6P+uLT5euFzSk4yGyLpjDQZPR3aGVmmHhByV2y+wcrULWMO+x3wJwEymhNGf7HFpt+f
Wqafk86mtzWUzdovpx07jXZ1Nwk94TjklxIoc0NUXM4r5Ihbyi+FE64ixtYCD7eV6ThA8O4qk7c7
gTQGnZUaGdhrxAcpIb/fgb13Tikr1ZAFWyUoQ0hJDtkttkQVJ4TKSPQ85mFNByOaNk0P25WOvVkn
Si/rSh6+Yn2Oex1Jja2kMQ8uN1DbMmHzoB+jFJ8rFxJ66DkF8CPZXB9Xwx5s35N1yE39DHOVR7jO
14rfM0FM67C1PK+jufJU16Bf7O1s3Ex2Inx/hrivYAEfHHrZ1O86Uz6yafQOZlIK8/NIlp6y1w3d
JFDGtMUXXq2lWKn2++zV9YoHRDtLrBRkte4mk7TI2U1YsxQHL6fAM4P5hO8eMdTY71VZsESfed2O
CErVKaWTUHCnRr4Bdyo6zInZiTRQW4YY8s69IjgQOI0RwOiluSRNRaL12SPKSSfw2Bg5DFGqWBPi
hGxN4VEc1acuRPxyJoDD9k+UoO+oj2WllGndBq/mKWCUyZ44/iHh4rkngpxBUv2FvucPsyM1TpjC
bDCcAMp9ouLsmxSXv32cDIEY4CmV0PGBwWPkz0S49uTzYjH7pDVsbf8fgALuQV6J2jUsDZP0bqDT
OpmzDSeZqWkDTQQhbSjdjRB40ohSnMCFMlmywHBxaPj9kxy7soEDb5iXlrk5xl2WDCaCkFQQJjkC
lCkcWRZPSj0vaVp8UE0GEwljSJFyd832GVpcI3gAK6GLjwQObrYD+69/KuH2WHO5HRVD38OuN7Cb
N5NFQ2p0IYsy7HJza5Z3Dpd3KzHwxKCD2o51AERQoBfdYAdi+KaWUMaPMavhAEutfx0KPwVX+w/2
78Sc/kJzNbOWTFNiN4iQOSV2urmemz5IgOa35cZmUz0EoYZScY7b4OQcUrdD26NF5EJNTTdH6gtg
nBaMpxFwNBAS5inIdTxdpmB0HkWXNMq/U2m8rsrvX0xFnrQXZOEBLadHhxr9gl8XihEXEke2i55T
egLY8AxeULDRN4wqgbHMT6ty5AcDv93WJyrZwxDlKJFpHzcb8YkuQGE3J9qEbV6xGpnbf6Nqz8dE
AmycKyCnFhahi9nzb2Lq/piis1oBWa9mVh+PsMEuYsUlsd5HJA8N1EAg5SmlFKGcANsB52md05KA
bgskdvFI7ad0R2BQ1OQ/d+HCApyR4LFXR+KQZ/O8yKyQDjv7cTDJBr5PHF305s8aLZOaIy+TwJ+Y
vxGzeY3c30Lzg9mvvyP+C9+jymlBT3bhMa/7W64rQXQQb+ZBswzcgRv2x2S8eudyxXNFW9+2iXoU
wHweUoN1UMu6s9JDyencl5GNhfrvgv4qU+1EaBfDyyGNkv4OQyTt0e7rRUvVBos8uguN6itQG/ul
VUbCk5BNI0DaT+lXCAftxSbgwz1O8ySLWX+igvKcO4T61m9vRFGICv/69QizdsFq6cSBXyvmXfjd
ZSfhkXmMXsbFvT38SPqrd8y0UCb0wypIBB6th3e1OQqCqLC8Rw0/4Q3/ed7HpnnHajbdyuna9fin
mR3hHiUkWfjlbaImkO/vEE+isjJM15NO7WOJsDdNQGk3X8lOZ6zMRbr8RFNLzeEIYrBHJkwPJYpB
wnmgon2xWEUxClfaPK1J7MHMvV/n0LTwvQBwgVM+xhHAHB+1DBvvAeYen1SFDe1yNLhv4GywbeDj
otbhXu9+MYfq6ylB5lDJM3hNYn79U/93Evic1RkC8nsgoT162FbKtRU26o8tmNfZHlsPAYSztMKr
MnD+gCqG02CGedsZb1LilGYtF8+CvWczQMuuIktH2gPjjxugHqRK9DRsdELAAXMetNf5C1JwZZao
Zu2o9ODHBUBKwIjb8zoRSG98VamI5xiUN6PCFQgKipMIxkJTOMVJ9ADjD4SSlluXewGDRZrIPHLn
Wz9twATEk7EDuL5Dysc4ZAUI0kPwWmnlE1t9WxzhSlzQl0PWHg7tkAKWLSiCQXHvhfhjnFIn9M4P
3es/70Z/iytXHjVnsWTt1X4LYUTNbF0kiM0UAPRZiW9mza4YfWMnVXYuZ+cYRa3WDcHe0Rt3seN3
7Y+Vmk7i/3y3PLP9sxJBugg58IRQq2AQKILAFeuL5PJHHrI0/hcE4dbs9cj54TJoJlI/NMLM+F8E
ivO0168Mthm/qLOR6Gw75dQyxJhGrup1UvDMPdhywamJRSiPE8zEGAEwa5eya28iYY6NpEc26O7B
dnytAgDkmBvgwdS9KHgRhK/PatUfRvQEKbki+QQPtVJ8MvR6TogHeCagXM979B47gmGmqamQo4Yd
lkiUkc8Om6B6FbLD0DZ78a/aq3yyxVmfGpBG4WSzmGK6GhNMkFyF/Bpa5ZnRoMftUrOkq6fnqSfO
RqCX1yDHtwQ7PBT4brmhtZ7OU7KT3dJo5LpdAqjZBDpGHwb+MmWKESyMo/43CcTNlkFvkwdGtAXQ
iWoC/Gjf2I1sC/uHYDI44qwKU3xDe3VUUyKBr35xg3tG1rgSrtTyDJuU23dVI1ev9+yTfMMM3qzJ
FluDEjdcnOR2lzkI3gM5flMRIyeZF1HBK+yMnYo8msHzOglrBMS+B5rHDKnKAYR8Vdmq+qTYyyq/
ckAbdhZ8MYb4XuQQ6P6z11l/i4eHqgykQ7D8/bFvakptpmmPkIi005jtu6R7fMT46YuezVW6Xd2H
yZNpIpiNre32RsvyBsopPkf4/9O8z5vtuhC9Kc4ovzufmf6MqLJsEUZn7e4ZEA4XQ/+dicDMbpmD
Bw+WMUDVwo9HUbNpeAg/2FRZ/MPT7/AP+gXXljc02X3XVr4g0QGnUPDVl7guvoGEl4hnz0F6Id3I
w9/SSovjK63Ci2oszvaA5X0TRHUA2W7FfPtBSKlxRfAKkDnCBrttXdtKlZGx8R8tAk2pM2hE89Rw
z2/AV7FWKWDoQUvMfGKvruvqeq12QKjJUaqeBEyXo798ftBVgKkIJKUOtiUzeyqQjj71tNOeMemd
SnKEqxLQUovQ2XXwOFDaWmyieRp1sFRLcYaS/OuiRJX71b8dizlSmX50srdiboCQPtp8VUbtfXb0
KTDyhh8OOR7wplVLl8IV5JTh1pNw8ebJYr8kynvRHNLnt9b9LqFFGFQCViWepQXVvjIBE8UcW3zi
8hVYlNk7K3JaHjbrQ/YHtLtO/ypSc1bjVLKO3DWkmxwWN4gFf55ZfQ+vRssq0exuBEh9eb+TfsNJ
+xJRlIphdWtYlWuHIYx61RFIM4xXUfU2aQhszmfebnKDtHnJ/ckRH81BsAtGjhSkhCHRCqwAxjWN
Mq6rZ4kVX6K1yVBDoDXz6aooc4bs3PHsttSLDNZ7Nx85MLvA0L4j5g4NjU3va4LuCDqGYvxqg0va
h6zqUkcjAEokEm/uBQ23x0cIfSy01MH7P+/rQnej121xYIrBVfh9mfJjExon/gbZoJ6rg/w3wqTC
5N7EE/K8BgQBL6+wnLDGD7oD0IPchu0WTq5yKnapi/oqXom48Eejhg329P345rv+URFtdNFF1xww
Ca8qH8R2f1ZvvGYPlr6F7X2myQCPMboMOIZvacdGFvY7mxidEZLS0yAFpwNB+pm2Z9W/cSJDttEt
oFWvU9ztVO4Xh85DOzsguP8ChSH80xMcqOasqerVaFl4I6PV6GXF2IP/Zgw0gbZJeRpx/YBxGVgw
pwT0j19Lj6rJF81a4FHxbWtHgDk6ZmIjS+RnZpiGv6DrGYomIeQxAtC2bt36uX9x0BIbNPcQaQkz
c/0DaCp2mmLk5my11xNxUC0/zZrlWJQhBYboZNMsrC9Bi/8PV+l7nkeesHtGbEIZs/XZmk6RH5UY
J8nvfugOyp5P3rCZZNX0xWFNtxvLUC3I1wrbslOIqa2nsW/2HUun0YlKAOlZZIidKyhBHRq54W8g
np7XlOQV5u+jAfRo8KbBmNrbUcVUJi05/9BuA0holBCrlL1bzX8+L1R1YIyFq9R7mc354nyayr9j
drIg5hPhe0Vm5kKfqRln2uKtRPdKjJkGxp9hiRtANKS+ijr4TbLscE9zR06bNap7XMF0wd8NYetr
6oThvfUPFbAXfokeNfbLOngXM4CQ02bAANpFECD47BDVZhPc4k97NaTOZCRHK2easUShKVJxuUoP
rgN3mXyQ0NjMmlYp5nHc74hgwLtx/K2ljfx61Eqg7wak87bQsiV7OLSQZZawt9KUDbDFXZNOutGa
UzXYkEP5ol+HKgZOZB/+K7fn3fiw4VNgNuxahn4PJpoJXGoHxIWTXP3Ku/yNIa1cWQtjlryCyx+r
1raO04gfUNKOKwKVgJr4OwIyxx/RTe21TLSuAiJ9Cileo6grQrdLq6HgDxYrQXzFNWuu5jRWMa6c
qglkMYTANuXs4BQfvLEYh6JPUof2U2pfWyN1PU+Lk8DckJFsvNw4ziQEIyq3MPof/NU9MLz6Hx07
qidj0foYYJDKCRLnA6jU6HyPMVf1mpylr1xAv5BXSHbJ8fZv6W/sDU5iuwCuv6dMlxEmINjVqfxb
nkiEWAZRy6GS+Opz34YpQvCOis4NGj0mtKwbaDADSw/YVYzGUbTy8RniLwgDJ0tuOW62yMu44QZD
+npQF/EwNQ/KQI7aOdxYIGQfeaXsGN0lTn2YNTCLr8pf5+siwHXnvI3HcnhIivLbUrxSQNrgiRa0
Z2t3QQ2kHVMhxXg/1bSz30FaCthF67AHeoZC2AwBLlNFhIKhSzQmxRPgdgLZMs9t390TiGHAki5i
focjpr490+iQ/h6N8jf6AvP2Gx/vwRbJxSgDvb6e+98znJxI2r5+iikjOiHfKgtBjXcSj4Zn0vht
1+FQzXPa805GxD3CMleROb8VjinETsM/kX1185LVeJTzhQitqX8pq6krZe/mfbj+7YqTxUx/Q0AF
d3z3bbEtwj1ImlXDp+IXKUqdfSEvz02RZ9vlIM3tazu2fQTo8Cfw08xl3+Z574ZvX1YIGTaBzGyF
h+8OPLFnV9f+feqIITFJz5skzHb/Uj1C53Y0VBG3KWuDUkvwHKzQA5c+t/Bf2OCpuVEgicFG10Zk
YDhb8SyUnmukIVN3ZULBm1oeyTESIhgDPNHugNQ36fhgwqW/SfF0NXFce8mYp4vGmrhvosek/URm
/zORfu+VMC/rBXmJ1jl6tOnmNaXAHS/b2cWqtDIKZkxtZm0RI+Vxv5oMNmCKe/eiKLgGSaDFGKUy
Q9Cl0Fu3vDWi4muVn4DAyhQVrjbwA3CN4KNZDFNVGoDvMbzdTU5krUpl80HcjdNh04t8z2ZTEHE/
IVXxqcJtUdltM+EuOWdRocHp9Xv4xUVC8TisEmgEsTql4LjzkGBgxcLcvhVuXB8v3J5A2G/VC0a+
ugCuSg6COVP+8m/R9KGivwHRxe6U4m/+1zMvKtybqkgTFt4Qg6cIsjjutg784WBJpO4L1KDRbOuN
ovLiPbQr3nOgmP4sGUrdeSc8qoYal33zkBnQYNTBvacFcmGk0NRKAbCXMuUeZylPTDAd2xkEUNVb
JgQ4rLcY/wLTcf+k66Bd3zqkx0fLtgyeWkzg8TIeqG+hqTfZN2QDHiuDSmfliwmaPrTSGf36hRsz
hZwLslsElbdlDVaPhPRr6Cn3bnWQ9Hz0QAx/SA17PZSL85iot6LYBbacYdVSTCgpZYci1F4+XoIf
SD7pcPfXQXf5Q2Pu8kTRHl0lh8QdccqbBEVufkkuQnCeeV7/0PKkVbOKaml4FXHsabyk0lJcj8d6
YIeMxjNkN5Z0PNUMsjnATMwsW6SahvSkZImO/Fzgscq7uLEt8wCAJRbZ6pTPeygdyEnjVDkSwqXv
Tf5wVppiuPHXZIL7bAtRWfWfCzyIewXaRdGH+oJL3xITS0cQEt39a5MR0pr593oGCT+UfY5W4cjP
iQktj/R3katg3AyhBwoepJQbx+RYZ27Q6SXu58wbbtZJtK0RPu/YPZgp5mlyyTyy6zFTNKXiaF2+
+GF9XtHp3aP/EVDPWsRR6yfLfXDL+mKlDoxRtiaqyGkol/Yn76JTrO+JOVlsV20NSU3Xo+TeMV4p
VSrbdOdr67JUolClK5DNcej8EtTVcML4I3vlHsMUDMk5XaVKMMiyUm2o0oeVlbtMq2hoOth6+nWu
R4D4r2ffXehUx74vlMkevst9bvmdzGHNwEUiue8nQvU088Qx/il6lSb7kvGdaS2cdAX8g/uKzEaB
WfT5EWxKHtokUE61io2M1VDXM6z1gJLkjXgOPin4Vj+nC41XloRbl3HAGixY1K2PNUAHS9GAFZI0
EngyoOmsKWXRlTlFWfppwffyxqk3h6HBWyyg+FWfq9CafMBk2xd+diBxoLRuPRDZzU/8AykCR37J
w+wHkqD7pLtKV8beDVi3nsUWxQCFKhDe0fbLXE+5zF8FfqRk2lQL6hKMrpZDaApET+uSeJ5XOuNq
uFaFsw7nTW0z1VYR3xXUgBmxPVtRlPA4TQx2VzGWP+wJlwnM0RagZK1DENfUtkhAQ3OkJpEJkM8s
xhyaxqJUuKWKy4pmjOgfwXKfl6wPy6LDuqaX/0jZ4h+Lq//UhJKD32CCPlK29lNYwdBT5wN0yybV
O5lVmM+UlJJPLLWnn0IDdQpVKVgnHrGKaGdFrbjOZTMS3lN9ALfFoR1HkFobhZ15EMiLsM8J5axv
Mz0blrjxAwu/wCcBefIQDJCvWEMQAP4roVunGufn/FuYJQLuN+U0/a2EYWwqMELshoMNXU95wE+w
56r8sDB/TnZHZrY9b1aNVbBF5tIq3LtLuDJAyhyvWkJcWBuPsXK9iUlc8QkKgxupLGoG9cdUXiFU
7pGmcaYSKH1jem7IJWbZFxV1K5xj6CJZ0+wEUCjspav9kSAFVTQGl6nPYYpfl3p7bigt8XHiN+bQ
bz3g9FROqxDNB9jBjQlgd6hsbGPQAnzKH2Huo6Iz8WkOM6JCrZdYs3xwCANkeGC2eXw8rFkkY8vR
/tNMgMhGZ79cgCjgQq4B1AiSJhbIrFvRUfyMvH0ST7isWOvWizi5wcypPxpXbnT0pZuoP+VQs5Te
m+JcS2DNmrPhfwVVimIN4MKx8eogjbQkndETJTtqQI85I/EJLMw7ydcjHrrU5U5fShyH90lHbtwG
YbLqS0tMXTrr5CiE4/8Ctn/lsu+ejoWgn5ERjFTPHgp3NUjRw+jHaz730dV55lwGELx3cxrkaiqJ
3U6Gwi0QlKMkEkDkegqaqrwNCF3M2ZouJoTPLQ38R9Bwd1rNt4z22Suyp7CNzOGpRULBjgUskmr/
Oox5xT18PQCYBFocneY7J5HseaxrUroVW7LG3ysYtmSzflpccWe7+n2TdEMJRF1NSS9OHl1/og0e
Oj/z4ctJOZUw6RR7eiwmLJw+9v+dUDLMygtZ3pfNs3WvE3dor7SoQyjAXAyhfHAOcSGYDX6AK4Bu
afBepHTCLuvQoHW1j0VUU+TvO772XxM4+3SnUC7GviwNVZest4NNmbY8WY91GOkwzuPS3aJRRXbj
A4VrJjOC4tPxLSftefyLXh23NPJjS++hc4RNAbmXJI6KTyo/GXuRblNqBZnYCYkb2wpPzyuwlqM3
yxaaROx0BgMN0hCXg/LfnAVSbt2bxkPXFLmzclWp3eoWkKSeetvcvjHlxRHn2YFwbosGrV102hsX
Sj/Zd8Np7YCZ6eZppVkPa7eXFN9bCMoTC9b723gmeBw5r5pFkKRILNHuU5OEx7w32GH5KHLkRmzl
/sNX60YZkw42Nc07CJu4hAgQ1m/jQuaGsNWeVAYLMZvxGzl6Wca5KnbH98ks9K984Ncdgu6bKQKY
Kn4g/pzkmun6RCf+2HSzF4YSKHxVsr92QiAmnvZwFwwO6O6YwpPA6T05I3C4AZ1ShtNGqglUvtj/
qFheAh4mQV0L/ic8pdIWjChJ4OkngdzSqOygCki+vb72Qc/P7LKmn+gOi4rDx9X1dJTDxVYOjv/3
DtZ8rzU5zHBD9vEyxhXJGcQFKP7HEVe5Jews6x0mxnOMHfao1YHV7eDP9pboh97dhLtD4DmB6DiR
cs8iGKVO/euP4/giArn2WW1UCJCpUu2vYP1SqnVNXshdwq+X2ejQdEGu+6QGqLJrlOcrjEzMitxi
CFmjFNQcu6kZmjVy8ArTkT9SMfXjZocUFVSqCG9Mica03VmjsPsl8Eql48tQfQ/OHwRfHp1i/xBa
xa9ds8rltz6wlDLGA1LLNJbVl+8taLq7dopQHn9zfAQj8j1w/HTGrHFJudpK83rKlC0xPdsyB9h3
QRXpvca78/u+U2Psx+efSy8tiTzcsGzCe9CiP3TFzCvpCcW0J3dZ7+NZ7BEkaMrsF1CKY4IRJvIA
sQWTENvbKfJrEmDGpBGTCvKOjfoDD2T/WZBcsa1GsN/29IBjWusjHkauG4NsmltkMakGCM8u1w/y
2ydP0/OrkJOCIr06gMNLvAlQrQoM9kwN/0teZD+QLTnxlG35a6fEpN2nktYKtgeeO4m3/0vmALP9
re/MLDZfsRq1MOXhccD1ksfOAdE8iAUWEX5h1KPxIku76pTioNjxHqw1rNZQnFJHZFdrVkkv0dHc
uV573Emu/RCvVLmLxcN/sdUGB+cYxYKAOHhFJSyEP1iQkNMISC8AqMhJcrZBFVu0qexZIqp6uX8h
HlJkBAmwcc5A/DFvvXF1Rl3o6RgwIfxafteQrrH6N3peRhNd5VGg7Nzzg+iXDC3SoMXJtYTjW7M0
GDgTgdCrGK/nlhal4C4scRjaszJ0MQ21853OxhYyHrE2FHTpp1j3SsvHLLgh6SIL9+YJCmI+CGIw
iGjium/RoPlqsNZIGkFhi9zNXJ5FaImEqCQlZMouR5I5kIkVvt3CRkdbHGMYifjlA82uzoDia6Ie
mHhLiMkXzjE3Jy2xJyL0Ej2G0juDtoarn7Gop8+Z63RoE3d85q5YhHO5gvFXg35sGFhH6Vdjngrf
K4s/LHfWm64ZEEO7rpl4QFSTKCS8jggzvdOGJogIp20ZY7hJ3aVaKeAd6VJCrKeonyInlR6J7ve0
4/8i8n0Scrzn6Gh1ZQWkPTGUEA/aIIIm2LV0puakDOyGku65DT3CtpsNNijv2UDlOKOgvrkHUvOC
G4LIBktnokc6rPpC3bP33NQ/Igj6Vco8YKfPiWwhuXv52TCn2tsErtbC/V9U3LVV3fBBlTBlEOjL
aCMzZYbz6SYENRQRqzsc/3sOex/pupLtxmzjGS7k8Uts9wCh+z4/Ad8kvC24tNGLd7Js9yS2ISU6
b1a+9yZI0RkTiAfS6/Dm6l+WlijKjs5M0DPGPOByxgd2K1he0EEqCVBShgZKliqXUGq1BVusC2qK
ubz0PbG6pJaBBbDl3Iry5yWkb+BxQl+VSO492tWNxi/CV6ZTKI6PzucxNObb0NbUQjoZEs00Rvcj
zSPc+hBdg5r1WZtq3L+oMEvJxWQ2PktqxTFWSznJ10FwR3Wb1ud2AVLQgNB031vEAj/XTv5xXPD5
qX06A/X7aKs7fpc4VuovmoxFaTXxVQUkc+WSCQMj7yrdH3qOGCRU/eWF4vQktXL7Cm0Rhem4zmHO
vdVRbNgH7guDsJ3GnF9u52D9OQSpHUGtq8jayx7wFE/aW9F78MOyoKDD1ERlKHaT/XQthET6CM6Z
dMz5gHrXDSWwijxc/S73SCR0PIomqUKEdiU/dFbg2AiNsPizbzdSYRAYwTQkt//PAe8GXDv9agAF
Y7rrHCF/JHpnjL2bIi4/ztn8Q7ISNa58ttJIRWtvT23xgRTMoqIcZ4qVOX2X7STGPLJRnMGDSgc/
PX3KG51DiHAFD3Jg5mKbSJKJhbASNhMck8HevCFD8Z/R5S0TZWCvytx4wZfT6kCL9NCyJ2W5ir+o
ID7UAOSIqTjUDMCI4eOUrpPpCkwrt90WueweoZEDBFKkIsAroTJ38GcYI4q+ltK6MQBxKPEcLXo9
PjgLedwHuXryNEnarITn59SJX0RYrEkXTmQ1Ci8qKiG//c49XvCdxHqH64F6xHfIzOBgcoEDlUPX
0dgbBvu0qF703huhYq/iaKHgIUFApUQfOxu1O133OiEXIog496cEddnNN87unU/s/uT1Gf87jKG7
8oje36eO8CqhF4fpcHURg0brud4dV3hwSSsmBGuQ52GivBbMm9RMWMPrCTLsC0w0Oh3OmRQrhnDq
rTgQUGl/Np1qo4RY7wSyZQu/3d8jiYXBzRRlGWnZnHkHSTO9SB3tvx//G4oYY87sqhQaGU0EnPJt
yNp/gtBlq4E8nsPMUT/vR7pHlgykrRYbrwIxjgdVTRN1rhUJelBtzvQlCqh3d+sm0htPtG4iuGvA
3FPGl2ODPae4lanuuVe8gr/LyZPrUkNp0qSEd0IUmks9G58VVsnVVZg6TmAhuh5keWD39qgyiaUM
iSetBykOHS9tZqUV9ETHOm4REPVKRXCI3TxLrh8iJS1MIVP1sr2xPxIB/4zD+iaC9ziVyCu8s+NG
TTorh9wdAUwTZjUqYKNwIFHlgPpN7uVLfqHH1H0l7lOT8V8sbKKsGkbXCE8oj4S3BH+THM9m9I6h
7bQl4P+arHAlEtjUeMuqr50xZo8Kq3bI1hL9v57+ktcNKDMiefTviOtsshHO/yQwSjMFKqT5ub0b
kOn/yjbpbWianXqJDc9DiouKMJlh4Ojl2qnlJW4Fk2US9KUJfhckm09GKvhgtqwUkdJjF9wl1bT8
sHYG85SkB/OnbyZh3XS+w6WZqwkigeglmkQDrJDYqhUJ7OAb3EfGuX8fq29x6rfbGtbANi+CdTMN
p6wmFFR92EK57c6bvK86pqkqMfqLSFomvF4p3L8w9iTDF0OmDJ4jjdP+x7b92a1qyZ7fMDXT4aYk
x1tfOLro8sKEiHECbDyDIf2O9J63arHNOj1MLZ216Ifz1ld8oDCEb1Gvn/8HsGdSlOREOgg4FeJU
v4lz4Gj6+pZjAYTeMzQ1pDthpaTEnDpHm2C9v3FqSMEqKOMBNji4p/EUNNu1cvJpx9T9oc+HJlNP
PuhQu5lTJE8p5YwKrDhfJlTXzNOuvXfSFnnqLI1rPOTocYMCY04dg6jHj9REDc0yUUVUGaNHY6v2
tw0zXqg4G6qx5d/JqxqAPqUBgBwVnoI1OYrqy3spQGlQ8Cc75EtdlBvVhCnILUCk0bM0s04My3y1
XMLG+ZyKoRMazLknJOg4SuTGT1Rsu7kz60N8mwtcoVUuIMCaaJdYjbC6sMc5PWChDC+arogxiM79
cUKLL3LceaS6U5UimcT2embhd4M5ep7vHfDOGExHtqUMW/QyyjJC20Dy6RLM7nhPivLQhXzB/3P/
SA9zVEhSXu5SvCsFBjpBp0qb+MkLn8vAK8waT+J1CgTIZ4MZhjJ3nK1Sg+MYVens2OVJ3rXSgn4O
DyxQ3UOo7axNNReaJnVPW4RG4/vIUmZTXnGNM4/c95WWqhk2Zxv66/cnxEcIFJrZCK1NskD0k2QL
NlZk1jCoX0dCziXQwu/hF52/f9oC3bb9N1ROrd6Pz+PdmYKWtEKH+eJJUnkUK3svXn623BE2/3PV
LNUob0J59yAipatoicZnefmPPFRyvivWyJl6JrpOW3bXfhxOrgq12+qMF4Q7vIZgOGVj5I7y6F+e
sjCFy0fqnCmIVWFz9ffOvQWXp7WigTz8+TEoH/4GwHtSx623YAnlOgenoVFv6dF8iwO/02+sEOSb
gcTXDdneKpYBhLVwnc5VpMK0cabjmvah3SatBBNkU1pgtkXxbj33yz0d81rvLdOLMo8y2HsdO5we
HhIihKn/Rcd6bz5cWynCLEy7ABRj+symAkRSJ6P+WM3ExKCBj1z2ls0ok2G/t2FQDcC9H8awq3L8
DP37m/PVPzVHmNjjnNvrRJ81QHZQugD3165wB8BFFuZ/3zq46yfG1deNPuVHrV4pnywr483hoVP/
zT5GfONiSwkMhqf0LPirj7CRJX/14RRdNvHf8YKtTqxP0gR5pHYO03n+CZQct8bf+O36mPnssgsK
Y6KPh4yiHhyX3snBEYU5mIXaanm7OeVu3278iJZw8Fzey2Dt5o79hD85XFakjhsCGSq7ElRd5S6M
ZAj4ZtoHCC23/PxcjNFLL6MAje4Bx+KKeXijwrNDMW3xGdYuoFXvD73Hve9fnIoNFlVOxvS2egd2
fdKWXOcWob2oKNHPFmsT3YWqxgQYAZBTKxrRhvgf3Cv2lunPbh/gbMQVXEz8X9DZ0Depl5WfQzQw
if1K94BrteYK/PY6MZ7r6FNjMd6GIFmuzZ1zyiHCDj9Vjmfw5rjSFbb7hju4SfvteYSSefIG1rtf
vO7bak7ObGT3RyezoZ+iG2fKRAFvA5Y4/cGJacN/wVFmXspmZqIGL1ma/aMnmfpmgLU5Wi24nlqn
E572bc53mh+2Oc5hUt7wYCg3MsjP1G3X2zbASFJXNymiwR3syz3tPVx2L697MOCjJacw695m8eFm
m/lQ4qAby7nwXKy3ccQiY2AaCL/2GpRjRo3/Mue1SAJ/Xv75JiW9YXqene8mWggnfI4Tu67l3p3j
9bsR0hQxU5VxsXu7LfuNrPwazXLpr7CLAmMiXX0x4L32l9i7AjhUraFW1qiR2hJwAexT75Jr9t8w
9H8xOHFa7uFu2Dy0QwcZupodv9V6Y1lTJNGpQ7qAJMX/36On+4zbjWdUonCqL8aJiQMZ29hrYMLq
x+CkgTF1b1Zu6yLR+XRR6OjKJ0OprbXiGm4CE5RcVFbY59SNyGiwA0dSurgF+MOBxuMe35pIXyT9
FuucrnFGaQq1fhE3TLogDfgSPI+3aKQiGpZSC7zpOEXbG6hxZ1EJs/H9Wk4mxD8BJFCBAfwTTYvm
MP/xyDzxmabKOkT4jqO16JkvlpmW+R5J5me49/vVGC3aW25dhIK+tmDW6JkX0U/n1qmQdxrtrQ1O
revpOiiKceK20eWSucScpmhyrYJwZD9oPI5szfDqhYmLqfnXRihthJqj2b0nRGneUUY8SxULu/ha
DtJqaFdrnfG7RKZQXEMCLsjTW0eJz25Ed7NFhz8uzfooqGuew+olF5XuoF8+ZqxNijQaMwWhjt3V
l/exuHuOrk4+aWLiX4ydq7hYXZrf1FJXO853aN3S3vs6kekHhhQimVFeepCYkiEmHl+h8kkNfFTP
gXRlqCATIPlOF4TEsKuAnzL8AVhMab7uZjTdUTYw0RHTM+z8mN95APdEPMSwkiK596FO/U1XwgkH
z389ftRncK5l30gGf0ObpUKkU/5yKL0Sgh3+O0WaEN6Gbp4RJmL8zc6cjnyHXpF5R+l4raP76oVW
IsJhA6cPQ/BIHi0o1uOm2SPdb7N4vXtOMymJM7g+YShsxMw5vOEJQdsUkqahuextrt11ekHboim7
Z3d1dRZwi8ci+7N+ds4tI6IME94060f0UxgONCglmRQKBH8yO+tOyrg7KE1pvOb+oQk2MwhbN/Bm
IqvDAfY0bMqhsEEeaxNR9u5JF/WGED1rqk84xf847l+go1oeNVkU1iiyco7OADZkGnTtvtAh1IL/
exgMaAppxkKh5ncrkZij2ZeyfOsfeKWFltP+5xrD87ehzxD3i1y/jGDuRC0sLiXyJhwft5ESqK9y
JecYmlDM5ocPrzNIWO6YPDmSoL8Q/0HZpoiBm3cWSTIje3gIo+NnVW9mKOCDqKaFFnE8lpB8npf4
VIu3vOfOa4qTyKnqkAsccKdugZU3JRiorTNt1GBW7iRPvgkWiHTd5M0TPabRasb9td4LmEfGS03/
ZxGxiADeyLb6X26ndUZilVjTYg4FYPdv1fhESHzxu1vb+smsvzOjOB/qbigNrpjTaQ/VP36rAvTf
fu6cigGqoJiEhhCligu67Xsxknz4SqMCLTOQVw0EJtJw0ThTF8g4pibivphQMMUujcHSFGol8wEt
mAaXebvZPn+beMQuuM2W4JomeU9FwtJ2ATLEMKv6D+AjlXnZ+14pUGSntFZDYUh9icHkZ1hNMe7S
y7tySwR9l8xWYKnoZ6enB2wuoAxWJHDPIeRDgH988JrHgWjXTE/3THM1Wv2yeCFqXrhGsn2XeP8g
72Dx1kl/VHvMj6DcXFGxkqxE9wJNFFG8U2GQnoLwrMT+ARbi8gMJJAn+ak7VnAsc/fSgzWQoqnW5
ilnO/RSORGafrR0J2ws+u08jao4qAjDGnzi97+CZL1z/PyjlYkIWM1Hrn6FO7R1CO1m576mpXW5P
6LwbC+PkoK+A4M3sPEZKb1MemUCfw+rbliY2kRUHd9BApvHO51XVUVpURENtcKN1AJGyhKavsYLY
2DsOtEsh+cqPnQp8lLMBvD3cjypDaY3Tyr374w41pZD5fBq3jzAHf7clVZZ10HuIh8m9/Q/79HCy
9uCX8U28DMgTeyO6k7gQxhUaZ7wTlXV0iRj6S1XtBmv3AM3j5B0aISEZf/l8Gba8xjqaYH2F3MB2
R8qRHAzRP/u3/bSbrIMpWX0YMbzEqUKsuAgfzhc7jATU3R0nj/NkKhNMavZ93f9RYrCkITlAJcOs
fxF7qYLThrxu8AqGSQLH2KpRYa9cxGbkVM9HKi3mszDKFCm/8t4asabLoM4/CW728S4clXmsWCCf
LaxR01YZ2gtpiZ+xuoZInG/4PmCk0+4w70s1VT5XruxYiub3o3TA/P3QE5cVEZiYUnJnfJc+Uyn3
Ip0O7Ao8M/0hPIhHrh3NySVy3cJ2Y6FlFvCXCzhMQ3zPqi0d1Zmfc5LulUYPqil/2rx9m/5spNk7
49WZ0WVlQHmSSEKOAlHQTxFVAQYUoQG801BzeE0fFzisA+vX7qkZ15oM9WQcQHt/S7+eRFMOIe03
2FXS1rJxNEYw8rBoggzjthx4RbmGekcinIZ7pQyWgduevYcR/Lh+aiArHnaVJvArhuHIPgBgyRrB
0MWkAaXw2pxPAQa08X3p4FyY3bPuUVr4KWeMJzTD1ntbKUYLL0jiM/MsmT6WsA77POxtigj3J530
nBSPwJyz0vXFVkKTc5xH3DGfW81T6IK+yBunQ0TKTBbiomIX+3VYSH4woIxBAUx7ElgPrRF6vl9n
ta4mLmuSrvImK6swVikIkXXCLTzzkkR70ta8ZZ8Q9AwdRERzIu1/j5r7FERGo+snzlCVCTsUJLv8
z/isUONPfqfIdtdIAWvHDUHhXn83g17k2/8f5wsX6hEIWK2gdkzbjJeDbimmvBU2lJpqo/pvmw29
Ztbd8D29l5B6QUg7DcHMJ558Lmlx9IZqAws3M5FnwlKpHuxMeuY3TP2sUeev726Lp3O0KDy3rw/S
eMnaFOIIz7fcqjlN/ta+D2/fM1GqI5FUz2aJs56W/962NqkRqkPiU0rmYcbvk6nyqPREJHdb7AuY
qUBENGNfhk/r4rv95ALk0wp5KZupR6i6/qDQmMV0Ib9rOmEl5eb3+kmggOFkFSbh5oZ0/IDC7TKZ
lkRaidwrfUsN8IMnNlnS0lTJ0iTTQk5dQQIQoSmE4vTeqeAB75FUDMqw2pAFty7XhoH3gPebCn/f
T1UiEJ0I9n1pGEkNRspC4ngZJ9dntU9xxMlGUU4F9lI6j3Y4qQ4wD4RR1LYNPGtzfFu+SSNNSd6C
Bj4dryaspFjH2QnRULAVhQ1fm65Q+TnrORBwb23d6n4TVpV2MopL4XiY2XEq6PpMR8Wm1BYGWs/P
Lvm7hWdn3dPUw9XmxsK9p8i3taOaLCILPBO8s9QLrpaDa1qVH3Gqv71NLGq2yEhfBscxYrLLtegD
8tKaZD1umhlkhvALD6jr8SP7Pr7TtTsB4+9umm5qU/2ueDBsR1Ha6zMPQ7SCdNmyWGNvHyHYk68N
puoINTr87dF2Hy3uJ0ha7c3++lQzv3WYI6LoEpExk1CEvlmDSxUhCA/+eg3xiHq3tuWL4pmONdgB
0u/J7tjwoK3CebfPsoEkzDvrEyyJNGwPs3i9XeG/Xef5hZUPSMKJxn3p9/ipyioLTIVMnR+dZ2OM
wpRXKfPGwwAspKSKl0qHf+73jIklMOsShFvjLjXzhKzUmnr5N7ujhzSV6CBWnTmvFUap8dyEV3mh
i9pf1dhTZLaDWstfWCHjsCwkyFAsBsIUI2HctUCaFlyFxjwi+DrPSR5NjhTh60v9lE4hE9V1YeNQ
QRVni71TmVmzUW4ngDO60F8+boKul8P9KHEvF/WJBsCaoGWEijWJ3lmbi06+bv0V/PkBLZr7xGi5
NFOyeVLU0dCwLZkO4m4ndGELSndTTD4TSZbK2s4VGq/AxsKynqHm9x+k7WXEknejWCloUqPeFEgU
W/TjMq5hMiTNKDUk+YZsXu0fITkBqWE2igIQBRfNKolLqi5jCb4d9dYqiMcNVa1BnfAECJZfX4D/
r4lnvuXEN6WvP0RD5GPwBSNwXmLq4X6IREOYd9CUZMdF08v2pMrLF/shnYfsLFCwr3QwR/t3Oaik
u4R5vmwvI0yAzaofxmuiyTvMZ9/ovIDWBbBlOCfPyZsrnkmVfN36i2+xofV6cAgiY2VrsonibK87
vJh9AmJG+Dr9JHiTO/rxLceKdk3+KGiBAW6X2rcT6i2U513RVnC6ZhVNoQMXGuc1onNLVkTkoMCI
b18PwKtIc5nudvwfjzcZPyU0d0nUKwFBOgo2h5mfLHznqS1GyWPK3qYsgPmtLIG2C4Rzc9jCPLa1
QHtBFaGVPC0ls38FWW8G7lJNc3kKMly4oJD3o+tSCB7wgUw6YjFbKxR/2zd8c4/G7m/9NRtVdJEp
+1VVF033p6C4ApnZLL66KeWwEtPL/3/GoTloPmuBHKFUlihkRu8EpLxEw0rdK5W725CxT/Njswjf
RwrhvH77TbEnRQyACWsaj5DvBjARLTAHuQ5guqne/CY4RYOIKamCAvlaJ7l9FbegXkjVOQN5LXQA
FXxeW6Iu77tQHG7lnEjsaseFnOGHpsDdQ4IyKCLeeMTB3UZSTrgRpAOfvwwxqwi2GEkIqv1CcBmf
W9/eipJj8H0a1kVgbBO1DFNfSGSGv1vU69q+VOUOmwz3ITeuY0FLN2FrYU1P7tNXOCqj61eDCY8y
qDnb24hCdppqpObvOdjWJ3OIbFWlGIlZpv2FDx7vv9O04VwIeZailZgOHiUy7OL/DYZpsVYuhPg5
oNHerEeo1W67bhRdJ8YrbHz3ak0NEk2zmoq8B01rFV7Z6vCRXD5QLDU3fy4VDWIkjP7uJfnoaKI0
PdA0MTxUvciFxSqCwOQCgBum9FU9Okig1MHc0JTK3jMbPnKLft5YtOsOIouIUJDKl36fxmIT8Isy
+2HpDknETzijQoCCHODfn9qC6y4CUbbD3mq/6VKJEZQPnmKwzsXz8pjR1orYmnRT7wmnfkTQb40Q
kzqcDKbOZv4xGhtdrs5QEyXcTy5MdtW25LHBJF5uE86wvu/41a5JPXc91wGNL7Mib/04f6r4UkS6
Q4YWuuBnCHfKKX7MVBF+SlDTbM+qs3ByfQTOIx/MtVXiaeHq2yFeizPG0U1RRrkOYWUUCB366PGP
Oa3oulz4IyWvQZivvVkYwqunyksvHFK7wUTtPoeKLsYt8ty6qHWzIE4xFXcXX2l7/LJHOjFeiW+h
XePeYPFZ6Mir0GTxJfd9sxItSHaCa6OFol8BE5aSanrW9QDX38xvb5ojs6UJ9Zb8SR00i169qPM8
ddme3c/g9lKW1WVs7IKd0pUGD5qPBPe7CRiFpp+FkA2peIe0X88VHyIDtfnO2zvh/TKAsJP7UaB5
nj4/CfhkDNYmUSMixG56B5ZzYFXvT2AIpqhcztum2NL8y+2zLZ4tlqAD4ksHqrfSvQym5Vu66+Pr
tcAXf8Qb9IaFpVEpFTmhgoMMPZjKdpjxZNiyQjH8a890z+exrObTRUU1VH+kVOFyeVC5NvC/ZvE1
bJSr3FC/h8/0OmKNDo0txS2pYoHiwUY7J4GTOOqQ/uhS6hhzpfaKiMs1e+LdVK0MyT6Rr5vANuDz
hrHahRlGyk77w+JSrVoe41UZYUxX6j4i0hiIjZfdQHlBxG4YfAA7m/4/UzFxYpOUKXK2LMM3cSjP
qe1TAPDZRjjm7YMiOwU/1FQS3wzDcy8ug9BPj8ofL2FMabpVH2mMYOYniRKQyYldcfXf+zIiH7nB
W8EDdL+MvlrmO2kLzb2/7Ct5lVooZ/JL08dC15LMu45v+DYedYaJL028U4HkYq8AGf2aSLcKvmuv
PfD/tcCJCKk7Af9IZ26cKAtW9aHdl9/M0grqsbKyksweQykNnzncqnJhFlqX1O5GkBoOZfvmXOtl
VG72e/wYR4LKPtZWf2imylg0Lx5oM7XEPHyiU2ko9yk1Ws/ZT2a8YLlBAnD8+e7YkAyMP+wEDfkM
xMfYLattqxey5jWI6gJdEs0PUNKCqOJtxC3Rw79yXigsLa3yYj+2jLfdypeXLCv4a6PWAh3jhGPo
kcghsrNm5a+KQvcfx/ZOvx291zOGp3rWOzMXPWlx1X+DMw3V2sfq2WDDhfN453+vdCsqyuoDOEjo
R4OS1e+G4cqjUP/3koZrjvT+fbr7XvGNYi97VEWWubirdhW4Azff8s3llTh9R611AE63isdMLvpw
5RMZJldmN8OVtRPEQMEhr/sGBAMhwNn+Lpz9S/yWHkmDuFbXyjJ95mKA+oeaK3hGPdgLcSlmWaAX
DVxHXX41K2zGxWdlZwxJ9SMoFuFSTd/JMU8S7VpepoVuGhesUSS6rTVpb0pp8q6R5aDAHDQtCHND
TaCu1MefxRA4gBwwcWHUEXxgqj7UHD6AUym032YIVCJW4zLnvAUPU0wIOOjw89zlwHa972CJqi3L
RhJI07vebnbLewOb74ha9OcTqEU9lOP86ZOvjv83Hi1fwhEh9makAQ/ipjCrZXrXkC2UOUZipndF
Bmg4lUb0x3nPkLGlwurJ5f5MNmb6RMpNwz0KnehnBkzh+863hMtitZ2czhur5IsMu/QixdorOnpw
OU9+Tgws8aVj80YbCbVYz5viqE8S6kG3fPoKnmihXhgSRY+ypqtmF33FlIQyDa7ww+LixxVNcDUo
6ERN2B4DU/RMBvHxCdqb32jv9h/6CNKaP6Vqf7e0LE8pg5KJn45pA6LBAPcGbEAm9BwDKDDdBADo
U+iCMyI39/Cl64YzZZmf3liJyX9XeVWjTgTwkE4Vg7TjhCnMJhred/xsYViIpobo/XBft5yTilqs
SOGTJucyv4lpfTukZfQ4NIJ56fBtv/aL5MAKdYcBfROwpuW66BTQYQPCQC0Ut8R+h82TGK25/njA
ya3e4lJXjrKlkK5fXcKlHhnpIv0uM9IwAOYnP4zjNgKTCfu+mn8NtwPV74aHh9bU/QmOB5t0gDJb
gU6lmO3DQA9KUOMzbammV75MaS0fSMIEgCcXiI69kj4NcEMxLny0x8ziPg/qgPxB63qLbrl8MFAV
kbZ+Jesf/uTVVrFlGj1/sjJu6vHh0NxqGBoKSnZctbBVM1VFhaRMle3CCPhtPfOTEJ3Ah3bycMRP
j+bHj1J/6QGWSLJHJUsZ9AKugQjj2jPF/MDh7iwPc4YSXj9CI3FnJy5Lxs2uENZeEkjSeYD+hstz
7p48JnykIFVTcDI1yZL9iuqjbo1l2NFIT88QrPJtz5K/EU6+9QxTL9j2PnXqPtSXAidWRVpwaq9u
Jc9g8iHuVdxZihUmwSJnisapiaij8vVPJG918wZgq/XQv4QQkEnmar6kkD6khGCEvkMj4t5LSkSq
vLOp2/ah6mdPEadZ/tVplpJn/lalxgNtgXDB6JNfYtHcLLy8gLThc2ztlajye+hGWoyh3B+wJcHc
72QQWyZ9hG/O/IKgi7zp4jG1nZes/PbwmwnUEmTTLygv0Fu8XEou9IA8UI1ffHARVn0EcCh10YuT
W4bqKNfnn3zQwCoz+Is2a8c+eUZMlR30x1xLhF43ohjJJVZZfl3DT5uWaRK0HWdnbHzv2ixIIQOe
YK5nAJ9iVliPTbkjN8YvF+7HysK05YvwRLCGmFzL6MLa9UEG/29T1ljaFYvUglGtgL7gxmA/uyOe
2Tbjf0v1vWKZ6Rkfk/eIqhecjTkbVLtKp3qw8cjlL0tMThCYTIGIt6/tNyNJEytAR/2ArQu748ap
ZGWvG13BKHdlELIJFSxK8gFvGyXpnls93ahJEupJUyymEPVFvxQNJtQZYnECo6wr2UoVSnXOd+NJ
GAwYRvO723HaWf4npUZfbFE5YSQn1mA8F500JwkMQeOGDhFJGgk6IJcXr4zaf0Q0rNM9AB/82cXH
hzTndxddkr3Xefyj+IIVJtlEMp1eB/w3VfDXeY2dV2fcQH3gSu3Bc8ME6krQB2YRGZHOpuzRHkED
fsCapMbzT3V6oku0fqs1YYNrT+aQRohHXlEMBSTQQCz8dfohU7hJa/16t1pQFbGGsxNlCWLWT9s9
gEiqcIUVmQWmgioadepOCU+STGl7Lw6iFyiVrndZzMarMeF0Lz5wj4c3Hyx6pxFok8lrO1lRz25G
T08bLR7AuMyIl0K18ozTRicDLn0c/Is8xKIPKfbS65w10OZkjoCRXra/gYKCjSKdJYL7ZY9c5sPV
v2uF0HpTQU14HTU1Y0migyh4gTbaQFrtODoAdIaFSBa4FUK8NxQ4/fF19OPPJ5eyPCiZRO2X8M+a
4Zel81Uk9Nr9A76sEN5Yg3TGIbZyeiJkMW5NMC2IL7otjUp8Pw6LEc5CGogskRg/Qcx2Vye1sY00
e5+MlDorjVrKSJR7/eA1GJF7dcW5IjZWu82+x8JYd5jZwQeBtdGL318x4l5sV8Z0hFSGsYuMWFRN
qMbuRnzN/TaBZumhpDkU675ItRDITZrMKk8vR2c81eNVPUuZz106iKabr/VZpNvPsdH/S6vFbYyQ
TD/NnHvIS11XWs2mz4+2tp4iwDGFCzrr9DYFAzjF/yM0hT43SH0XqRjPZnNLDUujnquPOi65NU5q
xeUjb8tyUgR+2Ew77T/6lq7SrlsGqVtLQQPIlUNP8+B0hPL/kcOCk9N0+vSapjmqunV1Mj/DgmFf
zZZtEI+tW5Sy5365aKrm/1GndfiHkizPVkEQTLBgZXH93WB1/PCxltOHz4TROuuzJBRqAoA67Eex
8VTE3S2U7Zwa57QhnJPvAtVWLCMGz58XrI8JAkxAkAHPEf4OBapSBkyXNF4f5w2GqJP8PzF84eCq
WjeaZunMcpxxxTK5IesHyDTqmpvEUQG0kFFB3/wf++RjESmw6Riy8Cp9uAvswNnNwyuxRvuLVo71
aNeLXduZiCT3Z5dbXYMjl4pOSgN6dog8M/e3iuqY3HpC49uaZCxCl2k/GA+TDEIvd/KdHrrzpwsa
luNXdYsl4J3HD5P5WsIEg2/dejHwAd/CugZ5ZuCYPDs31aI51WalPwKxocptmXAkW7x0oFlF3PST
4pFGOy5weWuIuOJmIC/ze3ULMAVQhaHMAahJapP1fvXqlM89jGFy0YSmqv53Pbx8Ws4IqvTA6tZM
+v5+5SAmkqIKjRnhYcDEfHpcbn5dzU6MP0gi10blWsVAdORh3s8XufIHH8vJ5jKOpLRFiklGFbmJ
j/m9lcLW5Jpgrf/7PUXDQ3KnF8La8H8K0JgJPQDHJevEp/SMJ3mpkAJs5vBh8huM1ENuQOF0iYsB
ZbzaJkLrpfASrW06H8Jc3qHDUvcH+SvJy0T4AYMBJhYXMJJ1aR0WsN/glEwZ82cKfQL0CoqMnxxU
VpbtRI4ty1Os1uFDmlfevMx6nYeFAaapJon2UdZprqKMIJje6IPLGa1XaEZ+wDg3vFe9iORnEfZu
qXwP9Qtpx0+x3MWh26i2StleysN7AtYJfOrpzkBUwdIzAAvuvHkMmcqAbtLEsv72fMga+Fjjs3bJ
nxLiBrkrcG2ugnmjp4e0w5/nLPgbWLbi36YlnAWOH81t9TYjw3J0irS1pQU8M9i3LwP+JdKhIl4Z
YX5DoDPC2Hp+Moe0k550dBVmxXv3mUhXwusarjPQEMmJ/hPzz2D4zj/VzO0JaHm3YYzoCCMx/WmK
Gjw9wDr9WliEBsGIjvMgX0di0cU5Bwq6LCXCohecX8rCgfo2lx6WD30ZwfY9ROdPRD/XRdiAm/ak
4nBna41LG5GPuYcOv5PfHXvRu+N4wRPb7KbwjSj5u2MAaylLYGP6ehJ82vy8Xqxosuhi13cEgjxo
0gFTSZj1+MQEWxMMofrN9TyooVYSVmZ1NJ1ge3ukt+VKnw97mGdMyI+MI/t+qae59fWImo4qbKeE
4DgPFsSTlh91B2ye6bGQinzM4pZse2iSqoErLypksKgorsPJwWWJH7v0D3+5V1AOEfxvsRBSMOJr
qcv6CC62GOpMC8kDI2W4/y6BPzyvQe6gF+NWn92ae1ElPreNyEH3dEN5rxv2yYgfg8+Y76s0veYp
zwZ2UJ60j8IgTcZbknhAMgcXcA998A1AI33epW3Ean3yktuc9ilfSUydo5wwQR5LtaoxbH9p6uv/
iFDxxFO66He3fkrrViOkmZWKNjL1WgUXirD1Aeq8VxZtSqEXN9viE244doLSyt4TyimcHhTIed5i
CcNi5LfgHVsRnRueu4grWkskzjhECZOhyNDyfx40hwgRaJkLt5D8kZD8fFzfLUYumYkn9NrhGvAL
H3Os167rQaRnpUVdZzhRK0XnFEJfHroS220MX0Wq+k3o7wqlkdQ2OGTqY+P2b6Vzrs75OYmwF+Wg
jEoWKUIAvcqHzSN+mWJ2+Q6D0QzIKCAT97yBI0X5vNQvDljRy2eh2o80Fhwya4lde7WmfGIbkyRh
RJXdUam00lJu4sffvPC0/Eg9KBMj0f6OTqQEVDweY2l9uYsta+lqngOQL14OL4XeTaIZrL12wscu
pRtGdkWLtzcqDmbPXfeDL9wP8QY4IXrXH1cEcHcMU339er3jbyWMxADfQt0MCrLGvCEhRd+/DpxP
0kdIUDkoedvqAl1CISDgHdeKJxX2IVpiwvehCc909KUZDCwF9qvVzxI7NXy3uTq1CczUd0ij/p1X
VJl/dTpX81E8+R1vRGPbbDKM3dsHasSstHli6bxkDRns8M7I1BnfAAg1bjW6B9vP+2q+aMeDLiOS
KLHz/sDuY+23rglRQA4g0wpZe7pmH/NaSGYTqLR6WaykkqFXBaYptw/39HC/6lDErHD33ONJWnzX
rNE6icFLORvuaC9AoH+vl4SJemv9EKxaqH8yb6CNQ1hh8O35nZ78gHVqA6SztnRMsdMSrSRoLTCb
/YbROQ+MmMGYB2w790h+lnc9o0v8tfseEw+CYmB11SWcTqdGlkrqVEQtAiQHgDY6YjzPxAhH+dIY
yaSnc+1GH4NvMmlvXTUKq3SE7YJ1LaYUs6o17O5LFPIoIfP9t0v86yvQDT3NzgerUW24zfDUE29y
O7qwsA81xMSLkBaxqjm3i7HIJ9GWXill3NnEIeNwqYPfFDLqT7NYWqyFKvCPktI47jFMSd3kb/3t
kdgY3iF0o0yspxH7Nu2iYeOU34Ua3FYdgdryR1+RUdBwkiFjkd0bMeuEHT71b87EoeKiCljpd5Qj
KF8lbjpC3wVknnUS1ZOyo+tEsRSgh05T2WuUwU0YpdZSw/VON16lQ/7t0I9WAtEMpDk7VnJ1ptka
dJ/IrwvZ4mKqGVmw9X2ChlfHZ6yzDRXwNLDuST9g/h5aWcijPdBy86MWR29624SXIYOJORksXwJQ
U4C/hHAT9bkQTcbhFKRrl+Ah8Fz6+Wxyfm6qAn0RbPMA/UGMUfZVa8wOMFlHogXPJiZHl2mSConE
9SiyPGqawPLfZERagbeaOs+bxZy+czHoq8rFchKG3OHGA+AK78MvFplXQesepB3BD6u8iGgt2Cx6
KWFzMizHU0f/nwcpDpRdP3JOj8R+R+cy519eiZe7RiAYhcNImcGdu4Rz4nHUk6xslKur5jefuK0d
3iZpl2PL1ZHT85UXWzjtqmlEAkk/QMvC49SI5JS97b5K8u1Ykr9Am71mJcrllmMrqEvSsoELZFte
ToIPoE36Exa2YRt/4HlbPDYfZpFIvDD6mqunxrYVRv2bXAbRcANjrgRsU3R9+FXf4AygvqRHNiD0
Bk/KBcKpUY4L6bmXHtniTnz5rAz/tcAIgJgCG/QQ0A3BrWO25hpzo3wve+znin1jhuHyE6kQQt0v
5VWNLuFTmyT89vPrG2Qa8v/DNz1P8zFlpVfO9iSEE4mpQT0wZ/JUo7qCQWPqGtwu2+/PEARHxNWM
8lQy+dMQvrgqWacMm9kztO39iO4ajKhF57k0gAfRNx+ivRo8eRwRxuyihtWbFqDfaDwQFluSDQpq
PfsX9PXabdhIwKHT07zwi179wL8qDFMoFQ5tbFMbfReRh7frS41K0vtn6iudqyEEZqa/7UDBUJUD
JqL02dRD8pzwyXTxt8pN4mNsPaPIwQh3xIaWs+z0eXMcEZFPn5OIyXB6QIXDYKIV3h/6reOOB/qc
DCK2Qz9dHpBzOOmYCiCd2odjQb7xFam13UWi36c+lnC6K97MMa454rUkyV8Ig3VX/gWzF9fTZAai
Nn1cwz36wPMUWX6W8oMyu0kOxn2+TlbWai+It/+b7U1stp6r6vHUH+vndXdTLaigL0TlzzxCDfqJ
VsisppiSQVOyoEeGIMkhFwNVRKY5Rkb7SiN66O2vSmbui52MSHw2ovbk7Jy7L7xte0GtnCYIoeIW
EwScFE4WSZjweXLhG6ok2zbFfDNyWTQfTtGq0/QcN2FpRNGjSgH2aXY9SIvd2P2JUHe9U51YMPMh
Jxjl8Pbi0iF8YSoktrR5Y22mwGs81zkjs1fgP544YKWu/iVcUYBtOfJ7akyqIwTUl+kiEKpMmwVR
4r2wbs4ovhjzsA82flP0W48S9cEi7fhRTgesmGOr4moTgmfQsc0JaOXZFYmjnNFQT6/uEmpKN8c+
7fxe+vEcPGiN+Me5VqV283yL3k7FWDy5C61FgYSbfq9VyaVj3ZvhEAYSsW2FszDTTkzHU4c+T6ns
neWKw1MivebTLFp6Zb6dFAjRVqbZGebgFDWVTuluOc8EEpGMYqjKq2eNRXq80m3JoVcH+Gca6btn
Gyd0WhNFOgLsCSf46bqzKyQPJAtz47tONrdOv1LUMPU6FbNEm1C/Cu+vfDjqCNWXJebb7hVN7Nxx
2FhPVjUdEj6Iutj20v/g2ZzFaYJnKRux/XlSmLFRfkZBhTT9hP19dnA6myMn+zf8dSzoezs8uh9J
cx8Dk2MDOdXYYnrhxy3tDzMTSArKr01RuP3w/JVVsyJ2gkYJcPnsjH+uz4uIqkIA4a72y9hp1RCh
dhT99g5avqYcWanWzSJBOw9kuU9dIB/mWMCFkJX04vBMkGkNhMKL4evqxf4TBSBcehYLn8z/QlDw
0nGJYtm/VudFeM4R74WrxDAkvMnWOKLYiTh8zKWOhwdgoD0bM3vvY1ykuca/+zqZLzEceaA90OZb
TdnxvXUR/FVWRI3ffmZiHuhpHIuKnIeZNSMA/OwcrXqCPCNmu13IJhOnqCgcUYEaxxOeoS2sR1gm
TEgY3O4nrVWytOCR4xJV2ro40yO6JUXUwX7gfTSG08Q3AGETvGZ/BzT4ScNnn6ud8R+ZF+i8y94l
rUM7oL1tun6+9R34NDXUL3k97kR47Wh/IUrMWjMR/5pbWOx9RULQK9PKvdDuRBlRrXmLj8hm9XM+
LKMp3BGjCL8qPGPlEVG6rLwnc8Gs9tKb0WK7EEzmqX15LbNWSuWmIj4L1/ekwvzZPeUshYA8onr3
FsTvNAh6DBZXiBTo3aXPEzjhrFEZC3XjfdKp0BglWVBShpO890BG9IOjt5GT3+8J617fQNY62iUV
XdGF6K6CV4PMQzasbFLAflyLCSxtvu1MCpz910ZBfGbrNhMMyuICx1MlVFigiqj1T8iYKc5an7L7
gl5Y38RD0rY5hDmj1rwxVlYmMwMW4LfI2F2f+IMw7mUYLKUgRsbXBVeFGpVPicmkeB7oRZbuOUu+
0jq/j0sMq4yGLo5XLMX5YxdsRMpU+vYyOblQ9aVw5VWSlOLme5cG4Jrc2f/EasBr4M7RfhmNVp6P
yHpjj2N6sLNzWHHhoms4CJT6xQywc65O+yaAvtnRyMhMqp8eA0Lk42w2/zy6AgRwKaSEMqLjtZP8
bgo8oSFQCkwR3omannt0KtX+FTSJy/4DoK6qqNrnXADdvSQlLwffOsukCgTVUtdcl0xDywlg+pJy
sjhzzOnXEIC4FnfXdF1xkqD50/07MRag2hyfGXUHxw/1jvTAEM+4KzlfRJ9fizSi6ymKUusBsFOq
CN88mRZvoDJQ9Ns+zlvdVAPojfCWpoIZ+E9YyHBlNfRbFWRhMTzwuafhgW0YIaUKbrvAf+s2TtMz
P5U0CtfWPwWxf4IU+luZZx96Hrdql8+94jmuORjJzPhEORf4GDjkgUoTFyMH6vos2Fk0yFovnkfR
4SnUVCmxUV21rppiQn0Kc4ZO5E5hf0ApQs73IJgplU/jXdcjXF7gYLkFh1cAHmeJN3xO1FwiPajo
gysrMGUilR44MORMIlpR0vXWEWycHnjkty4cI9H/KBVIpB2PG5EQ3RmWIoH7bkcazjY/JINSbvN7
yTF96UzhHjtwsnKUYjHsxPWd3PJzpVzISCM/Qu1zf1eHlNG6xPhLwjhyP+U6a3CpFrtq87TNcCoS
0qXVclvrGANlFMeCSG//RUAVGYyNuZQv308HxGcFY3DrafURNKcM6jPYCP1VHAkqnEpL1jvmFb6X
TnhTh7KzkIPIlnD4JI5F55meZk+5QIhKIfpOGHRD1jua0cotvA7JZqxaTd0SQ6iecfCicm2w8jBv
aYRVqKKs3Q0YTq6uixxHXiygJHq4HgiLfg39CRZABZeRplPX4vTBsbm/j99o1prf65TufkbmfWi7
8V6zacLnyIWG9N4QNlR+VjnR3gkZGdTVL3vDoWEHLmz0X0ooTswWMUUXLNlTWqNMltUWJvRG+bI4
6hsq/azJjDameHG6dFlI1imdYucYzV1V/SappOouDbhrG5YL3FItdkfhsyZH76fI4CLHO9VHOl5q
flCcCHXqPZvsxia6foY8DYAFtc9XHNzI5T9qyUZSBDyHz3KN4z0VAtNpERobYayRQI06unUQnZfa
6yra3CL0OA82u5KpU8gj7Xo4WNTv2s1ERCoBB3viVlspDDwfQtb0494Ia09bv4Ns5CxPGHzdQxd7
O7t0S1mn0fZlR5uJd2rPW9PeaK+nDY3BLr/3nukE09NHetKtGouIGT21pf1RK/bRriP1sAI+IEx2
JECiMKKV8wz3xj65CFZO7lW6EY8Oylz3+VJOaA+rZKmyOxv9J5Gj556vaW+P6BU9WidacXYCM+h5
jXhmlPc8DH5S5omEgB96bpJPMxIS71AubUamDKmuNg2f+xXuFRpMs59oLtcA9NyRRebwCrsbhJfj
wQz7FiCwkfYEwqk9Yh26SdqL1pwhwqvkj2jfnNvWMFldvzAv9bLuvJm+ziip+19QvMnpjmIL8hUy
6JyYlBJrIDFbhq+opcjblDoyW/8sbsjslh439+pTovChvggxepcj9vbfvXU4UkE3aHHq74qVcSsy
/BHlASs06UeQr0mjvw2p+Fdeosp7W18QLtEWxTLc912wiNWcyVmk31EXtwQNyxR8Lq3sVefYDaMC
sHqpqDfdZhoZUdgM4Q9wL4XbcRuVxjox2DDOPPXBeihMw7NN9VGbrwIl9Hq4pj+CI4WDkpIZ4NFn
mRmjHtynhTA6XZdTylN8gSqrcrSt0iEUZSAp3defAunp0Vwba9+oqOyWWx5Zpc2jjTvTq/b0xMcr
iYeAfCkRyeuNXjoZp6sk+/Zs73m5y2ySqRT0cbph7D5f0VyJeg9Xq5yhoWR+xFrJwQEZ/qphD6Y3
WqWcmDjHB8MMn/CwIQMJP3fuKZaUPL3DzZJfHXWuJU3G1hINHLvcgMY+by2L6j4vBF4JNEk8xbbf
rA5s82sBMqOWtCmdtzAxe2k8t7T2KInGVzzacmfeeE7gtO0zrG5K01bMT0Tjz9b0L+9nuTCU8QI8
tNFnZGNrYNHvvDPcRMHQ6c8VtgRhlqX6Jvsb3Ju2J8g6wwbLUeFxL2fcnxoRTiBz9jSgvh5woC2C
4Je61atrl7f8BDpdJ3xpFyo3+m2927lnhlMrHnJl0d3Khd7NDf7zIEdb9SF4k1vkyefHLkeCY0M9
Q8nOHg/cqNLDzEdgSuW+tNDV30chUQQmBrvCZuesYi2mHvVBnnhgUxsJKV2XH2Skl9ENTva3x+qK
DTFBKgIzoRuQVitJ2w0TSte92zYnR8VLyss+ORjm3hTQX9O170FCThyZzhZG6Bwhv6Z3ISRs2mzf
BNma/2nywoVDTWE0S4glbaromQfGAERtWLhMdTn09QWMV0KAlUgMHI8NLErxDnQ71OS/6MVSqA9S
dc08jq8Vx+P8stXCTMHOGpl74vKFcGNU/gqyshjJB2IHyGS7nuvjLK6izNT/XPQ+jWhYJMoSA+4g
uZExg1Gsddj8LufFfEhb5jsbMLj8hBEt23/8txayx/7qhQdf6HNiDmBm8vj293+CdTtXs3sOleoc
94+ha+SCLnje+ZMQcuqvVYANDNZJ5zLt+97ESluGkzFdpLj4KZhrn7limzMgelXvcJbmQqznN2Zn
luSP5p2yee5lgz3spVLCtuWehRIL+lYQaPOSrTURtAlG1g46drhy68J2R/au92UjplfwsfTkNRUp
ysEx+l44ZYykHemMDqNQ8R0f17jlgxb1MboODSIQFFUBB4M9ap/SrDa0d9KPho8q91ZWa5jOSt+A
ESGZrcPjEyqG7D1qY8Hi4FRyicMdSCF9UXQWaZPHRNESM4P41n5OGugIOllXgRR0jn8XSbSN+EYT
vAXRQ1ZD24cRbPM8aSRRZdqVB6kS6W3wmCoBG/R68pynTu1NLLLSkhUlp0cfoxxzkuq+KenHCMlu
ykEQfZpjfL5XIiHZKmjDWnwu+fQeS22URhxnFljiIM09zMHvCSeUQ9gUZpRjb6PTJfDIACusHaXT
8E5W4HG26IZ2xP3Y7zcN7dSgYphj/4NDlSVkCSTw32l6TQJDAfiFhRQjaiPRtwhjmLA2VfnOGCs+
9lLXJbvia6apVb0eUBx9xU8i9PKSl6hAzwQ5uWdeLY5h78DtJWWpkUI3bmBinUkXcK8yXwFlFvu6
SLvqJN1IhaBKwITgLWJuOfFuVUW0a34cuJ5UdkQx/6h8KJjP3NtZXtPWQtZmbZL2JAyfeDnz4e9+
r4IsaDH1npWq7xDHHvFOqMP6G/WSbntPpk+mLyqG/0ZeuPD1GgGloM/OCPY+34AEGRef9Fd5SIz/
LhuriNYda0akoN/VLPPh4rKaXLyGhPxhEc48DI8F6G234c4Lwi6agRUC/ruWaxNod4OSyX52IxG5
QbIb1YyzCuIYwavaOC7IgNP0XXWk7ddkgNPzCklBa+1QWNYNDurnD3MqNprFismmPXcRSdNeuLkE
Tj38Txy1Bliz5iWODg7fbBQ484oCTZ+PJcaknFSgKYttroYGVke9eH+vPMESN22g69z/v2T8eyii
GjypgGI4cyHWViCL3xEa/LP3uyfqgXxGhuclTs2e99vFYpRj8wOvfWfRjqMZVl0xlcFVGBgv018X
/Xf1XscXGyuQdbNtOpPPACLX/nxRRienn1MUuTOnrHPnAGLJMdiK5q43m7629kh7OF4UZ2zwfK1U
aXYp9Lp5yHrEsnsTEox4KuJwsvbY1+Smv+V71IoIdBVL6k+b9RUEm9LgVy29RqtSl3E2koiaKlnX
e9fyKvHwf+dvR7Z24i11Yc7x05PPbOJYP9SYnotEZr9NnCca0iCWY+/1wCeffXDdEuB0uGwXI4Xu
XtI45udmBSh74asYbONM1+eqYkYIFAZeyiOe/urWUvCHttR2dh+Zisqp/FsOJgHji6EvQFpRDBIP
yE6/6IKj7A2Fz/aaeAg0XQnIiiDYkY0aSID7dy0euFKwtvL840Vv3ijv3Ykwrrt/xpDJpfQ21LIW
kMiV63p/Df9NmCIy5nq7L60U5+nuCuYAIlZIOOMOrG6tB0huxC2C80NioUK3oo/FrJQU2zvgK4v6
qALn+kZuSOczOCL3xca7HRvb/hUWEs1MVl6FHIMHhC2PNK1xyQT+WTd8e1Lvu3m0EmWQHOPYfTbd
5GJDtGilYK+lRj4GLEjLA4om69Wide3RvuKzAMZhHuV7BG4wBmh0WXURR2StO4zHI98BVQNJcfRI
jnn708aeWiTS5kHHe1QloSptzU1i1628914TseRya+fkRjSUKH/+ys3v3nyEaICdfpgFw1w6yFBF
fjpw4El4DPasXzqAUzY797U/Lq9nUOc7Pftw+VQ+lr7lnu8rHEHAPSwehQxmKzocC0EgxbvZSmfy
a0+6VCcQYyqTwrMMnpdz/rkwwQ6Vo90M2eS7zUW0DhhAqYl1VzyYUp3qoaKFDywJVbxjUzxJ4Pi9
V+J8POS4vRHya+m6NgjiHioqsDoBNleLtZcbXybbqGfeSeiKeKKZOUlhnYysEDunBbgSrwWkd5kX
iWTzMYGh5TIe8CwvgLOENCOkjy3ZGoxaZcYuTpX5MOEL3Rd/pwluaOISMif90XFXQnnwmgVyKoN9
GX40PDER9nxlsGlJp6yK2I4QlqLg69OtMrVBw6SRva8zJpdJRFGCSGOG1x6NR92Rt35XVzvk5xQ8
30btvchhaXjsop7b4rONGHiMyHQmUsy05RGeNkl2X21Mty3KVG/S8TdPP0Lzn8iUvDIlje3jzoCR
EGYd4UEm0WJtdDC/nrXJE+eh+9xsInemzOAxG9kks74/FMfvDjpEwh4pXmlkHPBget+pbyNKhTEz
p+qfn91FsMGOLCJmqyzQWgKa+lXyGd7EBh+OGnNor0Fb8uB4MvUyM523Edi4/y8fm7OiTXSZ9aXn
lMnlZ5imWZmsCloBv+eOfKWa8rHu7G4NlUoLV464ECJhaHYQzjIl3ZzY8eZskmVUF9qQjQJDJrdg
Dule8g8PBsK115RaOa+Gy1J0GkpnZWS/eFJBtmL9GGPK3XcHR2TdIdE5cBX8L6ZLps/x+kb95M9E
h6ypIqMEoCM+YB16b6xwFwWEO4vbNyqbifiwVrzCor66w40Z2al1D/7dXQkzBfFLra6P5Cx5ekKQ
Ep/UlkMYbHkGPAisEEmyxwA4pQlHeTF6sqeDzYA26Q5SxYKDkakcOmiA0k/cU4N8WAz+T2Pohsz7
KYqF5DuL1o7DNhvgYlqvE7LfoKiOFOTVH+K0+X52JoYHo9t+6w3HQ2DLIKXiW7LrPcpwLK/7Jhwj
DJK/2TcJXFNOMtzsrpkoMSK+GZHptITJM4Bhu5Ow3ZAu8otNd6xcTPcOMxOhV90PN4wZxJ8VsNAb
ole6g6CpKS3SM2GpsosvfMXNxt1pcSYoXEt1EwSbox2HP4BXuxmU1eMHGdaZGD/jea3YBHofNMaC
vyGeMIyzqSYWo5zYrg/AelEqbeEcYaCWzoG+ZEueAWIaAeuwq6vBHuv+G9iuzJSDT2TFrB/Lwa0w
Xeo5kRMafcFZVn0VNHmpQ16STjKWm4c4EoJV7OAuj/mbhXSM3ITqw5tYjOXpvvY0itIdng5DGPrW
RLIwwEOkvhxIXO1NY9lC3E1xVx2igr925QPZHgn9z1If0IllKrmEMF0SUtd2g9fpMgaYYvxaTcTl
ZcrUOKkMbjA8ttCQwEqBj9pktqY9Bx6LSUnRkmjIcFfEaLWWapKNJPsyyXXM8eA4uPzrWFu3KhGl
dD34Lny7F0n7HEKimyv9HhPYZqgQGnsXuHYK2psLDb4/IJtmWT4BMy00OjBrIpMgUQiwCVS9ZV/B
KrBTg8G+GFFOnoFQSqqPBRq5dT7qv+Y2BVxClm1nXfODJStD0NkS/444paYbZg/Qv6NICmoJJIc5
6dLVhHAdnV5HULBoe3G9BQlId1OxjGz3tJAj7CVI60VPUqmIHSlJLUwr6gU+bNCtvwd4J+LSF83T
o3WTtC/Pg2Q87kKe70IwZlvtNV/Qb2xyOmsFTI4AdG6EnMR0/CdvrGkgoIDCLx2oC5EePqir+jwA
3YNYPrHiiWHq284uWekl2aC2s7/pXOQ6Und0jb1q7XRz21z3KbB/gbgtBhjZtWByJn1mLJQS9B4t
o+etToIP295T7yR6WQE5qTKXqy9ioAEDSvLg+oIFcqq8tD1w0RtR7lN4u84PhUy3ps8qc6jvs8JR
W7QQAy3IFMMPeJNG1bUwE1FPxTivFINbX33ENPk6d47kA9X6HEbuBRdL+DkTYR0GrbCEoKpoPUgu
8CQNyJOCAhd2Qoo0W26Q6g2twx+XYp0XjzxXtjVG1YfC0lcgJZYkq1aAOjhZwRBTb4m5BXium/5a
DoyudDK21Jt4pqOPTPySH7Tl0c5jJ3/Ps25wMGBG8cAfj7eGGnLVLA6zR1hh1Z/sQxTDM9L5Ahub
3FlgNLC0QpObY57KVdpap3lJiMcZ0NiJmx6/Xd1lsZxxjdEvT/C5KEVpBQHyvyoutmqCkVqaMP1K
PW9AaWSOduKXNWppRSdsg7RGBFLVKdaEgQPQKf4S0vPpnxRb9uUe3dPnnKZTFaF6f1eddyUTDPgz
Y/kymT1skP/fakSilvxpHkElqCSczM5E+8sFgWuV+/qcVv8z5DSDyOJ3zDuXKqvb4Dnvhnq9OoUN
PO7hL/9RcxfaYLR4CfGkyGhjkvbL4j/qCimyQGuFSwAL6O3MuR6SumY/u025PNVabRlw1ld9yHSX
sv3zyVsj5U9ZJkVUpPc5v/jqHbl8xSEEjTk6ZFIUZPBaph6xQ1xLMkjtvzWqoorZn8B4AHFrZJ5p
tQWKHe48EnpK1Ci2mjNauWhJwdqlO7LLJbIPEuf0IzO3AVVo2pA2Fg8mfx5s6bzOrS1eTrsBWwHi
+eJKTu8fQXxVuLKLAnT7oordEyrocFawxoOMZM+cqSe3PJExcAYjE8a6Q04qNu4H18iN3E69lcdc
ocPAhf9p24X/XTA6TASzbEzRY3OA7QdE2qSAiYp5SLnZvPS/kYo2gPfNR4bYLTYM8r/vvbh27IH7
f4BBOsg1RJPhEVTO0P549wXwOsRyY9LM7ZKNCJZQzunHOu0fXfHljbzPyekF+PVSfNwmKKHx2QVC
PJJ7Fsv5Xg1bkfjkW3DFTSKMnchUd2s9s1kLmTPuOCNO3aJg5zANRYNfPHvVgkpWxq3Y8sL4Vcdo
w8EEdEP/eXasfkWcle6m9I9OdrM+AzJEdthHxYxeJkNnreYpOYNuP3R954FNw5q3VL9xDjBa/Jju
e+eEuErMF3TVW+zkNe2J6UOEtVBHVH9hnL0J7gWhB15kZ6ox/CKmz/sxWjq5EFeytTfxnC/qBCBO
47gbjEnXNBEnUWYk46pOYtfQjaoxNqrl+//4DTnIcIMsTB1Nl8wyTKLlUDGv6+b3f6lsYPl1vF59
I9JvgWK+AgaatlxS/2NoGjGW5Hi+x8n0ft1eIRiF3JX+eaglAoasr3s3C7/76gwvG8t/s+3lEfio
bZcaEmBBt+EDPsEGVWEnlfljTtiQ7VYFLLesT+tzw5YJP8K7a4vTQDeFlFHVZCO0MsPvkR+pOCYw
oBYAmNSXeXiW73uKG9juauvVGE2tch5KyALHD1Km4PtKetkso/q2PFvP7Eh3Ai3buxNDEfI85Fzd
3Ai38a+rXYx2XgWL4/T6nJBlPQukJ1oALSXT2NBXkvuI93hyzMxOgM2/MZZYK94E2PByBkFew4+K
Y3ZOAEXLHQRhY8qNjA/SoUAveyT411pxpNlZ63EOAK3c9m0qMRhYQpgabXyI/O3fsTaGUHayGiYj
GLiQmXO+wGN5cIyFD6PX2JPZR55bZdiigtBVCB9nWkxw7+2SikMysBu9pYXce3f03nK2Cha4joZV
S6POcOk5NgUBXBP4lXpU65dCipdWygZ32Nw3zOIaz/JK7cTf6ljkzAKC0xSQm4h+kD40zi4RcT6H
uyjXqM4hgzPMEAGl+LPTvPudgdr0cQSlNJddHFXekIvmGoLi6/Znv6qvJn/dcthfkoUXwPZUj2Yg
5iWEpDUjPfs7TLHVbQ27xSNVcbrekcMmPaRNwEV5LKEiv45aOXbCS5OcDoFaDsUGCUv588EGnJ6w
grzrDCT60vm1c8Ws+fN3rRi8omcTrdk4ShEv0B36Tfd8PgRJc1TbGMLpCfrfGZKwc4OJ7Zxbcr76
3eO/iTwdoeF9epTTzI8kGFbSy9gQhtOinLLdHnevoKDxPY+jcHqERBKj/GYJY8Me1gQtkHMr/aJB
bBSHr8x9FfE8VcZKpNpbcWcakJYevm6poqInBQ/54fkYwVZ+6G8I5lweIjFptyoUq/9YD6C0PYD4
DjCZ8fXZPNnXpaXafKav5amXA3Ec1poCnOeiVvMR8RexQaXr1rQPWAaxFjtoDvjAJrH4SvGxVqdm
n02z2O3cc/vA6tL8Dn3p2z8vyXP7TqnOFv3KwoXBoFVbULfXyC9tDCQHhDJHuvWOeWh5hN32edr4
Aomk36MxMHXh0lD2N3LUVh77Upbdmu79OVKfFf15LOWPcUpxz9NV4/mvoHZEkdBuOzf6BZN2j+eB
ZBXJzcaPTKwTv3iHmZeD/xgl8hxXwIP/DbVmyglu1+aGK1wq8Vpp5tL2C1SSV8GGAR3xWpxqdskO
1AFOoEeE1M39U6YQ7Dh7jtRKBhAsDn7qUF7xxT4ngkBeXQwLcurpM+KMETFPogApWUUWhsDLY68v
JhHTewAkOEJ3a93xWrKhN8IGuz9RlcHJzUuCf+tYKlXNt4HmzgZ6TWg8YEng7TSscGX5bQsL0FdG
b/bPPzhv/O/BKeldsS5moYTjREjChdYzL+a+o7xyuC6sH/TV7xxBITHpwbyuj8v0EV6uGK56AzNy
wr97Xz+QZCbj6fpg3AtXl+fZaS3WDhcJlHy37KK5Qd4yHdzQyIZOq5PJstRfJhLPVjZSlujFNwXK
l4wbazB11YILk0QPT4lzvMJqIOOkjKH0bOJIf26WXsbvhLQ4+aKAGHwtQN10vpdgcKJYAWl4qOks
Ac5y1aox1XiNsU6lr6nc0r6dApC/rfh4pncNh0sXCt3Zbjbs3M/KbWIxxEPJbwOAxp3GWqlZv0lH
ht2W1wlARiAAIOY32HVRUJA4yliKE18DDG3ATIPBrs+0LBuArDl7v/lBrT3psNa7oATqlgYdLNyF
bPL6iQZs4OeOPABFx5HAqEbPzWlK5KM1G77FSzhaSvcpTgfh6xAcLJG0DCqpamRQ0l9s8ZWxJEVI
m+VWGzA7IBMsYM+HCybmAql9IvcBWubGdLDbMO19Wb1kcMUdNR6TdUwISwXUrgVSNUfdHcfw7bht
BQZFl6Sc7ygh6EYlYIFQFYNyMFwQ5EAm98KgTBfK00GEhRSvuwIE5D0pkGyis03mk+zDbsRRJPH3
UFHyJ43BdRkHkYLNUV0KwLHqMRSnjD5aWHEiCo/bD2ddbZlrklikWm95VT32I6DHxGY3jzqc2+wK
zagQdlYro63bV/LfXphnRG2Vcb2VsHHPicAjQs5jZVq9ST36ssodufwid1YQO9F55S7q4wc04O4O
wN2TszbLjko6ag3+6nz3f4lR2pn6PLngYEbo9oOOMBRiHD6k1rVMebfNTT6pwn/pzrA2V9i/YYob
Zw98/hBGC89+CEIKDejQr5GLQ+gBhmGkB54lEZYmdd1BrWf+IwjhCXgGP3APdBalR6lXBHGL90su
lXc3xZwwzOjaPCvT3BL9IiMsh/pN1Yg3Lf2FnGR3zAkCDooOYUZOZvDBD0/hgL0zpOX6mVYFpX1W
ogdbeT6vsERboYMef7uS2CvkCb33mG/BNIKi8UkqndsebCmNPFegT/EDbJ2rDk+bfsE2Kvl9zvDA
G2piiA5ifQtaFOLkEFnooyOI53cdNePKQ93/ldw5/axX12Kz//Y2Zf1BVob3biCkWE/y9xZWfNTu
BsX3LEZzYur1txA4JFkgHTnANrkC5XiTCGwPsy6J2yPoWI9IbQFfQ2f99Biv0WxyOcnHN+wXDEyK
/+M2bqrNoh+NiBpk9/zI3FVZcJliBkFf8JCqq516fuhHbeYRDH8Xvge5zk++4SGS9KEPVqURcPLf
0f+fYQU3pJmh4Gat3ol957r3RmU6PIO3BqLR691vO4f4iE9qeZyYaexf20FOXaoXlypRxXUwfIwo
ciPkIHhgcWh9mWHaPV/xNmgXx477ExwA6Xr8Q0gGS+nHfptvnvUws46pGeHyAauvtsKGXGgW8a7+
/EM8cEuZ5HRS8ItVbV3OvUI2mak6SU0W8Ous9jM4W+vSq1D7TLjd3as3z4vP+7mjTtWBLXZSgTGR
TN9Cd3XqwkJFqmGQ/nJkgzI4SJ/Z8WsoCMDwxlsPgYTaR+ulooiZATE1mYcmQDFtyraujdUe1JHI
l0CMzNW5V1S9RMNCeLMTZKEnSTk+CpsbC5jY0KXLjlzO7ia843OjcB4tCVAp+4E5OIt2WJiv67a1
l51OzTx2lks+XlGr2SqYZnWCE5g06Re95IbgYG9GrX/XMDq/VRybrOpAxkSnrdyCv1iX3cpcCfkK
aPZX1KuC9GR0TAn3/Hj+AaQa9Q1EtFs3S1EhetZL0WiYfNgcUgKm4t7TwHUBGncfpI60b5qik60q
/KLUCo6dZTCPA/yuZUTz0ZPuzjd5PCBjJLJeqmsGfpAe4UiVK91+g9c2a7VA51us8n+w7jqZ/7PA
iqXEQg19eAxicgsA2xczgSpSPNZjbJaTjk+Hk4crlW3435KwYxPefTmk8TMYzu/0SPV0S/1hmVAw
7dCUK2FhGn5HXclUtLCYps+5cWwZ3eCSdfNnqYDvIOm/YjzCAQMPn0askXThT4M1Re76onB/FLoB
0N5JuPGxZAbxnbUcURo3lpdG7x9j3ARuZROoT+ICHiMSrUg9OUPiR+vCfa6Falw7EziKdvn3Z8fB
eNYGh3OtsPjjy2B4TLLvpbncZ6dHKXSWvjS6ZYs6uSMrC3eN/B1sHPkfj6srObcv7RFV60DLbn/3
TAHrPF40uwtphaiWRCpp29MpnznlqNdzwz0vMEpRa1G8rYRBUTAAZOAq/t2c1g9S1qSRQw4ZC8XF
E1ZJ3mIomq752U0NnoAFyPZp7zchCmF0NBFzd8oTFqz6xw7GuYWT9RpZfcwLVq251ATxU5bwIjAW
cpCw8okCtnj/txl7xeXqFYkOiG+sHyusF6SoX+uLAIllsTdfd8Hr5ik3i+Zl2CvZxO+yjdsMwhV0
KA2sjO8mM+R0NYcS6Nw3Qy1r/L3vJcZaTIXyMKNEje42F7+CDRIj8Gv+h5+Y1EascFXnKuWUpf8a
SlPC7nPatsGJoEiTLsjlrCWQeeSjUrrg7uB0kxeRTHCpVU6Cy+QjUoNT1VoFtgoxQBN+AP6YjWEZ
OsWsQmdCW1lswD/NUIXoRzru5OxHkdnu9Lmpe8jdY0Om7xB8xwMFq7F3IsQ/PGTIjkxplqyVc3Bv
j9Jy0ef/SgamNEmnCNiAVo2/lB9Z4T3NDGfe9WsI1s2n3WWlPliyX+gMPKxWQs8ISV8+uKTMWDcg
ZwrxbWVqGqnq+8rIBFmjvYwR4QSJx+5grydZQkMBsuEN65UmEW6REJE0KryQNY3wz+BTZRJLLZW1
JvSsO3C6B0sQJxavgX5qAphw0xAQsltuhuz7f1zGGVaZzuPtbt+54KckaWeHg4h3/oZ+i/4WVuly
co5SSsXCd8NgnPl0kHUbLswhvz+uzoXKFkfG65/gY5O3sR56o4gHm1oUEaR53tpdn0AtHHfPdwcz
LTMOGswCjihp5wsEAv0msaAEOCOgGTugl39Jcooc3XT/CWoPqwMC624yKP+JUTRjuIPzBe+nMR9c
d/+6+4Y3gB1uboZ0bwr+ngeRP/XDRDHI0NMIWz8E7rWTFE8bkhrHsLXF1/vGCjOjNk8votmtXrSX
+oKSJ3Sj95b4EhkYKDO1jmH0W7T1JFBPEUCW9ZcK15c0530T4FD8R+3dCmdZLYs0EnVMFHqHrZxw
E/wqMayVtcTOMv0g481r3CYbusSi/znUZI/A/epCCiglYemcw6nvjqSEzcOTCii4RvK1zRPE1yrC
escab/xLFyXf1uJ82AZAd4EQQP/5t0LpEL3SULifdR31w5yeymYf7aJQBhdp1q+buGKFMBfy8hY5
v0WZ+U5jHIc6olvWQ7GbPXlgSIhIz/gBJLEx3PIzu3TC834lrwLJPKztW3bWLOQr9git+F5MgQ/B
TgUP9FhWwCrFf8obPmjGxBE/C++3eq8tO5E/6crItqNcVWZvU31PW7tC7qwCwWKy9ehQ/0GjOgD6
f3n+rH0vd2w1vs7oSeQnk8+IrGnV2a8oWsUcywDtU92JGeOqWhU8n2FZQS3qBV6e92RijtXuqdFb
1qrunlYVNvGtsSbOL82Od7H4t6ApDp8QlzhJGT6AV5qauHkLgpxMGtaMn+VuJzIsZNjHyBy+j/0N
eshGs5gos3TV3cdKy93l93A0jOkCnMC8HPBmsI7HO4wKGgBjL3grKrhp6GyyshkhE87kFbLle0VJ
4VY/taF0ECGjoVjN//NjESzNdV4lQBQ4bCcuHk36+3M8cszESfIXvX/pLvgmRQkwJmsuCtC7qRmJ
LhGRoO8SM119RbN7Lzn5Asz2Nn9A51T+5wrMgIxnCHaZRkGBTJA8pmFc7pff8lfiHjJmkvHRaRPT
aq5RSo/0MFFU/a3mjbd0b0GpjkPILdg25Tf1MbcPIDW0SWd/E46+BJG0gHTU0YUxc3yUHlR2k/X6
eA3mgCsT3iuPJhftWowVC8DnXvohXLgRO6kvGC+wQJLJyEmFWCjsX28E4xWSoKcyn9p+OGz9K0i4
Lc14eybNFPYlCrNHSh5T7oAtyo2Ouaqa/x9QpiH0Dp+o3wg6YuqlERwbppbpZqVUwCk/umcz1vbG
nOLbACUgES46KRvI6RH9uhJKjeG4PutUcOcr7EhullareLM6rAHsBKKt31PTWcpAiNUKWSs47l6n
0w2l4heYSBrr1Kau1WvbgXReZxoRMTHurNFN5olw0m/cql33DXNXK8wTYUdlGhhTIY/C2XhYgPw/
R4NL2WUAJFfnimxB/nRONDIIa2HFLW9BiX7Z0Odpij5fdBEmwe+vOhSIX8KrvF/PqZw2DYmcjbae
5DWwp8Um4o1HxDzF0xOpBDcSo3B0ZNS+nz8mXO+nh7dcE67Y7FScihBl+cAR8K45gbcLJ9xHl9k5
mXOXQ4IOL5oZb+JeHCV73dTaI/UVJx2f6ZgKMFjjeT+nAnM7eSrEtlB5AZ5kYTBqUP0BHYePgXKj
+7Yyv4rUDjU3QvlgeNt7PCR/yYz37AzxJQqL8iAMCLTb5sJUl+Ro9asqNQqTkC/Du7vMqKGuaIMA
oW2rvO2pw/cGqYTfgPIfdeP2EVxqP3dFlGSRmGGxT0xKtVWPqrm984tPPq+UiIaPNObehoi0ZoXx
vhLhDFhf+yBEJqyOVaVy4SqbmCtjmsRgFKqFQD+CJoeP2gEhpY9WE7Ve9/w+ISkXvUInV+7VvwNf
/Xy06Y/jPPJ4G2Apc03o5M082bz7kdMGtg0z3G3Skephlb2XwrKoYnnJBDFVTrJLUHn/jqlBRyLu
CMLFrkOIh/wlNsCkWXRr0YJUrKBA3+BZU2pxG7CW3z05bOSxPuICEfzgpXrmGoyCnCpapION5CKc
uYwCemvrGonWLbEcygu7ItjRMwEYHA01S2FFuTVw8LMxeyFkZdYfmgFNFxnge3M+rQdAqniagiRO
NDXHWu/Vca8BzoOKXs9jbSIYoGfwKMKSg6ESPAV11up/vXPrCBHNQOucA5DvGwXz6i9aCvMunyZe
wIF2M/TMqElukn1Nxs+eSo9kqwQqVJFiwsowHunimQ5XrbCOgUuphY0mJRC5Z9NCBVQH9Li0c29k
Pkem1nWz5j9ZNhw78Gvh8lhjGHGtjVcyWMeO2+iPEGUX++gzQwqdvUQYWuDUeJ6yQL7fLNR8vZ1B
IHVKF6z3b3mIVO9jBQX91frsQaj6cplyZBHBMWenKPs9iZZhap5YbP1CRvSvHhUJsThcweRWK2nx
yef27KLTZw43EVWdldzNGaWsSfmuJQHCV7duPE8MW4hZ+hH8gXMFGX5WGXT3nNPCNRTKKm0OUMcb
qcTORDiy+4h02Hlty+/DO60k+4Zpr6+eBU49m79IZsnpnCsUAi8B5xn1cVc3LJqr4kpzKdb/XBid
YF+At9VsEc3wSK+uVQuCBRoMuftCkLn1t9sVNt36RshkvjSkvuQFveFKSbZttSX7kCY9r+cq2gMC
52DDqCZW7FYgNMxo4igl+Ek66um0GH6sv8os270o2nxHNkHC3SPF3e476RIh6tFekxo2KTyY+kgI
1/ZQU+Wyv8zfj+rQrMQ1sd6MtD5xDfuly5tZy2heZ3aZ9P0hf9HMcdmE5Jrs8COQNZddRNZwrMBa
eJxqE7rQjckg8QjtaME99y5jWcZiWL1nMHXjeMTYNtAlr/kOvL3SY2J/+CyUGh3JTnN3mhi/t/pq
Aq6zMu4yvODIV5UM3Ln4YVqdH7tp2eSKQPorZlG223iTYDJc6JcQkmZVeHaf+lZgvb/KcyKnTOjB
XU7dMWlXdLkfEoK0ZQ5wQ56LJkVnPZuRuvYSqZDWI/69xyqFPNPeAKfppiEABK2WHZSn7iFzO1Bs
GDvXuXRTelZprjgA75XYf6QmLPQcPO2LrSFzTHik+kWUX4CLQ/GVZDl+/0FFdbQ+Z2+WZ8chxXoq
xHhhOb2Cuy2ba0QhcV9NkGChqPngdQkQQy0KxPRH/JOEvP3d7utACj1QR84potkCwjEm+s2jPI3g
ZvatJMw+AMd7Pq5LsP5IHcbiPrxDc9kQG6gvBXKjyTSaGGX1AGfXYO6RQ72nw45AOjvsV/2LyZfJ
oVgY5mgxk66snsQ3dOM5ad8pRhyvw31dLF3JFcPQ7YJeDOJIItDwruV4BV3+DhpUZf/IRIKwCUT0
kfvJD0NasrIDZwixC7nPLdLkzCLGkpOg7G5vOBLV6CNPBiuqyQdM+/KB5tNt0vFsiTRE/ayeGNf6
WSHkfC2JHwmgo9VxNn5ezqG/rr06XqxIVk3BjAMDs32l2L8THrN8J+WHME6KmLCJxJ8nQ6ACmJWR
CXTBuI/X6rN9tyHcwNDiBQr4xFgSh3edBw4iexwvgivTQBC1ofr3SA3GOqxvVs1XWx2K+Zu9udof
p9ClVn2DSQXd+wftHUca72ciy7fn0fw50Mk06Qwye5EKswHGKwAN8GJmQLQzUpuLwQVtGxe4PBRp
FSnuo5mjninQHCMWHNLDRbA+eBKvNn/PaRdVjQv6GkHIlMmF0MHZyUrvHuH3Y5CMbsxSM4jedghi
HxBPH9KT3luySsOdeWwNDIYsOlPDcbgngS8w8wBabCww0w6YaX9ztuKlOWBdGxTVFI0B3gYwaW/O
bOfQftxciDJYAipitSa7HjAZWhRsSlH5e6PEcv4yT6cN5q+GmYoQulms1MVac0vM4kadcWCzBhmH
Y5sGQZtt41g4Qp7VKg9f9YVDt3xZOXkp1iqTt6zANSmV/X3WdkE8+3BPYyaxMtWuhlW34dHGs8nV
TKUHozGdTW4U0Vz5SFr70/dOka7hFJ9GxY+wbndMxJeBCvLAYRkfIZCptXzj0idXDeO/xwaR5zfE
Wk+J+U2w8FwXk3rBusAhhptE4jKzRt0spSkyqGm6Jhje/khvnalnBCd3OKatE1Y3G/fK3/D7VFyv
4reGcZoMPSku0XyVygmjuQObc+vUAMGTnj8D/MNwrhF1U0na1TmC7K4hcLZNaFXPHN2ro3yqC4hX
+UP7f9THyYrgpa07JGGNGF23ClRtSoZ0pwKOUT9lh6/QLBt2I2J/7ZFgE3ShH8kgjywORcvmfqCk
n5XGKKxqU5ue81zRqK3mCQUS39O9hK97APbBEUTMw2SlqrLCaV7aLf+zcRXlkWN+eRmdHz8DgPDc
Scz0rkUTm7v3Ncc9MzrT2wc3OQOveVMj4GXWUgnKVshQ6UC1SxfbQssSSZ2jo85LxvFq96xy/TYQ
05P6l2/NC2Xv3Z72NSVGz+HKV12qrmuMfvO4SYYz73OgwTBekqw9Ry3yL32g55sbzDGO7jqw6jJ0
nIZvVOU6vBysYOX78eR0FmU7vMlCqhi8rns8l+UzQr3NkZmnCXNbhjeRMOFc5rwSTRXbJvbeW1aC
Perq3l1lakwceEcYsfM4TMRnOur6WCzI4evka3kDep/OEDd20eYzgu/wLVO84fwD/livpZGIX2W3
yUqdkkg6JC0n+KEVKLFP8ODtgCIkKiyye/Uk23598L1pzqySt8IxGJkf8CY/Vvf4Br5CGwyc9s00
2laUrYce9Rs7cY3zaNq+YaHLUJdyPiHdbdkHBIIb7Juw9rX5vq3Q0DK87ZNxTTOVCveNFHQaPJ8f
chtNEX1jvLqv9QvzEcrYTpfzohZ2rWpgD5abr4SNHEX8gotiroDEoC/fWmbFbicviwzvCqbObFeu
syayMD2c7xntyhPIJPf2zHZ5SuaEJhj3+sem/XCZSqU/vOG9VG6TFuXkMIsphwP0IsoKLYsnXdiX
qqzn2qPXKFytEuxybhIF+xjfLqtV7Gaa4XGyBJgTU0+/FH+pE22ZSGi0nUhgO7OsPzujWsmN9MD2
eUpcRbR2A0XDPgx1MKkK2PVNfjJ79KZFvpSNzSI3zattJeoCCsRPwbraA5dyQakS0hAvNMMXe+BS
+27ybwRhIOWrlfZa+QFM6aMCZTwWKpDN1saMl9W14PvLGMwb9BIF52094xTxbwYcGPgTM1G4nfxJ
CeFGgpXvE5s6W69skNVLUw9IIjmLDRo8c5cgnjsPicOu9xNZ7F2P1aTHAbsYqDhlqSsRmV8/ijHC
SBFZqb0LxmEVe2DFcF9D5KRvclp+r2CiCWBet3phOQYT9LqUbWiF3fgrocj5+jHwWx8+LOq1fFLV
7eJFpM16ObONg7G9iYsobxml9ASJ+aEYzfAB5wBPuucEGMggJNItJUfPESHj1nut8QbvMSi+cxw+
Dasciue22TRFfaFs9k2YM8kp2tRbeEk0IaMz+ZOn3fb6roVWaq3GFv5Dd/EbinfdB9JwSMrpY3lz
3fsRzif0SHU1+m0EGjVRbMPEEuf+8MXhm9VWoLoy1CanxXkUB/yhxhUzDZk/edLioT/QOSyAW2BP
G4/tPEPOhVtKTEF8XVjhGYQfdi7cT45FEjCbtPvCKeII0MfkTHWhA0+gqjCFSTzqqFNTpJ2tekjk
74WOF+cDcno8JnOZAgj+v9nOvE0O22EqsEwX72vawwjMm41pEl1ih/FxIHoHYkH2PuYi/Q+v/pEx
scnnTIFJu1+foR+7NuBaMhJjue6E2ilxm89O4q6ypcB/9AYB5BvykE6y0uc6lZjqQv3Mp6bdM8Ry
XOUsYQgMVUbc88gGWCYGHrB7KqL5Dh1wdqpjUv+c2rRNx4ERMiUN97oTuGGNfHbcIF+2h5yzp6xV
z+FljlZyV51nLi4tbQGf/Jl3qUKMoZSXZ1KbV4b2N1ERZBCLMaQtUClhhy7yWsbjBdKkzotJGviL
g948hV2GRgiXmdDPZ6dJz0qBle7Yw1b4A9z0DOp7DP4sMy5P/WrPHXucZ6Dbj3co30vrcrcsCa9Y
zpmkG4DaKHP7mrBFRtcfXbRQoJ4URIqoubfWrrgK2UtriOg/C1600actKbvSy3T/duObWOecvjaL
9u4IZqZH3OdeFZv+R0rxjkj0V1yw5MoGGTUr7ZAmJkhhQwFBvR7kTIO0KOmeEggUO8PsSzyPNJhn
ffEU6Q2Bp88PKR8mF+LHH1unAm3c90M5mn+ZuM4KsXYPy8KwV/lXxSE/+0hdEIWmWy20W6c1ATx4
+b6Ox/2fLBxt6oWltfYt6lEgmqI5EBFnbGHLYVP7/d2Ccxr44FlhRXR7JPqOppDOzpdRlDLIzUdr
4jbfBD3OMEXwGqY34Ia1/AMKBrqNO1RH67aTty+0P1YKJdWs8xAmRuVKMm8mvNHIVaPGIWbT3bUy
uza4j/dmLB2nMF+bGIRLx5rXN+B/9vIUrDxXbJ4n4E6l9k9ZFfle1J8Zl51ceyXxNBc42m+oV09C
7IJenERc3PwnJNo95RoSVRyC2PMO/D7e1d1A43PSKGZnS3QqxoJA4dndu+gxbJ+se2ytd8C0oGIi
xy4zzyOXzQs5+wIPVPK9xbe/uPxsETld83fbXoeZgAIcRWJ9NQbi5uhuCU+d86k1jUBaz4RLLMeZ
M8fPbKyfUbCyMd1Tu6JW5MqbykoEYyJd/UpTgCcyVbYRuzzrAIFKOhi+HXBdnOX9E+/MNm2os8My
BmRKrGst+Vxl3MBoBvGf/D1Jw89gaCvWZa0Y9q6EerCTSGGbxfVHsdRN7AjK7kHyNgGqfx1Zk4O3
U7zgmsFiakfS9GTphIoLFhHXAhzBYDCCBqKC3sF1ovlp8Yrx0Nb/gQbl7rKmFpezZx7A3xp+MPpn
CVYScHTofZfTd6MVIrIzHg4v2IPEcweYU1AOFCJk3qnDdc3Hcg5h7AnStH05lhiVGRqhMtOse0hJ
lRhhYdvFZO9Bvm8kSP46RIuywnwetIDwCyli1rHz6oLHSb38B6Br9ejW0en/JU3dIQCyu3wfJu4Z
YTlfD4k7uF/UtuTgWh3cwkkoJYipB4/B/UP8MxXdKQ9DsWc4hgaMvxq9c95uPuofjNCC9dv6J9OB
Rkr5zxe7LUr7FNfxU3/KH66LFoDQbDE7OzMGXzIpOI1OCww4pxgP7BGlG71fh7/kAd86C+pRcojR
tZ7t9zJVp4OSTxqWjjBXWyLI39B5k2BMZOqCVJvYbiD/k5qhrnULevLcy6BDYRreIfbPgaIKcm8Z
nrhPBz3EThcXxXRq2cU0EnhWNfddWIod40RoXwBJIlw61oGpY+CoSXU/oiGUcubkK4E0JYw8mGa0
ZGkmbBAmlfxh1pBX6gwq6ERopBHrlHjESTVyZEDGWa9cwnBIqNFqRcV1HGUNUxB76Nds/WCFmQrk
fzhLM+kJeX7J0heiPD+4BD72omkHBKj10+yiZUDv7brOOKp3xlgCUP+B0vkqrzRm/cA/dPevXsIf
R/ygvBO8rDHhLYrXOabXSOrvPkw6hILitQsqCS+OggZcyWQsiZNHqoY9/IakMexcJz2FLryvY6q1
1U/WmtIyw4rmmhKoP4FC+bYSUOZgMnzQa4NUTquieW2GkFWhJymtkwrCg/4pnhCVHASywlWcoDcr
30Edc60cAQ6xG1HmZ0SEIRgWmMs8noxZwoxuiOHQMyjims/CypNfTSrYsIJnHnbbCWfVTYOmsZNT
EwPTQX4Mv0x2kHCRvYncd7TH6VC69hCWRdeKxAJopVfxuIOrKntYhwakKYXXYjdYLe4zq1qW0bt+
S8rcyyIaYpzsD5z1YW8AVPbLOKYmhrCojB35lqQQ7QjXO/3vPNP8DI+nTwTas257IEttOfCmlwtM
tm3huTVybCR7psygzU/0s6kbQ8lrhz45FoFP76SW73ClB5OZoUNvcBT9DTCkRDnk2/40SVSEcudB
tPH0heTdeOkRzNg+qxeusx8mSiYrnF6OpfFw+YrLlxD8aHPXzq4/SKGie8eNQXKOQxUtR859aLn6
v7GYVu+bDaWXDgSJWw2eghnc734CgpkcMFjrpV9/WQQbuoF+q8DFQV8/8i725H8D8adUBX1WAg/G
W59JPXU9NFk2gEd2Ts7WZ86a2TzveGijWiMYXgFKQyAkUqCwiXkXqhFSaIHKI6AgljtiFQZrURtN
EnsH5UiMEAcEbNp3vWda9DYR6aXpOp/HGGHDBQffMMmyu9bR9oddp/2CNijwmACMCiHl2P9EoSK0
AZXgL8LZ6cBD7Ah9pnKLBrh486mgZ5NNvwS58HolJ67/AF59HPzRE+hkdtJ1PuFpjH8osL1Wl5UW
V7pMB9b8g1NIxEn1zf5qERrExXQmmwateAPIoY3xJax2UGsLEbsIXwEeHvOjNRd3QVs/EpO0EbsG
7j0icvFAgYjxPZx8Pezn56gmUrxIvkE30IPvsCTdgE1/JrYB0ke2mdLTT2vP4fG0Z3S5SYJGYAU4
2Ib0XTe75dfo6rOGlaS6QhZDONYIof/v+S2QWIn9Ee3dGSXzsr9NFtUi7deQHFlNaN8nK1BL6SU/
TYqLul37H8qzJsJKVF8qljwWdLLkJn8UUWCtZTKtRNtw1UQ2yMvXm98M3f4JQHZGgtkJV6Dq4Wav
m6XNdGtKRhfrng/zmKnvXnm7CbOgrtWzWrqUfh2bTw3jUwMPctC+HwOuq0+600HeaO0fC1KgcgbZ
04tK5v2x+gUtIPgq+WEOH+FE5/KEkQAZ4ieb5lALCpzNbYN1McZg6Es7u68w0RJGr0d6P9nLFBdp
R4fAY13pOsflwFnlQqX9NyT+uLwfIXy/LirQzvi0m7FKEdHoJByR9CNofUb67D/eDlJGBxk7v0ZP
Z/UMbBIssC/Ma5udQMmnkZNyIpLmTd1adt9L86o5cwlZh9X32d4qZ0wRqIwKDfpOtwt4izFSu7wW
Z24Y8GAf7c+87Clxa8jWcYtR1SgdjGr1EiXiB9Q6Ppp3WAasXWO1hEcrXT//9qiZi+OyLyH/SPCB
SS1boXB8cS2DzceaRx9xedOS8aJl6TCblotDBVp4+mz/tjBxrvW1Kd8TgZFjF/rEHn16FZlL3N3a
kl1vVRIHxk4BX0BWH6yVlpx8ozipJtlyD4D19Bc6BCMltOtlk/Ygw7WfihTDF0XbH8Qh9vKMmPm0
OlZUhtnQXw+jOkG8XvBp6yG8s8phSZDbsFCUhyPYVs8mihmrsxH48MAYgcQ+KzdAfNW4uEzOMIDZ
bFv70g7avrt2keU3SaiOZekv7UqiNVH64R35nFK4ZbPzN8ECvrVxrI7xlc2N47CNbegHcaNRMNMA
4E/oWdMAOxf6oNbNq1zCX+UVSFe9NU01Kpyiaa5esg0rbudcYj3YpQ1sG9uBzbfIbnZNCDDP6y1y
HDQNcjXQZEsLZSWzHDmLoyySouhJm5HZACGL1AfHj2zK6AdO9I5LXIGBNThrQyTBELuntSPaN8vS
mOIaVz8F4I6094kOaQTp89+tzx+PHcsopcxxD/b4SZ9rrFWjCitmDY1vjNMZzdFEOxzP02HBO0fl
Vf2+zznWcB6zEicyAz4a2t3TE5Th6am4VRm9CHm5scl503b4mOaW2KFPSgnbuWYPLAnGtt5Bxyty
eTYlBQtOYmitMztfsd3Zj6FaOTLdnMgX/qCnhKXUWIhuI1ZjmuNsvqSz+AdQiD75//oUXlJtwITb
KFKnOQ494iB6C2iMJ4QwHkMCfIg52rV/VCcrv/cD+zdTPw/OVDBXS6pCuM7Yb6V5hWzyjy2NDvOE
x0QvMZzpTDBWeHKvHgLVCt0Gu9gDz3hSVIrH5CMUxjWtSnluyGHHza3l8aqdtCsrgJn5/RqjJLFt
3icHs0KEgCRY1VOWHhXRRZzsAr5JgncLMuap9ojqUf2yugX0jTDYhIR7nomaETxI1fD5OVVCNx4y
c6GyLnpJloEjfNuAMWGWpQFR6lk5xI92E5hWZux4nWjTJFJqoJrHtcDb3rNmx41ERt9gXBL3eE7V
lA8xzQXue9+pxG9mR7+WdJ8QgKXI4gQ/ntSveNKlxaWOX+KHDQJaq+/1EHojy6ChDuDiG4qFKHvy
P0M9N9tNOeCimW29/KMN/yVUx4bIealg1Wvv/g0VXtoRKCpQEwwXaCIEJJyLkahZz8kwXWCsjFqP
U1HpBpUyetqWDW1hNcnyiwrNJobwx4G5h7ephrgV8atCIuCQDbSmPEX2iymTszHh3QAe/AHXuPFC
8PbsZO/tnkugDlWIJwv1y8im+PzBJKCM2HYqzpLUDvGUu/KO+2Gen/HJNbtH2B9pW3Bo52v4dcjm
QIlTDwwMJVMx/3EhcTLL8MUlj2yyQ5gSspl3VBW/uMxooBvds5WiGVfAhEbvnm4BuxMb2lSFeWaS
YqsSjr5ta97AUSZSqBNSSxUcNPN7WyOCR+ZnSiJnmW2HdA4E6bKjd7EQA/eUKCvFB/gjYEJUtdnF
horRAClZmgp228879jh0aMa/hzMztFZqNktgW2utkEegJqHeyhb9XflbLu/VKdh+HPwE8l/7jfwW
uqNj2p8byEL5MMk/lyV3nPlNtW5Q00VNhjs27m4AEGsqAox+i5sxdXMYBOqszm5Np5pypsl9fXlY
6xVA7x/Pwuewcdb7yHkZm+9AjDtN+hfxS3eGzo9sqFZwiQqwQLeIJMTcL4ddgnwCS3nt4Rya88Vo
xb6skDIexmHrdv5jehkK7Hit8hAJ25SCoVDCd/k+oMzKUxtCb1rnumm5oa3K2dCyezjak/sJxg8V
fSXk+bEd2bVJFTbSTp6E+ci6rBIEp+MXyxphkVOshKbIGZc51yCCRMJ04UOV5UwVPu8ThfB3QGwz
5Oo0XdvNbZsABhj6mdplZkdLJdiYFOINwVNTXo+EsEOs0uCayIQJSHHJ/AS4u+W4kPf2k09wuZy9
TCwQuyssM1JS9lVla6dhm6N4evcfQwrVAFnhklWPMIO5AZXitQP5r3KtfzrSmIfaX+vu/ov+nST1
W3PBvw3n7Wff2wPY7apEzcFPGaQ7OZ9gRRcnSnMDAZTkT+w3QTuRzQSTiT10bPMkGyIDsbj/taiQ
2cN0FeIUupf2jQA6o/8/imDDbwRhIx/xofUNZMqnDX2gm9lpE3uTivtFs7fVs7V+lH/AArZ1mBtQ
dMiGU55h7aSj+VN/BWz5LmlbZ5QzyOFybqwtKSTNgHbDpEdaZmRkcpIEPijrXRUnAoEv/mb5ca5q
Ka/6qMIXnMhT/IkYJP7+p5GMljQJyaFR1ViWBw5qL7yAthgC2MNyW8FyHZMvSfy+l0G2jz8Bcp0r
ZHMEAUvxxQS8U+gap1aZXEKSD5NxmIL0MRs6AGV2PXPiCIBRyb5UHg+oTNsagxAzAUb56/xdjgqT
V0dwG3A4twVsgY8zQ4GEXsmndTyX4jHmpekwkomitOuKAVoqhYVhRMuOMIqukC3g5L0nxuzro1ne
Vdeab7Db3A+Qy94OPAyoQjNmYXYT4UM26G640S7ru2/WCbbx3HEb7ZJr6XOmvSPitPz+NmFsDks+
CHp/wqS3usBuCE2knHA+LLiGAQslHtq8nyKgnAgE0rp+T4yzziaeWn5IF+qN1jaltTaat+FDDQ+G
rvWjjwJN10w4x22+Bw4GOd3MZj2t8sMJ+hVaWgpfJRvY5JBETijEb/8a6NtWsNITUhWssXNWUKtb
C37k5YQQCSgY6CaquHFm+XbvhaO1SzACxN51locyjxEowEFwRNAJFRh/Tku3pKcIO7pdUJztNMNe
iC8o6DPPQH2RlZW3vKZEtiAZnX93/xpfdOxNL/rmNELthLM4cva56m8dFChCjjibTuPEVYn6q4MQ
JNBJyY+bd7lPLzJ0pCIDYnQh1HhyPPWIRovZK+OBiNnseSZvYCn6yGzmTF4Mlzr8nmBe1NoK3xIb
leKCUV4L/H3Kk+mkv3gueHq/AONC+G7qvfpGuRaQM3jqU7Y++RiWqlemexAMMsAbdSG2ItNZl1L8
a8ZAQJSVkBe+82qyJW5d43a8OKx8eHb+VvCpRSuUt143wqXdGAgN1jlOFb9SGSBgsumOPSNQv7on
Bk2c1z0Urw8T6jNgcCaowxZuN7u7sDSJBpSe3PuueSH0JK+xdKpAf50Wb0HY570tfpEZlgi7iHwW
yodT++NestDROyvZbZbpo/o53UkhJ7H2WrVpAlhIOu/+IpLPcGIki7+U11tX90ouJAyWmJWpvMfM
x0uRhB4ZasTV1O+EAROhJ5FKmXW2HGDHUU1KJF2Y7xxxakqq9r2M57I+YnvmdsSSMLOAxhY7HXCt
I2Eh4vudO00CPOSHUcjHhKjhnEYKAWyoNfJ5T1600/RRy6zyKQA2MkGOOjPmUHKeIGazeisaOxw0
JM+FSrzVQxG7NV8kepJEB6im4xxJdzBA6tJshoFgFSwc7inR6Xi5z46u4AcH1HlsispKPUJ3SacY
ISC6wGyEVzgQzMAXusYVcBQE30LQHAMAF2+t93/n0SWk60wEFOSIozR1uTxj+G17r6MvAAWTO9eP
y4eoS2iWUL9I2kpnQ58ANMp4pXpIAuQqYm9C6ubEWuh/CApTAYMB8QBVlHWbc0sCgAs1Xi75af0K
5GbjlP/BALv1zGAzFEfwIpU+AF8J/fVBAbmY0ttPzW537Q+yLGpzqXFefwzMiZBikeap81NdVr4p
F2Vi3IqF+mqvkZu9X6NQ9cM+AG88rmxlpvKUG7JYVfbczgbeBZL6iDV6e6LZgA8ZpHZZHqWvTIZ2
wCH607KyrtrLC7SssKh0UiCy+LJcONdICJNfYhedTzWcwDJJOvxKvO6czHTXe2T5OgYAd0Ws5tvZ
qmrjzFPYtMpCocam+wkfIBdBWT8CVf1NpQp9qpfhRYGpFw8zK7L3eQUji7w2h5jHaMUvSYG+znCL
4sVzdAaGrGbus9dcJldJmFV3bAkM/SNMTRm+JaXJYcLmAjJacYsWpGlx4Equ/M3PD/wU1N0EUV95
8iDif3ghLpZeqzCeOjYWuJVOTm5uQ274FAY6WBWSqQW3o0LuMEbiivHCpkDZA8/2iQXd0q+yt/fv
FLqHqgZ1Sjy8a7TmQ9nhEhgKdighSivRlqU04S95rm+axzEHjeqYJDCy5csom9setb0GfT1evlJ/
Epkjr2jdir+TLc4/wa3/+3N3fcij86sXf7k7YrIepfOgw5lVB7aAiVztLzZR/Ok6mEaqmNRDVKMk
qlAz7eq8n/0QNIQRGbB5/DplFLje2HQUJiYQQ6QqCB4/xMc4da6kRDoNK84VZpV0Wr5NqPGP86IE
U9uPmOM9rwL7lI9Zp5ffV1tEjfY8PZ/LaQ8H/rtqM4YotLXwz80QbYWphmO06ZfgQmJsgR2/6R9x
m8LdbYJEUPWc+1P6zSXkUxXdHba7ArFLVdkWwM+RCM8768GgeDk1ganU8MizpALAWTkufyFaTur5
QeD3X3C+obfxY0pACS0sdoHVCZhmLiLqmXtQf9ydFB+28wgSupjSlu/XoSxAt4KxgqR+tQ7ATAmI
J/k1bl6RvVpsFw9/2Z9oXVIrD9YRXXqaRgOyygp0We8/b/V7wpo4YcKjaXMZw8zSfOM11QyFnXIw
z+7NtLk6Dn8jS2GXsz5BCmnIBrR7nk6CjUPL/3UDxynLRbXEqvTAI64p4J06BmhQuZi0z7SW9nlo
ZyXU9rwan7HzuLm5r8B1Jz9I7HTvUiwZ53NAymkToutlUxoIdvGaqAitOCw6yDbTpz3siy9nuFMx
Igbdl46wSY47rywZ6fZfTC84oeRVKI9oTviAdDlTV51ErVH+85UHSmEFOk9nrU2gDO76+R2en1Bb
tQ8+ZHrmXURsXE14PZ5eSBcvCVOuohQ9n5T/LltI5+CjATk2aU66/9xbG/Qtl62VDMSjk2Y20jk+
XbT7ScWRf+H98cpfU0AywvBKXUNM1LXPgFyfLIoOfueWMnNZT81NIoNkvNo+srmY97+9lWYueRWN
uVQ7vBcomCbWlGJFIhdQWA48kH9zz3+3I9DdaDSmtAC5JeAlaSVn5Sng5QEmRDh6fOQ/J74hwaZW
HyU9RDL1R5JKL78yc29UBFoXRvo2VqHCacplbIVjlPZtjuWqHXHdebDHsZ61M0NccxTPV6dXR8g0
W6jaC91hok+NTXuFC+z3H3HCNrhUVFYeO0RMnMuZlnevIQP9N/mTDDgHwnA3nUiF9N5VLx1mfiHh
w02ZT/6UtWwRB6vksNb7KJLm1DLrKA4aaIF8PbRuMdMBAfwapVBm8iym7TdqncjGIG+vpqD4SKQ+
nnDhv+9hpBSr4V+MnlMoEM1gIL1QGAx0JLTfsrpHU+8Q93TosVRanowyHXc/sSH2c7XnGYsOXklk
LLYcLCfIiNG/5DRQbYePylAquAv9S5/D3lDFSpUvAskqsBbTYR4LnBo3crFhs5NEZ/nVKuv1wsKx
h5Ogdz5rsBQXnnHkrpJ11HjfqYo9CO8DL92T6PlyymBgwm3MBI/9tAV8P8upzT7Ef/HPOLhSFExI
bCj+i2WzMe3cpLfsp+xlz7SpENLHoGSU5SeO/w2hn/l4tL4hTjg3/1R0BjPL3SW98i816fv/3+c5
l8zmQEY0/3EWV/gxsX1u1IQ21fM4t4ly7Q7o7q07oZY8W64wqKtXwXKuHYpKDO5T7jw2/RELnKWf
Br47ney/OF5agrKwTNextSU6481ftbUJlceSBqxZFyU/i0/RSQt2NAMUhafwsTzVd/R1/moqWJJ0
Y8rrG2gWfmvG4/FLqpTMBcsnaSgX7qzDURk1dUB605ZTQ2VQGAN2JnM1exoplQ/uVXqWfqZ+0xu8
pyLHkD+y+hKt9qcF5fFcFVGxHuAywbsDp+OM38QvyWYCm4EOb7k8jQI993DlGMfQu2G7wPlYCH+q
gwUHt1/6nrSneksZR0QBs/75W6kDPF16Zj7TuPByHaQCBXZjZeh4fox88Ml3psTtJsLtXUuWnRH2
vJWPiWiD1SetMayKbZgFS0T2otf1fTiMBn4HLirxcT2e/3yC34zxTRea12c8J/m5Cjz5Qds4qGNy
ehOu3tBdC5gFl/2mZieuqHWpo5F7tAUiLzjaPYi9ujvDkAmPNN6cm1IfbPXBLv4aAlvGBa0VOAbQ
JQSuP3k3rJz8khfh+7kjL1re+0ydJ1AB/eWxmMdb3wAMXWJM3aBZ/7AII4u5E51LXFnZaFAcR3eD
66pd7B3NqE8kzOHx3M09Dd7T8LyHoBYjfYE7Rxi92ImK/H89EwsV6Gbhll21KMl8y+J639PSULN4
a48xobBRmIp9wmCRP4y0GmDnDUZs+QslM8reWqBPqlDJ4Hss62mgv+cnMA1qsW7RHbfkynEM/DWh
bNuOfION72cbRnO5yBURtCnChsSreOdmrXdLYp92NbK+qb81LxkFax+rQKhlVuq/d3tXXgSY98mN
yrZr8r+rcaiG5BjbAZ+H3l3pe/JeD+RiEtqwp7A1QRhdmgF8ixYuWLOAk//YZC3up+GnoiDauPfX
P8aCtJ5uuhJMZLA5qzRuqd5+f360LxW/cgJolNXvxUS8fiYqYnf6uNIUrsGDqcJywjtyYBxGavtz
Vl30Vrn1zWoolEXB8LG+4+/hukOSMZbWbTbaOB4J1lVKK4cGkBGcVtKBwuKQd8gdg4jzH+XIkmv1
ebpt6BVBLptqBjP0omfpSo/dm42Sh58qv/mz4KxSJH1C3kxmPY5WTVPVNw6Y72OHkNuOfkLLQbO1
Wp3prhLGL9gnI+EF4zbZm2rXVQLenqqfuuOLGeibT7Q52t9OcbG/tJHrkvDuqVaZBCi/cdl8qeHC
DXmXEnJ3z2F3fRPlugoBQhhzlkknvRSRG66jO4SJd4Ge3wKBy2raRXzPETATsHcw6ptj2pCc9f3t
7hTs9h7AVOAGZ6xsLMzrOHbe4xCQgR4tJKBEBpfE8CM6vYmhExZCz7/A/T2adsiGq1cwc3nZeNH8
X6EgQvZUTvPraj2SdZhlv84YNsdvKtyDZn9zrQJtF8iBhbvz1oXDGgIvcR03PAHDbprywU0bOs98
MwlKHElEmmM+7xW8bxzr2D3T9jRbt31DpCZEIiX4B9MEkTh2XLXi78ab0HspAOZb0VnwmKa0TIDX
+2giAPWB8CJLZIENA0FipJiUQHzx8OtGiBVjOoxKtmp7nDprSm/fBpJjigSdfZ5E5ilNz0AiKSEO
3UlCxJdAMfznXK1MpOS5Gwg66sL94QdHVn3sehtFSm3OMBuWLxgrADSuaXAy8ZE6Aay9589/qlTA
PEAOIC123hozylgx/NxOE7J1mTnbERvBaS5cfx/TefRgAHULd/c37tOIqgELI61GiP/ERuvM+vBr
AxwzJAujUK6LnwQFecle+CT6QprNIN4KuWcfHcyju9illftQNdtKMTmMSPlmmhozoXzzibOw8l+1
q4t8PQdJBWXceASetEmkhPx4BZbXBsalHonfQUAQnD/ddszLVKL4c3WVxu235WYIqWE+WnhoFt1u
8iAfsB/02T+O5jXwcpVQhGc1eed3oyPYEgARsDyoUOvByl0HUP52H5XFqIgjdAPHQdHTC/9NnExS
jMc81veqmNYFiC0AmWU96B1fZ1sCb/LNYInqiO77TYDviJ057M8SYVAo9j3UP4zjKmLmkw0Hw9RA
HdkuH4t8Awb0+wfSVZpTtBs6mTQfHtV1MPbTumpQgSRmZrsMCYk/hVSA++nBFRcMi6CAgofhh4Q2
qszCJNZ2VyaAvS+Pou+jd04bjqnvBsjeXQyq3Lu0eLyEaz9PocNrKn0Xx9DZUjhzxS6NydfyUP/4
UDGxeMTGKKdLMUXb2zvls75oMcZlAA9zOnNvFW8PIkSTSU9GmDRHKjq4/3ZXEc1aBs046mEKJeAK
R4omw6sA5hlApk5UIN1VosUb/0naYeOPAP73ZRdG7tu1YyIMuWqZl4f5y/BYWufleUu7hd+7KxpH
tEHKEy1kgnjhuYghKGljrIQ4y/ww4KoXjxh6AiBgID8ubfkbO9pT7wsGwzff+xldbjCOkIHs/5NE
lViaqfQHkB2e9GyCfti8GWYRFnNnxvfv5NpNObsrioQxSfw8SCesnJm5NXgomtIbpckkmr5y4sjA
r6urxeXOA2bGOtinuw3QO7dbLXXOIUnzE3Kj+Ymdsy7qNjkG0kdIxlM50v+uUOUBNQEn3GwwUvAA
F6EncF76Kg2U72VJOkQqHZG9hT6ONAxEcOgiTdgr+TzpzClFxuZrGWfsfBwBgOpfyfmfObToa+8I
RwKRXr4zSeyNThNV5ZB35C1hpjuEelLEuoOyixbIfBqKJCNqdvLGyog5psm4t26Gctjtuxy91tiS
QB9kGCvHl+IYQC81okeS+mrwTZdrRR/tTPZncQ0oDtyABDa78BtZwKtqmqdgo4ExLH7PUfjjknNp
2ewxx1LwWufg8e6+OR5BW+A6DgBcMXjMpbFlwMlFRGxMXn9ElDBFBS91n8QZHkaqFZAkxK+Ufhgl
LAby0ut3L22ALkTi6YAwZQf92gdHhrhQISFLgRsJimSj6/1F9o2ZoR1Jc3WfM+DJMqullzWNVHac
voRYSzUjRepAzUdtvYTNtVrjmvy8yu+SOoiY7ySPr/svCu0xbaG9dzT7GOPQvQfNwOknYgR8UFpo
rpG54SY8pXrIIZM+8cj8gMVRK3aUuWjCWOByDkCcUqwCniP4JhlfoGVeMRlAaFcZfPhvuK859ksR
cCH1rPh5v0J80uIIMyaGsT/i3LH6KQr6/Wh0ZK4+vQnrj3Xrep0QZUcb0QWZV0+CnbrI8bXzyn5C
tCPGdifjNjvEcoobpQBINzM+9+MrS83a9mTsGelyhZxAs1G+MaedWWZDf6DndSgj6KlgfqBl8WPA
jbWE5Nq0Gv/LBZa344W1ydLxGiG/r7z69Hb0Zqgrigyz6042G+2nPgyqoCyYni6CC6vDtRfbNyeO
gtQnyqXUQqBIMvgnL1CILB4P8PScICHPk178PhMBf+uERK5gBpgPpm4qY+4Y3uSkjlb0Od+7wfb8
j/DHLUPZHribodZYxjNL8IuNoIoEChh6qRNs4lGcd4ULubseVTPaZisYpRCafbt13f0l88EWa4PU
cqdbFxXoPglzIoB/29D81g0FBQVuX95VLnd8DouGSq1xdMR99abKK93Xsc5lSb+Xvj7CQTlpX2oD
jhTkWtVq4Pi41UoD/hrwJHOrr1+eV8djM2m0lOvtfWAvHDaCjxczQLqsMe85Mp61J7HhwtD/F0T6
WkmLXgiihDe9jqWX3p3kmbNecXvg52PJKPL2m3jH4AMGW3BTv4UlpbD7Mw2HmQiwjAT7WR7Pw8FC
eugAARWdcFOOSQzGyApD6pkx71zk+jCYo2EIUNMxBcV2YzSPbz7a1Kqef0GNQdy64nrz7ReIk4kA
Mdg/0HspHO3bOD6l7rvQjS2GSt3lwM1wVINmzSPpVlIwz+/VxswwiHT1WcvLW1D6dFP2yc8CvFMp
eDFDtm0rTszGdAY1/hqtWRJZptyW9gl56gH81P+nxXdrlC3XCBmzd5MwFdKxpR6aPRnPnW/Ho0Om
6XdXAD8nrl3bVZXY4rr5Mr+rBT2UjmpdG4eD56CGZPJSuBhTsXCL+yY6qd39NupiCCQatcrAJze9
Zbv1Inqk+CYUWyTYmVOoU4oLNzHwEeY054ftcQsk7qx5uR+4cfWWrEBJD1xF1pJARmUUBOq6nb0K
1DGTL9uEPqZ4QD9SAtXfEB0/rNS7ItC8scOCS8bfuWHnXlCTeYeFzn4j1Qs+PKb4OkSNBaKpmG3T
tDlPs5m7rolrLAQXxa0nkgAAlvNyndQBnxDSJ18KpbzQ25PL0/JzIqPUYYw8l2rjD8E/nHpYMV2n
Bj1XDSghsnTcoatJnPn9hLe4AguZZspUFQwrLd6Z0SlfreoAQgId60wwt3nbcWMk5x5P8ZbGfQJh
q6EbhDNbnz4sHQ+MQK+6hWwD6poTgxlXrWHmM29AY5VCXd+nggGphe6fpjJl5jZWy+hyK3/IiZar
N6IZ99i5aj/Zzaa/eu6LwxXb6YButp1Da7xrw3kaa33iCJHBG8AJZ2HDxgrogl7A2/7TmhNh6B4n
YV/uyfDjw5YdsHPwZ4d9dWz1IrSDBHWkBfS/f4rxJ/vZSQFBBnVf4X1XcIseT6aD4hSM67Pid9PO
ujkB6UP182ETYCmfTvjh9CU8EOvyXAUQqqMscr5mZ2Ng9ppFQ+38iPdDTVzNEsmX4Xmda7xbBtp8
abqdUGyS7/dnthbvRHuoIxJYcXUlLGuUl/7wSQVYL8A9yw6mf1/UIKSk9mvNM0JKd7/OlNr4rIWD
kVF8FurhODn5pvrvT/PT7xfbmv9KoXzKA09QzPJjfQJkFQZQXBzphJJLMUwytSbNVZw9yDLA3z4U
7kAi/dMd8XgOCCsuBeBz3QWA3rVlzs0sMFvqV/HwSWeYZcgdZjoNtJ3xSq7ZKNMvDkj3ePIngdl0
3QVCxywC/CzGhyHNmCwysGOOUePAFPoI/Dcic+7FZAlY/8rOGYyLiJSUZigpa6ndY8cA6ZV7uWUJ
jVreE7HIQrWi48knBm/HtrVQBxhQJ5W2H+TSbkuwlOqHFI5YzjlTBoeLwPD/A8KT1w0DSXX6w0C3
8X6JBAoYQqCZBfFTQPbWvrNBHzRXssyY87PmBU77n/JvAYBgj27eHtQlKSmIB2VkstBs+NioTlkz
0tl+513HxqglVTUqgxGu+9FqBHLsJhZ4m32gtnKoYS1OTYEIBW8zykuxLNxoobeuL93ETj/DtBTT
tsCV31q68PMnfA++PBObac93GhUBiCg/akTpvbDdOF2eOwwd9AkRD+pwB+ODj6WBEffNg9mDzafZ
AdQTlYGyikog7yoLFgSiTwUaLoeXkpddxe1akCn90LSXy4VoOx6CC8iOPSx6MZgJX8Fkm6cwTfu3
29w9lLgFc7kRMxoFoic/YGf8c3dUuhtygljkXZrQ3Oevi1thf7ouRjnPJuOyCNnIwm/zKhEzb7og
APCSgRXdzAkVnCU9MSe9IrjEhI1wPflodtWwT58vLUM0xv9Di6RDtvdzlhMliUsYJIn0L8FUeI+P
ewRUvja94OyrBLdxB/lobQ0Crm6itt3zdLGMcnwrwlDWX3IKTDyIE2jknYTdhRSHwn0uqKOHu2Ny
uMw5SmVby2cQLRExppue69EjepzB6hyTqr+5GnXnx8rGTbyUMB+1dYQbz6EQOd9duzTO7RlMy1bi
Rw8e35eeGwNaI9ZersFFzkLc/2bCILQAgLvsF6ywPV0OX1jzA4XwLvQhIw2T6B5yPNNjwEQ4Ryo+
haXTMlL9Qq7tFKOH17cq9q6J1gyMYjU8aWyaeWvjT0kL7l7NePyWuCaxQrj+oXYhHxNypicUKId+
iACpX8Q7RRj4VA8mzYtugSr8h++vAEb8ayk6AkQ5SY4ePsljbpwt/DMzQjWuO3X848/v3R3QZmGq
5QN1Sboc7xuWqkos+m1Ompp5tFiNyt1MdUJ9ARXQz0797TzlRGKa+/UHuyuBHdLjNRYnHVI+UZb1
9Sjm0/MqWC43ZiAXjScMEMnwZPMF8ZymFYmD7rK3OH9/1RIbmP+03CFJ1TZAtdr/hymfSICVgLYw
K3d/SEVAP9aRoD5g234H4P+0JGfX/vzlMrQJMDsWZhfGcKDM/vutHubd8slgUoS9I12nnNpeJM7z
Bs3iagTp41GOE48sUnL3wR+2SQyaf+rpzlZ4sd5WryT28mPnrraQEbZpAqaOvKlpL9RUwsM4+PY8
znU/6eEhGCFfCITi7aRdLubxEUFhb+yF/COMd1ZWAGGFNO2cL0U+T8EFBgUOLMA+QL1PaxQJ8BPx
lPmz69xrql2MP41VYcO6j876qLA9c3qWiOU+rCClYVMC58TYM184V8Yfmd/9lBcNQ+6JDC3soQ8h
1SziUozzcBQL7VxASOg6z+qx0DFxAQxKbfHHGI015M6NNzTOkItRe/qFI8Her3pW8xe1IIOltA5m
OZ8DNGFvXIMv5haxySXsP6XyCp0YZND5XTdmqTAmQDCtuzNLnbhmFlJjvC0Lz/OCSNv/26hMswFA
R5nISOnAgPBBns4dqoRR7LQDOYhntsbJTWiB41KUZ6JTuw6hGdpUSLveqGUvr/P2KW3VxNHQEkWM
roRCKJQThlsmbX+sRs6t/pB0lKuHfc1caJDU9i/B+GSrCV+2DlX3dnux5Clhwot9X+zcZ6BUmcJe
kzwnj5OVHefo3rmxTI+zcATRTxILn/cJtTKcCilutYDfJJgKD1Mp4Ggmj+G+cALZ1bXDOS8vu6dy
IOQ+XbJRggf45N1nJ8cR1LjXqnY9pMCiF7nw2c4lW9Yiaihf4r4BJPOs07vKkA9mwlF9ZIXvHoZ0
HYUPWUxNytUKmqqQc498SsQde9xM82FSWu7qOx2uRqfsG78ayGj/+mKAS1XTpNJnJyCZISE1r6vv
UkRY3UOduEQjxvuyRuJF09H+OzcfE29yiW+KyzHM536L6BtUHJTarsRy7RRGv+TXSHXJTqhXi3K4
sjHt7WyYI/fGvs9XqH2/Jm5a+SP/wMM02agPDf3x2kcIOuG0LnZUeMrmKhfi4KbKMXltOnABi028
q/uAjPhBYqXpkYW/zReiMg82ZeNhSEm7qELTR+varmHWEAmqxYX/iU1XZQN/L2rNkQvU1vGKa4rj
tYoPBgSBBoI8l10C0e2CHBAbY/adnqwP/Wzh980FUe45Zcp2loEtdIvhh1etebu8N1Fc9pNHBQM3
rb/CdxZ8n9H/DJjEKZVOGgnudlEJyWOZ0MkorVjbBiVkgQifFbjxy338T6JDqzN7Em2BBV0h3apV
aygvRQxmcZd2/YBEVSMqTs5OHt9AAKMPshIAaOA24ctmYTI4PYEl/eK7ooV02+cAoRN0Uq3I4THj
D6wd9tRynhcjDy1zWbFmR+kCSXmQhUVd0/OlMH6mQ/R52WnIpFqLJ7x5qDTL9thFwafwTWtcRLHz
KogdvsgErNHmO2RAoEz1IwiISTsQ7VETc1c8So6y7W9Njx70xpi26T5hCcZ804K4MOZYY6Li81mh
czwMafLtck4STagIzMylOj9QhCpqLB55Jdk4hxu6tI4ANSVTxlhp/CfWe15Q8DCCOeiWs0A11fjr
SzabUQxA8gWiDxTJDf8/FdlXQxOZehZkETc0du26yFpzWYhYuA0C2g2G8ejFAqnaPxh4LWAn2GAQ
+fANI3iboXb2mdLaDAj2wVP08h+mb4JI49b91VumVr/JmXV+8xS6pdOvmOY65GRoqhdzc2IgNJFq
ms/t41BICljOkjXJd23O4rHsRJJb/HRXcQpOE6wj01TgTqkkTOTDRr+mmR2ovX4DXZ+DOwRvWeSN
JCxzQkj12C1rIV5uwore+0VbUYwFGvXfclidoLHipkbs5QJXjAq2PAPlcgh0yc8wa03JBptmMntI
ezh+JX/7gAJz1mrZlfyIOqe/lBMy0PJ7ulHJmqLNjBDsKPfkvv1O3SFvbkUIxxjt5/LBQmaWsmhL
UvthEHtBz1SWKiGPW8Qi9pJS5XN6kBkQUKMSlA9jxHl4CSnN7Dk2P3RYh+skWg8zoxJmn/7mxlgz
X5J0hqAwiBjPxTWPWYJRJCDg9ihcRZljhC8VR4imy0oSQXd9w0elH2dAUx+jLaLOuy03ubJ3/sC5
7dnUucLChElHVVYgje8kerUaz6mdngGv0ogC9Xty5RbByjZ5yR/E2Z6YoYRL3mGCsN0zNUvd2p2w
vzoULAuflBbK/+GU+OhVa4QPbkomESE8RcOzrcihydhY0pGbJSPJpYQaiQ3Otyq1WAWs1ypfGPBr
RwiQbaBCvBGanF8gJ0cQYqnWPlsY4BoA/y6BHdXXq/N+NjSVOXAJRDlJUC28z9SuOMVMCy4J/1na
hwwG7DR4xZNM4xKFU694E/z5EEBd8FbZepsYbSpfZ6NC92wyoGg+1YJ+iW6V95FIf6RMMJ39JZsB
+LFvIyy4DiqGkX6cjvpouIWiXWGjvvvT+G1mOq7uNeIRNQFDQ9pQaMertqLuD8Rcd/ilMvhVn/tz
6z0Cvfm3IGibDodjfLsrj3v8Qt0betThHYbq8eRPQqE2uxSLiDVP3947ajPy3OYn/zP6oWqfQUux
xllYVGM6e73qyiLbyGTMLj7Mb2RkxNy7EiEJDy3BWLEGPo4aOrdRGPs/CmamH2X+LoIDCodvT0H9
TQ9sY4jNCIvpaum+VUg6nXuGzGzRD7+Xf0CiOeglCGGIbQ1IowgY8DB5EMVd6n6D8XHardZuLqsP
4NCPB4e2dEYKY3d1uph/TNIJMlwCx3j8UD4y3QRP4cLlkPQN7vWig5mnu8CJljoB8z46O37lUfrT
JWPGUkrqyy04+DqxQVc4wpoJVD7AtpPt8fQg0mrtI/xszePXCHoLb518wmHic3c8tbCSTnsScL95
7jgFEbWDhyGZkCtuDbA5vWeVxTytJlrW5ZxpxcmOJ7O0Ph+LCB7RP4CwO+VJzHZW9/WNC1z+13Gg
9oB2Bur4+9+g5EhBiRH8XuPAibIFCgtdL9gUcTZxEoMuykTrcvZrkx+nJHD7TkjZ0qGMNAfFSp0g
T18zdyWlZLWl5ydE4JSxg6cefHqWVkkk9dViy+j+nGJ8vg59gQJ41/yhfTIWZBZaKeYn4c/2tXeG
X2i+KBttLMuZu+pEVkIIMahpzI0xhw6k2/Q8aNN77K3eEZNWN1NkkGHBjRvkM07NUC+ld1le1Y52
QnhmnBcSBOOJD/5hvoMW66xA3LQ46x0HUpCGvaQUgj6LDHLbB3MDTNz150TNIt1u9AM77cchdcYx
K3voYg3CjOFjtV8iBuRyCjHjn0xfAHX9xxliBMSBoEwhSHHPim1TLiJDarCHJihp3QLpF+I/Y/yV
JdX3GdpPScmyKoT43iubv3RkmXbxIUNGuK7I5q1pGykNXCLe6b4AvS6i+yDXADsU/cdCWKZI/M5E
y2ae6ojRhv8cEol3UFzDQHEKg6FKhgi2l8UmgWd+hN3tO0SHv4G+Rk3sJB+BR+1REUAGHoxMq+39
iMb4LkQkBFtWDrqBvP3aH6bekzz2I9AiiveOAKoEaKxi9W8R6bxaicus2KT01ZcJe2jsgqk0Mq8c
YZWmwi7E6SzFdIbgpiaMRjgU8ICHvbTk+JScvfoAuX4j++KN/EMQzRYKa6mbSken6IJVzFgGKEdz
B1kFnrGmMNkpDrtYpj9ng7Yge0gfRbNRhB6NfxISFhmphYnNqBRoNWTZqhgr0McitRMjXiBVGA+k
JrpzAMLWnhjAyZtQGa/1B66q6odX1qg2U1y5SDbRYbu3KJNCJuNTuWgOoUUDsdNfzawf2Ej9IUjA
9mdLAnTNoUGvgmhOvrOQ+W2KD05taO8wJj6N2LEnMrRZip+ShYcqglepB64oHw0qVhja3LznbtjR
Tq63mKBkGZjWvMcP27O2TgXVIxR+9EBaXj0LvFbU8TFKXgR4M1KS3K2HGc44dO6mH3/haMnMFL32
eJYfhUaciEAoim8PGiEbx55ZVWiHbfpIZPali7fTBtu4dENFQwj6HcQwjG4bPqJks3iY1+dQ/YII
mBuEpz0psJaD9vkRAd6apHoDUNx6YpmDM99vCvd4s8c8xs9L81U0TVtMBTfGwvChE0LJZsC2ZJZS
Lya5ZpxYGEOBnUqsvjqSMo0UiopvtWhHB7O72A6NM491qf+QGd4h7SEa07noGwTshVecl0pJyUTz
XdddAM/vFXbSRTJWFZj8HBD/y4D6KWZjewJeshWpkhZCtgE/2Rwbzc6KnZJUPNOZYl8C4DtyMP/E
iIYHiss8bAUl2PoyOlMWGjCscotYvGiBPO9vkY6aWlDjgLWFrDl/xDGqnCxxOiAcLdU7taN7wD6A
DU7gXMG1AUGYR6dUFgJVm+fZuSXczej4Pz9hNv5Zv2fZflrwGnXm4fmXUZgwsVU6VxdemBQ2CYmU
Q9clWOVGIrmejt1StXvu1gDQIvDsJ3CALticSUD1ObW6WgOKIVdnIWd2UWDnvz7xzkdik3144FmG
2Hrl9CwF9FMtJaBfBZu8Mt1Wz5+qc8/0dXkpwUAqJAxAn+HR648QrgTTm3VkEZV81pZOz09u1XSG
csSSpjFzFPYRu0qMJUlJRvJaQdKN5KDhp76KKZ9kgF2Mo9gQ6yRqksGB08epWKATg/FUAaaQ//mg
cuCbnh0gUwfNvTxoYVUgJaVFHwqA4+WQjE3s47dJYSlOd5k/+duNxs8h4WaTWD7JvM3mTemIn5gZ
UNCaPPX7tB3gyfe4Fv03UyZFPc5RL2yfsXN9POjsAX04PbgKg6Jvy7uPaVNISzK7KAu6Dy8MqFNo
3LK4moLGq7doA4QW/5PoTWNYJoJxZE2IU2Gf9EFXJmsTOm/sTRHMSrhXPOs6drTGnZiP7JuVcbti
9XIbReweMiQfYEy5vgvDSuitiSPN6A3GYewDroWwYVnah8oQXQBMmImSXb984EunW7k7QBZ9HJ5v
tpTzVBNiuRlEmGvYiUUDsrJOqKNnsH6DMtMO61+2h16IOAvD6XeETUVNXvLMXLrHZCTrXIyihPlc
UwjZM9SYf6IYCxGWgOqAc5iiUU17dc+apN/z1Bh0UEg0p0iobyBepg4QJ5DLNXjqL9Kzt0Ho7fW9
0PnJItvvbaaNEvhwIq1tWpxP01bW00Ux0KtVjuiI8XbyRZEC+M6LCSUPdczgj+/qtCGV3dZiQ7tN
/QdQyoINokaFwgCbEChfT8g+8wd8fqd4h7gPQwqoewpQg8aP1Jg1tnWUxlribRd6UCjEU7Kut+t8
LcwR4gWayFTzXSzjyCvUJXfzBHPcUZpqm/ZHjSW4sOoHNBJRL7roCLfXA8GsGljz1xZKPJOsM1xj
vOSRfyUXSigV9u38IiLb0BtteMvfcP9zBtKfJwYa++NIqhR+yMFraDjvU/SqKVIZL1SXECrqHq3C
FE2smKRXokZYzHP5wr2U2OD6LOrNVXCjoCzbLPqar6FUU8UTP42QEe9kjVOrNboo7TS1/gTL0+1d
AKjpTmR3KCC8FtklzrY+s81Lg8ofw92+hRtUsiDRfw/hRpIVdx6VACcnuXpEuXD0escUv/Aaf0kD
BMHDOcAVYlGMnKM3yCUp1ciUvtabIroX3l99v3wVwbd0R5jCr6B9dB9sJ6RxMeA7mR2FPQEBPhvP
d5jl1CuvbFa4vH1m5IYfmLJ62xlKYkjAoT/Kq6sNZ78O2Gl3ZOXtFbk8uxcx1XgDsTuwa3Af5eSD
tGBcfbV15CNqQpe4XEAeRbtwyIj6rA3SKPXs71b50wJwPXUi3sDo4l+yVk3jlFU2Gf3teEVwjZJD
cSrjeMksmFa3E4nn1Ke8yTrIBqfTUd5TJoiKujpd3KT9S69u1T+fFUwDMLkiIvXyk1HqXN0hyRDa
7VYkjEFz3wewAieWBqzRiDlvaDWxHsXmesSvGCC9KpRsVKzoZk/uC2YMxQcVSgzr5WNXVE4paxHN
UfWO//Jg9HRf7AV0vDs5obYC8jyvh8s/V9SbMgt+2UUXHyLhc0emTxs333kpeLrkRptWVkcCWqjj
zzz1G2Uq6CDqK+WGSRdiSbgTkGCJlpjqAoijY+pCSb6pqUHPgRo6IvRsX+O1XWy4zINlGZeZPWSp
ZmLtAj3WCP0rwW9n//pNBCuF6DZbJppK/BNriOFBup6LPuYasCLyGMUuq4zSr63wwQ7JWOkTpwWG
Zf+hendB90H96wtabLDvhBe0ilqjh2kbM8eQMWU/8HUHjt+26yp9aHyrjB9b7MZ4KbEpcyYiPZYR
89Fl5HvU4E7qzKjU+etwAv3rM+l9cWDohCI35gyxgBnJlaTtoXPYOhoajGzXdrQY5BOhEccRZGmG
DVBxElPbYhXzBKtz3Epc0vdLWztT5D/zl/1HmA4A7LHNWHXQZsbwK+XbwakXNZBwjfpalp1cot4m
T4Z9Cx198E1hvvwSNbR/n42RBjBZbt0FcPWaHoIDml8g6WHAr+gOYbhdKThn3szH3Lyw3Gq+t4ea
cSugyU/DuMB5Bn7hvv7FNwzh5QqtAjbc2Z5PLSPt8uvkMUrh2TTb1k1cyLCquCwnCMFTd1lTDUd1
r+2U0gP+v2nuVeHYShs4H6pwckXiXTT52Zu10co7Nwrjv9DuEzHHprOmt0hY/XIQ2KQPPHeiXH9B
prxh3lQvGLHv2t7W2q6jgzDd2j3sKGGulylZw1abAhX40lnLhYAbyPHspCt4GzxK202/tgBe3ith
7uEoZBpc4gnUJLMjqqsMjh1ejFVx9zduhf/wtPRJvV1oD5YMgCONrofjVI2mKXRlaOZpslPXfP1m
JDDZUKDCwps71GlJpPDC3n6cF9vQoB3u5w0rYG8XgKWHuslpFqYb4+ok4u4vXcI3dJ0UASt6gNo4
woGcl22NDKkwk82V+K+lqAz5+N+QR0kdvFI4cGYBeu4c6/se7Dw+vQd/LdrjQA9CjbOw7fOvUuPU
bFo9AL8WxcEnXNGlGTwkLh4mpx1cVuHSZRR5eSrDWaThmN/LmFERScB5pcw1s2JSo9LeD9G74te5
v2NxlJQzVDPmOMBMnT42I006Pl93+TpsI7Y89GWmtabp3O7FAaQgEab3XDs7/BsimDArIhnNjSQG
xvOouTYOSsL8+3B0h0F7ygDb6UvZsOHgDhlr5ESrqQCs1TLRK0GuFpKH4eLWJqon8oLxsh/bUMWp
8397Sas1GO+lxyPr19Fzl6s2SHUyx0H8WjeZZa/+WiGogsH/pPpjA/+aetcoY6+EQjv0aSkY85NR
OJ70Ma7fi/6iNoIN3HEAHGYIecP/XIecaqiLKMg0FwOIR6i5XjZ5Y4KPFfKHC8V29gpiFsCoOlwa
DPaeZE8CGkMKD4zZzlKaVziNZEHOJsIIQzkGtZ9rv4axTL31GfTH/t4ocXbqiCDOqjQwAv8Zlxr0
l5FZ53pouYQtxw+UAOadfK4jqY9rj0ZkNRuJzavOk3IzPeHcaupNqzeINrgNyjCGBlvXWK2zveHz
HW8Lv851EPFelunbqK7bS+O7AIZha0VfO00icikGFTChfmE7bJlE4kpJbrQxaFEIZNYOCMSL8TSQ
0O5ak9+Rap7yPxPoHvXwWqExq7ztn8umQgUyAIp7OjTKyj13iVfA2C51Hb/w1emVzbHy08NDmD9O
cot48uSItQx3GAPHQ4D2dcb5WDljTuma2oAEshHDxXfc8t+IvGBRL3n7+yG9Lt9XOoU3sGbgWVWa
Almov0wCcaaq9A1HAQETBplFYAMokOfmHZL9JiwkHwwU8obe/Ns9ySt6tssD5jZmoc/p2tjPAxH7
JL5akA9yTypI8pbdiow74KgsB9qZlK2fYPhNKrawyNZfDRY2w2EJaB5F7Q2tCk05T73TYU1Kputk
+CdEmstzTYpTVBmT4ne4nZLyW/AVJYNu78cl/NCJNEKJi8MqvlN07BcvFBSYdL5eJyF10BnMNCYi
DWIY8Zp1fBuN1yoa03rwQCtmlY1ZqFCCB+dyEoYH9pIcZotDFr9dUdHrFN8wsBpZZ6/iTB+PIq+d
agynOlNrgmkTj3mlchT4rinq6BjIWosBj71Laoaq5YK4MM1djDFUGzCtFPZVECG7td4R8B4Evyjc
NZoufy/Pf9OT5XIUjcQNz4REm/ScU0txOPzuizvadnBorTFOZO6mJrAE8tqoU76JOVzVr9FEYhUe
b99jv0RQ/qmOIUJbt5Tv0BQQEKRVDJkZNkY81irxI8j/jnUnLpj4GAlLOMPVWYXuv2ZcUTM0ug1O
OqMzsqYPydypUOG/hPl4ZEJQZSuntywWf94q9N7B8DW1feOqmgSA13aS1SHb9z7kWr5L0e2G2DKU
O8/RNGP1VDya6U9Ne4jfVZMIx3qfI7XfAkJrvwf722gwLRFPnqb62QvrRv1HJZAT/vD0AALhPR0x
2ehsNuF7aw9cjeIVNaYji7Aw5pkT8Y5C//yVpDwSZwNVbvlpix1/9ZFNIsUkNaeuSNT+8OSJkMSa
o95AMbVW+ceJj7TI525iR5sFvIUP9OJElsfyCOW7XAE/apnmbKkcY2QGrqSldyd+eqvmE0cy36Fg
5vaIXIcc6piFtBbhmaqG0ZCxAtQTDkvxtNXyvkGVwahsoxisrwV1fzrSjX7pCmmw/2ctD7hPrdqz
0qI67yiGrTHzd1+9cbUDSQ7Zsr0gmMb19LBdpuV/6PGPmqU5VIifPXe8n9PkzjTTB2N/iZfOOWkZ
mIPrjVpKV4xAW/8mQTR80GxDU6EDiV4LYBKXeA/eym0oERCbaOlRauqzg+pRIvBialKHIgfzTd8W
VO+W1yi/O6/acxsMYo8qFzKYFgI89q3EEOtpeuvGlHxd9ZY8qyrFvuXGfS2Z7pX/t+XaBI2BquwE
FGcQoE8wYUDQpBJsfWT4fMZQmDzZVMp7BexElv4sjHyBvhgB2JSKEeLaDhCwndoSUnio1F9L3xq5
Ki3K1nBBaw2cdOn4OLlCwzCXyPGm24Oi7RulZSoVO1tVsG7gYIaRW14WMDmGUeWojwfpmSC7B6Rv
+tzyRZOwMmhSLp3UuIFKmCAQww+KkUDwXFIF4Fd1EIMc84bailyfbbaK4P6AU9AU9m2AIAlKQEgB
8WphPYoNIwjqJVPjc/eshZlxcTPr9ZdVu/jp94BtFbac9Kw9DV/XsRSdfD8hNOzDYr05CJPkXUsY
Fk5PobFHRi0aKS4pCShboSBBlNBLY8ocLbCFUd18+1XG4bVN4QyQY98FO9FUf87VMX+2OqXegdey
YqhDBcP1hCgKOgBW60xC3cNQSxZ1zPRk5gzT+amOx8eRhcZ6OhT2WSbKNAs+EIzqUla+wofqmaE2
DzPeXD1ic9PmusfTQzQ+uoYBW6QACDIh+WNuYXRLJk5BrBI8JcpOjbbix48s+Oijs1FJYcRJUdjz
UKcmbmjkZvY0CEvASTjIkivY+V0KgFQzAchpAnNoJjlSTnwLVmXYADANb1KO7wVSyrQzRT+nO+zX
PfjgeOMQIArQNc1HY2Ae/c5J4foYzBfG5BU/wKDBkrGXuUfAodoFhXx24yoeNkZdXdCp9mM2Hw7x
5lJKVwxxFh2igThbj4cURKy+OGPN6X7AYxZBtFvA07Qpbk21TZpWq4qdYBbwX/CpI9DDjwkFMp4G
3SGeHiLy5UUix21oZvk+tTXslHSwCgt5+DWy2wxOsr+KoC/L3rp0jNEXC/B8v6YM3wbuy2EKMYH3
q48awVZWkDeW4GjzBvc6cjZwRIuz7n/5jCza3gn+/EBJXWE0pUM/nLbrGe6COMfUZj94MlDtvBR4
hILKF2NdzJlMhQt7mmb1xsXfBWTar8adXoGS9ksEfLpBplK4kgZsVJcOJ/6Tg70fLEIYNKgzltFp
CSJYYZtJapW139qL2K5Jx7tGGY9kUDNaYxBcQM4yonhpz5PtmnDAHLIjVPBjdAM8k5jePMgSWAoC
JmjxbQeucfQsS7UCeR9mjwUeiFPpsaYYuFAjah2X0ntdERixW8NP3ZyK2rPEVX+Gfo5sVnuLP3C/
Iui36tXPHrO9ufrTyt6HsJFIFVxv4I2ATLosCAjf9bcGMmkaQO4sGOrD4j2g1Ugfe7lq8PbmRaJk
4rVx1442bBCZVat2wyuGcPOGXX+V7D16g/zlImgEWUTJjbnnjYzoFonMQDp/F54z0ea6i6pjwVKa
+38R7LvAXRdlYoquoZu3miQg2CyXVPgGdfcUjtbrCWEtCgKdGsZxeHDbrfbMz8zMdipwDSY0YtDX
cAUQo0B8zE4BYj1GmpAOcXc5VJ5SDYEuHNfB7shjHM5K5EnNmjE4YYUTsawszQlZAQ1R0lO/yuNW
2RDq/U4V0O5gIJlqCPHUHjQ8XZkq1upLkwJ8rEXAlEXbrWnN3eeuxwSa8AE4meBppC1HixSvNq0a
C2EB0Movt5GAaRTW8IGgyAgw8SeUE5N1T6C50IHOxnS0Rf2a+AyVeew4XfZDqYvi3LLhJ2xg0wMZ
632vicK29p+Adfg8WVzC95KPB/7FMN4K0sk0JqWYnjxeb0VEjju8LuEpUA0f2xyNOV2kJQSrWZvn
LTbQ9mUDT0+IvhDvd8p2grbOdkesFJo6VK3P9X7m+tTtYjm02+dPqlE4LS6tATRwO2C3XVc4ywYT
5LRobqp0GzHN6qwSsYiRsEAQsElF71pvqb/66L+IhLFHvFHE36T599o74U0K2jmwA6cb4UIKIT/I
em5xuvrODWQrZZorKqc1WbVo2wP0tV9RnEiGhOgqAo+zG4p4zReCgL77yqMcFYZyEtLnaG0r5gww
sjZ1rLXgXHgx8NgJW1Kq9jAgkP0I6+Jl1Xf+e6FoSwpUqfLFaAeX8bT+kPWK/IPege2ry+D0UiKF
Wx6XwT1YnFPnR1+FI7A7E3wnwxI9JzSL5lOZOHVyT1whsghjPK48JbL5kL8y8RREcX+fNiq4e5bV
VR0qkwSsaHNEV4fCpT/oncFGQ9DVWBUASnHCEnKzVcvFYnY7jhilysYxG9Thp9+GlzQ3YAyEJK4X
FiEMOSG21yQgohPJaMf25Ca8UiQswnZhzlrv5TkFr5w90D2cAHXZeoEHOnf/atHTBNqPCIAXQpnJ
ZYK06lvfq4XtNipUlfGkY0HGudU/0zGMr59OCKD9jYY2WZh4mez02slkPiaVgJC4YFkoCtRz1K1v
vM61iin6rz8XP4BKOIMzLvQJq1sGLlGhSYfKwE4RDHAtwGFmKo4NCh8GCIE/vIy6+ixGfFNv6/53
USR5Y3oXed7HcoiNOJlghsHA98PDe2idLom9Zs9xxtn30ZKsXp4Se0Mt0sPU4Zg+qbjOGKaerD5B
Y5v4eXsjKweijs4HJlJ8o5M4wvcVaJ17AXru2c2TvvhYCcCvB20BYT+TtvkqYUL+6VW3H6uvrQSf
vp2KMDJlONpdRg9KHtJPn3+zFxvfBMKCJrqeA9qRzc6GDrqjUwg0MNk0CwocTAEYADFvo6u7/EyU
6PslGK/TllCLCjiZSz4D10q2jeMyYJ+6eqGl9t5KV4h9l44V/L2n3xzYf1VZCDR1UOuHsnVN72xh
Q1ekDNnWSHfjJM9wNAYDEyDGaqz1/CAZgxwA0c2t08+ZsIDJ/DPqGHXrDraOolluoSXWQM8mO69C
WCZl4NEZ62KodnbsYHn2hkYh8zEvGPJ2MkB+IDoQf16vYqdEqb+GFBQCRSeZ6a6AXEhmoCjKzJie
7/mFgCHZg8vLsUZkIm1AxQM8UnlEKIVFRijuld5bMcYnUn+2iAC4muX3WA5tx7vnDuv4iAzCoxv6
aUIc6rONbMDMJOmhFzcKWPD6HZNssM0SsqNFfVkAecYDQ4YQ7VoFy/SOPAvbiqJ6KHclDEMDtTMv
5Yev7YJIKCYdh1xsB5wVV9Gu3s0PrQdOSa0rcYNFPA2aAWQbzCPwMYd0cCDQQoVzzFxle4ckXanD
bDw8kXJC8y6UzGQCk7wNF6ESc1dLsISOppCigpGlFehO5TsM5rLeNxhaa2EGeKnfWUNX33IFab4+
Fl2z/FYvUNwmzKiCHnxnQbADoUJCSdolVd9dnZTuuMwX+H8Xo20iZ5m5BJh+aIlKZk4u3n6zjOc4
TpfL3vj0WVd/JiaTGCCbHEwUnvsIM4CCd88Q0s208rJS5jIpThkM4ixE0HomnCnlLJfsbRw8LoSH
CUCigVB6hieQ6Pj0TJxgquR5XronFhuk515CrCQjqKtIbMj8UPo7an/b51Pk8rIfR11ZosteeQI2
D89myZ5MDnYfC10l38VEe8RdA8WSo/xDftlzp1Lxr1trchFS+8+bMaBNybhBzZeiy9etRHNc5wfM
ySSG6iEP1k7sh4u1CSkU/Qfr+1SngG7khuplHzi2qqrktQtzm/ScQHo3PzlsT0UJQHFZq+LrY23F
OR8d1FdiMF+rDYZy2GkhZQkPCgXXwPrAQ4wqLLkTPQMbiN34hL700Crltf/lEqOg/ATd22WJXyp2
UPoepemi1krRRIAwmXSTC/7rOvCwVqzDtEhYcHMWESin+Kwslxn11DEErGiYAuoJyMM+3YhHbqUw
1+wkrB73LKa7NzUeqVJaWuTyjyuwHCPu2CoBhiwlFg030mCyPbJ2SYYP1e9GmyhB766LyNPxYLWC
1XHDVRTl2DwvNyivF40mxz25lZp7lgN8BU2dVGCnwwVQf0WqjVDwNmXqPuQTUjwCyymh/l9UeFqf
5umoJWiQoipYqtzC2/TA9G0rbpMFNjLsC+4+gRldo7Iu0NCYhcIK1gpRKtW+YApm2S4BeK8OpLlY
DRwYHeOLtm3WzOrLPwJ84U5dstkOnCId6WJv5AdnBh28UHx9PlkYM2k3Nf8bsNa7bIYTpC4tkSun
Lhs+jaFRD5Cd9AohtG4Iqeg0/3MDBcNBaFyQNkXsDc/XuNmVNWYUY927TGYw8JRsjc0jnbDfeS3K
uMaGwHH5K4PNLXgUoFvWdFNS8/y3jb4cga4+oQ95KTMytddiuVRjz79e99jB5k1b++6oDDcMdnMF
nZIdMCjd0OMR9M4Noovn9FrNncxUc/UHSbyLYbjb/NRjezpxVWK6g72xFKzA4SkBNYjk4gWjPQRo
g1fHUWgsYpqC/k8DwmYN0ap0v5QE7WONPQGfOSLkFlm9C2aaC0IqA6tBCg4TBOtHGt/BeRG0YxJf
C/pUmYWHZ07OCr3P0kM4wu4dpQEVMAQIJaqpHo3iiz2o8lbOXIkIgBdgIbSFF2OYo/grVuLvRQnX
RlRpgS/wOYaAIjphYtf88QMy6Ee7BlPgcGOxFgtKPkAtCK3XdSeP44siBXnRiiwQVAlM4NfMUXUS
f+SiwhdIjY2X6w33G7zaVc9abbXSAQ2ciR6CNOIUpZIjFnjsWzKkNxeN8vUxNiGrZGA24/c9s6CD
MeAq0HN6f2cRWazS9dX8/w9OGUza/hUWf1kZNrmfJ/GdEBuDhMKCyQJ1g5n2wsLXApNDaw/mZHug
eSF2EKdfk0CU2Thjwk5Zkzms+QcxGl6yKeUMqOX08AeWV1NNhublafXWpZMUmoCpD7Z+7dYO8A/E
5DS55uCIEP4/k2/G3T5JYx4nz97IPPdOAKWWNBq1NlzITS9rmfHk/CT3hrPIxjYRDlZ9Ri1lSlo+
GMDm5VZcMGDS272t7TaEiLY/N8nt4iHB1P9t800jXi+u6l+PhQ0NQkNRG66Ua57Jf22RrQxbH2NI
t5aPWAEKNGTCsHgoHp+Lr9U9JVWrdJsR4mPPBzpIiut3CwuoLW82hpjp67Qv4xSf17Kz/e0XUciD
1tGAlDFTz/Gr3rb6+VBKSkRGE0a922iTXJSLnbWgGN6g0Otj6SHAQGPcBFParslpTgMp8oPbJFtC
6yknxJeuuU94wN50KFhspuBLcKvZetNo2RwGhhywIS7u1rfsaAbVZkezwCE5oAVSaUbYDAiaRR3A
3NIxDsrp4q7Hz1v5uRN6aDyM1mc0yXKdZnjJJ1wCBXZ4QMs/c2tX+QifbHy6rtYL8Ntn4rznX9e3
WIAYmonJNvQdqHtifngyiMKD84L41hLniHikU4WgSxTyh4hMs7qtPhx3CKv9S1vXtFSUw6UmXiZy
0hZ0Q0gpRRWnz3UTRzOxllKmB65JIGsIl/bbuVDSxf3dAWptp3quUC44nlwg4figaxDlcso9Qckc
JI9wKwFFBnrf6XM/KINFf5GbkbJcbAT2DezviJmvgQqLP504Gqxx3F19lQVYkaITmmrpyplY8vGs
Bil/p4B2EHC8DocMWD5pOQdsMPUxh6L6dWs7FAnekWSsmWaWQEj42vQSnIJf6sny6WyeDgnMoIay
PH04qqfOWN+Y4a302rgrQ7iwtRq8ffa3w1QhIK0Od8JLyrJxrM0+dbW1Q/dUBWe6+w/xnCQ0GhOn
YSugMSs8bC3m0h1c6jVn+o6niYZyN+1Pvr+1Vq7Bg1rNzPxsfp+enlz3Vs2uFIpw8pPhK2u71SoU
2bzGVe6Pj+42/N98/55D7Kw1OAydgZQikpN14yJKnH8LH7Pwj93ToR6BRhIgagkw/T03qFXs49G9
iW5EPfZBhosarfblHsM2YOdDqjgWx61VGQt3HyV/3i8OW6deoImSPDivUwafQX1LoEMQW5KzLI/Q
8LRbhyr6mkRYRgAJ3/x1mJg7nOy/YRf7Vo2Ea+rrHi3uc5yVjFPKsR6NExJcCzQMH+3ytZZWCkV8
ftcQQjpvASBW1B/m0L+6g1+JmI2704ru9gC8kUScq7cn0T3fMQkmEoNCY0HpF7B+Wt5g+s0xrQQj
I3bfGdqJAYNo5nARRoS7rSn/IhmtB5UK5hYJ4RYmYt4qSfz79Ifk/az8Mvlu2xJM3trYnOI7eXKs
/UPIat1AA0+Hq6lqIiEcGFsdcv+b9xt7P3F6/Lqq5OIxhuiQ2OQtmICld76IfzoaKGV9Pm/vJKqv
86VuIBWSpxlmWOT9vabv32KNl4nV9mgS0iTrhGlLfpmSzP9KpaR/8qhXaommDEUKaerrJkfYpWts
8iP1vNJbSzYxzRD+lkgy+N51jEC8w2eLGvWXWLqERd7UVMaE33f5hZH6X+V2ft1vzjAm41aQ/vuY
5CU6Ki0Bm5sY7X/I5P7A4KjiykGJN1zeyQ9iGDcuDM88lHyJR4NG6D2JAk3Q5obawozjW2RcRUL5
Ej51fDvXmk+DSF267ciwblo+SdNb1unEkH0ukeaI22kFkR2b7P1E552JmLihbcKHMmTNODvNL345
pUHImMRClSqfC9ICLnEuMSC5Dvk39Xdk2ALiDjl+ufJhtckTyNOnR9YBh2V6jjpoRgFsdCdVUA5M
Vb/H8blet41jaVj6/F7zMazZDx8igSG1NTBKXf/PWRtqQDVkxR+upqksx8U+UtZJ6zYSb7V/nnaI
5YsHe16rz7LyNl8uggU3/cxm4OVhELb8ewY8nIYMdUqbLB/pZemV94El6dBqXOxs+Ewk4SEv/w0r
gFcy/S6k2bRDK4CemzHxS+Rv2XcsQoc3j8r/rcRfVZ66tecx9sE/IlbBYvMJVnxkSTf0aoKsKOgO
T/FLo57vniRmutbDeKfZpdHZBMP76vYi2YbN/wim6rlXtmmCGVftCGYba5V/wbLnClajHlA+IMl+
I0hQyBdE5UtsjlVIj2xSHewT9I+lCzxysMD4Y5+02YyRUFFSxfwo++oih6uluOvngpILfU6uGPTL
B+5YFaTE+ETo4STqi4uxZU5Dg0neVbnpjQeblOlGAYvZAUVt3WOy4jLDMNO5u4lWH5IOdxbL3scW
bFIlcIZgNTNykIm/Otv6xlEtWsabVztcoYPjBG3AFQipgBWemmXJ2MNwTEX9gbnVvFkd6MPZwFgA
U8vWAYgrU/2Eg62ZrOIQRoT+OJyfXMD86ggHDEv7Vm7tmPiqAzH8G7qt3irSgCP5yfw2krhr8TeG
rIVqS1XS+tUS+wz/QEzWx1l+oKbEcwu6sZCepHV8kEm8VckN/s0KG8dDqv9DVB2R6TLLf5A7tW17
V6rbcqOqFj0JyQJJfy6+IIrwrF/OLKUwTzwY6IkDkGpidcKc8thyNjHWkiZpo2VzpAUPqZ/4lq0w
ueo/dVWbzuPrdYFhBn891bt7iafu4FLvN/1MbiP5a3IeKjy+IyXRUW5KVmuLabYQ7bcs+Dxxc5ob
AUxxvp5a6HSf8uzkz07/830cj6GSrldrKJXsHA49j/E1HSWCFJP5mb8FRWDKOoiyJJjT5EUp6FHX
b8EuwLm5KqVsFIJLs5LInkqFfHUA4xxYaw7A0LmRSj0Jm1Jf8+f7uVOK6rnLhR7ILGl6Fue0QRV5
E5veFBcIxgtnEgZa1fL5tmiGFPaSmxm0Hzl/Gkidp7PdcBRJ/X4ivVeiHGXcFXuUy3cnUdZO9EdR
5KQlikNXc2YMDj0l+cUBcrR2kGs5zRjqJIUlimpi/riWBxvJnIYi0ZPovK4W3sAQvKEDYjbm9oW1
R4v5GIJ7b7jJ2XbddTVmilWtFqbURRQLjRy1oEeDyf+gT7kkZYzDu6A+Ml4aqIS6azKWdrAuvpAu
xg/ufHxUmW9crOo6v5gAvyWNQcS2GhuNCOWL8+3mcC0ZG7J6cXN2d1/KV1yYJfh1KExB3ICmy/vN
2gxYM5qEK7BMTOvkmG9qNdj7Xi+IWi5qxt7NidBq7AoZzoyiYyti5VXm7ITb3UstXSRG0GmSntQ0
4rtJ2FcZaHYEZHURQe1ViS7rVPXfrVZjQlMb//olnreLDAeGquFWH9aToMnK0ZzGgn5V81zftlgK
d/2pzJaLvxHEMO48102KteQXExu3o53ma8iK0K55Afzk/Qoopvua3hWaE9gaYvhpjoFYLZlnsqsT
6gF37kg6N+uykTgcThcOkDsqh6tBznLIemunAwjFj+rN5BLu0/VliIGX7lrXBR+iQoojGmAVnMnL
V/MHl2FxXdwP4/KZdYP02JuGprLZ8FciCh7H34lDUsyf9UMpkJ+Wbn32vNHDsTORxIBioLIuci2g
Ul7QGI4D7bfgxyAv2NIHwOO6QuPGeV7vRa/Vj7tNG+tapsgrrR5EGmKlJOx+cqhblOJ62h8kA/nY
CFBrSgLGVe3iWGFgaz1Q9EhMeI/XwCVDEe4azSRF70xUS6wBEGYstZROdld3J78nvwxOK7NJidwr
KzB+oB1vdXfQoi9B0n0UldG19usl5CvTBvws5dpZjjCGirUISOY/DlablxnOAfL2PP9Sswo2UkJG
ExCZ4HE9IfWlCV+3CiV52VeKAFJwCCqU15ezBioX6IG8cKGQ0C2E3RADritI6n+8bjfrjbP4BtNx
cCr9e+nA7lJAY+9KPrfXoqU49boiFDk997DKlhLvLLGzBK9+GQFb3b1DSm+QVWosvK6Lun+iK1+w
delDXAKeIVL7j4RI6KwQasBVA+NKZR9p0fZdQvL7zjb993L+vRPZ4sNlgNYYNINQgHrFYpTIn7O/
TtjTgF2q6pFK+3e+plu9bzM/CbX5Tp44gNfphEps/5KOrq5qjaCCwIqnYbiZ271NESLGkffYcd1O
IMAVcrSMVvNsRTwNiYbjl1Dl0RwL8RPTTH2UCqGnaFH40/ud1Ii5bvpduhT/LGe6fSQMW5OBzt5R
EDm9H7KbnepEKKA+l1GoqWmRsWS7HTAlV9s+i7NwpAl1PGQTQUqBqR4zYJv3gbzGqKXjvMHLvA5O
G84SLtYE2svILS3Az5LBz10B8CLtX+BIic4kln6mwer1cx0bEUIQXn862tuCyPsF6uPSdGKirz4W
NdyhDQ64JGisMUc28/cedxPCvhIwFltZ3buEDIwOKW4ge17v7QoqKcMoaufZcDlMu/Hk2GIncV4q
e9nLZ730rqJayqDMwnPoe2NbjBhuaZnjSKL4rwOLA3k5xSYcz59Kw5NPAjGZdWedD2tdut4ser0W
O9IGfF6M3WSdnTNqlNS5xavTo1OxhkP7qao7qY7cEyQn/Hbo7ztwO06A9ZPHgF0DKi2JX7wPfwH2
GO4IyGw9lSD1DSriHY9Swp6Wf5gj2e9n9dNkIdhCl9wliy4wmcRMWAUN3CV+euVKaN6zyCgO1MoP
FqxPkv6D1CPLQJAX3ecDV/1C3Izqh83DdxZ/UZSVpjocbaAwOstdOQir0aU+twbqEdjF/Skv5PHT
4WSnMqEGslZ3pTS+Y+BfzSzevlGIgL1B2wY+Z5IxWP95JvX1e/GmiDABfGRo3JbCnJcQ2FNm5dca
8Hbay/dtmkkvp+LOALBDAwx+y7brR3lNJxCAaQET/SYoyUaxxmbYIUumq9hA2S8dOWFYBf82Fcu4
iYQ8XTBluEfKphDe9FfdjPPMWrCzBo0iDFQsPJ0AQzWvi4/KOpTqqjB529sEejdfZm3kPmKtKx9I
/q7+igLa4YaZv109rK76gTWgl3s6xqq4e7Pjl4jdGp5p5ET9SASVDSfP2LeFklv+POhpkBUYCeTy
VaxmV1vd98DHxNsdmVMpzc1hbPwm5jwkw7VdR4vvHei2G/IEqBA+SFmlnEdBwfu5svE5K5Fie/SI
/0Ugun5dXMq/Gh8Y3gmeHn07T/wtxfmyn4eXrlzFn0Z1T55yz5GIHIHay4I6LZmPuOwhDT89d81t
+lqLezuNY7B1Id+HpKZ0D3KuDg/Q+34QTmumQp9imFRa5yPeXNAA3dgQklbVm8TD3L+UTjlvAVAz
Rfj34lbFSonZtfzs+Fk0b8LTCaznw5jroRhhK9RcFogiqTrJvs3Pn3rgpxOc+qdLboH4ASKhpPqv
KcQ6NLSXCKBU+zVvJEUGOS0kt+pceFKAnTtbYtMxM11qWmQMm92UNeHUgnZUapCjPGO97xhCE3pK
rc/MmMVA4rWjDQUR5esDvA9hsNNYpWmijZLa1ASTGQs8lGn7DtKnAhU30t4SF9+mtc4h5lwfVbDC
lJuwvKPZ/2Lx8Cd4j9TpA157XPHD/Vm5dRqIWFFTdMUv/Rt3hZmvtktmxsZn47Zqqi3ysftsnonG
xziw3smSeKel8vddOsiWAO6g9MDqcrguBFpRl/dzQ/0qgVWW4PqpqgIvOclWR1GjYVc4z3zg0ge8
cTf6QpPuuNBH3S2uphzbSxiS4OBmLJ5Gox+y49AirAWweVA9ru4wp7xcDpFCjAN+Id+N7AwIj3QX
MU81Wp3GqooLyL2EKYM7eGadJC1v8E/98z9YwCW4sNos32Qd1PlZKKTjbnJ+nAGT12ZSgBkDkujo
itOscVfpgGnJbhOfWTzEWa8945lojhxATYPlsWNa3D4bUAzRmkS4bgqTssqna6bG0NVo2yytshe+
XUnryXAw8hxg7bvVC9jFj8GYpodPevshO795nYIipTqqejtoCDm9Dl+d1AkPs2T6+g6O8FUan8d5
Q3XaqstAysmvcwhpHdNFzk34zocwIwbwjIH3wpf5rdLVoDCyQzU3U/ABytf5pisdpoboZ37Sd6Yw
XGroN1JpryirBiIPvHIiq92+cW3fFeXmOYYP7wPeS10WU1yD+FLq6z77NbC2kPCEzXUiNvWn4y4f
up2ifbd7a3kG5h+0CPLwjl6LMV8aLcP9yuZDxU+j+UZxeoFvIBGFL8As7JynihlDzbX+haQPHeSW
NWwypLnxglozdKLNbCc6VjObPw8Zk1yuulKvsQ075TrkI7nxDd7+luTqyO1r78o7ma+lKPb0orLT
9JA0f4LjhEnC/vpR+RrqFayCEc+EM2XvLbz0Dlfj3TKKlwUuHExTUxwrb0UzxFdKuDuZfJqmgn2E
uXArqOz+cQ4cctaPQ2CnXEoCl00WwE8eoB2piHoLnPwYMDI2hps0z4kkKvkTXR/8F8N1PVB0+oZr
0mGxgfP3PwcKU3bBLGU16TKxYbLg4DtdR3vrOoYrfctWuRRN3p9T69gIur9Ni2Baj7jrqxSRKOES
Jg3oKpwaADlT0jQfpoqId0+o1IpKHqkUakV2MNbdP8JRcShaRSCIen97Lk9if8Y1UbpS9d9bQU7n
VP0oLW5eULLfPfX/p8gJXvOtq1V+/pp+ymKmfH713+qdN4RIO9Oh9WdwNGrJn94RdLcbRKHaO3Wi
SEePSD78UL8hRnqnV1F6t0252ui7KKevncuxQCmbJqw+GYvtNLRJBpF65mIDJw4YjQRGCmAJOlZ/
KIKEkKdukf24QSqZIn0EyxZg8w/9QEWgNY+NWjKYCIlBwl5TTJp21IilLus+LUS+XB53ma950qfN
jbee2gQ/K6/oD8Ja+o1SoNr6dE6u70yKMIKA4LaWcsgyCFjPv0Uh1XB6Y41iyW3+kSDdaXFudn+Y
EuBHWNTOU9r500AS2UKd+z/L2I86FcTMQlV0VX1jMSMV8yme0sbjJKMElQ/AT5n3weGX5nRLLuG/
bXzdkNIYw99lfQl/5tPrITo1mnhYqrlSuLeM7F3b4SxikkmCkRSclXBwNQxyR5ifhsaLRHtz5wUu
7lc9qTwuoAangWYVhbVn7PK6HQUxl7VVbOMkTVFHEjOUdZKOJPX8RhIY3HMu5ZB7NZ5iGobvqKSd
GThyuFDYj7Uyoszdi59DhjDrikO6O45M1NY2zSqCxZbIuzcst0GlRHqEfuQxomll76dw6L7dQepW
A39KOp1komyAOirao1HKMNScXj1T1RkJwCPJDhXRFaQYuDwhulyKD3K0XIfwuuiDig5Ro6KGzwKK
piSi9qiONkFP3onP7m8e5l9vRgA/dsagLAfx2Y3SQhh9ysOP1KiVGgZ66U4SX4cwNK1QiVoqfUpi
5AjTrjxCA77/W1WYKHuMvQnu8fRXiOHpjWYAzELKEXG6IZapcx7zmChA0hvqa9cw5G1sN3Mv9dw9
Iy/KzyQ11i475ZLvcRZWx4YXgna/KOvkA35YoTjWaSj9BB7IvGe2kIFeq5GDbg1r46kxcrLC+SP0
EtgHYgEVAX6C90AeZ159AyPKkyDcZ3vbRtoGvddcPGdvO+QecFVWBvmVHVcnB1i9aP4rzJ56XBvs
MbbamgGyF2djL9IIjOo/vvuE9Njewr2ImOeMD6lFkn82ROA02PU6xw2LN1SrJklsK9zMtBRoqQkp
PZkUgmooBRO05xnkbc9bDLdwmdm1oeEAMO5yaqrciOXqaLiXnJEoHu3caM+n+62G/qtZjQKNJJoW
cD7T8pcu4/ndJPe1rrbW1KVmmWooACqtF0norB9ufcHoYajaD44nqe1pSrQ8rmLfP6niB6qmuCnG
wttl1eE4INwD4sjDAhUB3WxPku7GjvAg0d/HvFz5WD8LpodhHOi77G3HbGMSoPMsBU5hpueVp1qR
LUipCh6cqoljMwRkbmUKCmVzQDRg+k1y41Gd21wHp5AbfJ5xSl9piaJT4edFMVDQolhP84Ozn0K0
zPSGjX9DbEOL83wqT1wP+Kv4i5faC3654f2qYzYxhMu3j5bdgJOP8BJOGuaq2Ma3IzzvBBt74mOi
/wdzUoumMpOnhV+uRWiyyncwOIVJrar5Pc7W/qe7EhsPJNQC28751XeiMn+T9dTgd5K/rptOZqUd
zg3+NmvoS2LbK8F2Miey2bPgTzkKYQFgu4Evv3A/oLNFwM+A9bi/rjqWS4c8XjPFb79Hhp4PydeW
ZrXHC+p7v4dHZl7VpZx7kHYBswsO0LzEW2ylqvfsGdemaWg/KEXIIe5det4fMV+HVNmc0hydsOVK
6dv6dlL7vmUQCUfGG9THIg+Vh0QNqPuUH7KCwa3M5AGDqLUD+3X0/oBlMU21uo+6WRkJXpk2FOFo
idPX9aTjidpsmK8bG1u8DFYvgkLJ7GpGxxoSgLffUWwWgoNrk6RFyZuJffmy7h0qtvc3GKrHvHfh
OAsHAfY06VSMCSKlcnPi1O+wrKpIPOpKs923gFnsjrT3qPrWXWcg/KshcOp5fWPQWDYZiyGwiKQS
DPgGRsdbuaxa+WmIyOOiwlWRkBk+p67Urz4/9hoLWD9gT2emQ3j3Zw9fOMBp++zlh9OMh3pJI++5
USLsNo8Il+07aS7b5wKrkv5iTKJYtE1g2Ds8V6Nr0+j6gW2wbShntXvC3/P+ERMX84ybqzcLDuac
Zet42B/Zqufx52O6pUFxm0bDuh9XJw8ynd+QbWp2V87GvjekiSe5UW6RlUVi3Kg/wzM864JsXhUg
7aFoCaWEO9LYVi9rQmaA6IS0thOyEVo2PONnxL47DcEPQXFl5wqF8+K3BMxU4sm7nV1mYSLfp0Gc
7WvElTdhvNBZSQZQwy14PtGrKq6i4fRdNn3LSqLoFDR4+4IPVThAHo0S7fTUDTiZDtub2cqjsPQl
yyqWsMySO6ZBk0pdgrVkjT1fOb21bSyhP8/AzuY3EWhAlgGsPaNK3netbW+dJn5BMk2pRck0Zdri
R3ils8LNi3mJF6zgrhijWFWeEOs5sAED/bhrE2f5Z2eXP1pXReffbZzyQFm2txXj2z2u9Rdz2jxV
NiHxzOJxhGGMa079CjEX+fVPOJoclqgnRd0pJkw/XrMNr+oVObchxb8WrkhmzLvRDqFR6zx/UxPI
99/QFsoYv6QOJyTikmFu1U/+nb2GTpVFiK141OBHoQajcrylHW62LSVaXv1h3vQA4u6/fLjw9RHe
50IwU5mLnBLO7HIkl6Z6PoQ4L+CZusjUZ+iyEQrroyiw5mdzIiH46bDyEt253nzVl1IRpvXjQLW9
KMuT7i+Qb6BB+ILhX593H56xSgkpKXjnDpvkkvZXWgk3qGt0LsLU64xdRscOR0L++Sc+z1vRi7Sv
p/4fB/92jpv7YhF6jm5hB4tuubt5xJw1IIt9RBadPPVJI2MxIzyv3oVp4AOmxOd0usVDmoyjHjmH
gGoCjgiKlRa005OcS+dYrJe/aD5Y9RrJUmzsTiRKmiKwqzdlDCs/09P6Lhc52Jn1QGHDPJlLOzNW
nMvaLlXT0DDBv5Ob7PDlH6sYro01qm4UGVc/uicbaZexUG4t5ZPcDVllzJ8aSD06xFeg/ydxmFJV
/JFk8IJjuu/086Pu0M2Q92XrjRAH8lelmCxZFD7Gs5e8cpSmqD88WFdmJsVggmleZcNAFpIilNXJ
9cZow49NeQWhuBiP7BJaelDBw5Xj8f+anIvjTceFFlwFxstLYW4qDPCASFNqS3jXj92w/QKEDyHl
qDgI2Rjf2+ITZBtfa9678I7o9LR1hH3Oe8ES8zoDnpnPD9p8ySH26dAkrjegoOgC2NKgov2Ndgtp
fe2aZkJCeMWBFpeTTGvD5FBBdX1ivOKioz+oksiFbuMZkRdq06r7C+dwANcmrefdX15UVGqgTQ7Y
y0ntK18QtoaOcjIOyJcjie4xqEcb+O7TF2GABBhwZOoxcx4KPT3zwuSFqGRi6NJrEDAJwFKuVg19
m7pKZIdwzXc9iuRBhfwkZgZUFbx0o1XhNmxio8DCXVMtjYlLa6Wgqqwi1fxQZJB8C8yUVkNt60dg
VmFDXzv39/fDELtkmqx+/Z67JtHm84I6FNhi7mFEZfwjDGOwzFKB3fqgHctekEC2X7VXmUKjxUSM
mls9h1zxftPEomN4FzBHjzVF5hK1o93NUnlA0SIzc26mb9RE1pCmiTKzdL7gZEPCXfpnGmTHNiqW
Q/F99ZtDxso2KUXqdBroNx0niSd3SJRZ1PsN/uXUVcfrMH/bA4b6ypozQjggfNPN0kgv7o0I4Ayo
EQJk83sYK5KcuWYcSqccIwPCkkDNLDiOPKApU/g6fPxHIYYTzBmSkyKvgRjlagtk8ThnoyTjSAsT
6SvL4luwhr5WNUdkZg4qUzIGPRxhKxY/RYvgQVD5Bca3ILZ+LslZvyWLXcnJrE1IaIj5VkNbNSgy
aZpTkHcw8UdvsPJVlF80oUn/oPwnXBX6ZaNmUaslu6yVx1GBxNOKYaFBGLIFg0b7wDnVxwowu3LY
2KVaU2m8A/b7sIs11pRWkdL1CBj/8nNsTl24hO0iBjdMyQ2okblNCZ7y56yvZD0Lo8wta8i9LrsS
rmLURnk5VcUxXwVhJ7mWdyHaDf6QmYUFRUx0+SecrIZ+c9DNZjXtskIqo3htdOZA5NwI/xEDBZSM
mG7hYHTNtTorXI16FtmHlRT9nrqDRIc0fo2ZWYZyrEGaXaLH2yqr5RQ65HIbw6G7RXX27tdt+B4h
DihhVBeDcHTMYDxP4hEPX4zoY+JMtEdMGKK6gsF5v9lURaAteZhFSPz4l/o2AKH08FkIpu3BzOxx
Fes5EAnJcPS9f4wwCE1Rqvkaj4Da9tyhsPUp5Ro4VMuVcc8BTOg8PGXtSa6ls7rOsm+2RdvSRXmN
a0ak8lIBZVM84uWnPI+sc7SKK/YsrWcKYqJowHmMZduu5Sn6KaqaKpTKm0VPlGNDctN+FMItiysM
hsa5J15xg/rutP8/gRPsaIiwDFPG8BSpy8gy1sewiu/pPCalyYg/CW2Reeu1xlMrBF5PSUunsMjV
rrsZ77aFvH9rPFSpR/BQTdGB86JXv0Odod+TP2QJsiC0npAnOSByhqlrJbphFnJ9TrEkcosdmnmV
OqdOu2HnG204EcgFcm8ZyVLeOAidFmW6Mtd/Hd91Mv/mJcgXH+pYk0t3UARG07IxAgZxQO4mjOQ0
vDvmobuj9wu86QkN/EZa48lrUDCWS9GkvGPYV0a5GeqW4fjJBZ1R84zmr0Z3jIEefyOWjhXJB39a
56IbXEKbBARW9h6RHzHHAWJME6sSvRda7r3xDDvpQlSd8yYn1sd6IU+jv1zQ1jHbLXKoW/S5qKkJ
lrbCLapSgnUEoV7DNRHFTh3KVMSCoEQ15zFHY2v+qlLMBAFcLC0UMXgcwNxWcnV9NHJ4hwAygPSu
VD9g7XancICQXdaS8b9YVBRbIjkwrBWPehSSahlcDUwL2hbk9huQ2PcTxpjVfJ+tpGDSRMBykOPv
MeZMsX4BIGyoOYLtcLlHBVlwLkXrBAbBtafqD3iPA6O16rO/pz7xVLKhU6QudA1PcwBK30rkNDSW
fS4qY/5w35ZWwPJn+mZNbAZSicYgFcTL2wOKXfIZ6Ncje7ts13bpBh9w9657FieTLEV5cSJoHe23
7AlHxASMG4Obdnsg3qUoiT3JdVDpyrJ7FiPtuKTj+WyO+6HGcRlvnDZ1Kx8rjnu01ZovnHLOq+rd
2a/IeVYZuqrZ0NpT1LF+YZSspz4HSaPEjIaCptSOx1Nb1KD+1QlGNKjO4V+XWwyCqpPnPdCmNc9e
6Xec4t6ivmGmigPdaYDcKAbWCCQp2JV0fFJxAgBAWRkpBH/TAWQOLeZF4duv51nDHvnc90mxRbGj
6TExkor7anEbw68met6nvRixpHXSY5j0k5wf3NZRmAeX8NVgtTqFe4tO42KLu/KOiRPuM5K455CI
nZ+7Gtdz3/esV64uTgL1mu0Jf5TquGM1zWOWoUxPp/h1qWc+gESnFLtj95ObZFcQ9kU2PvxT07yw
xoM0CDYEH02KfEqs/4MQTIx1idBqsCektWpPFcAGSnEHDkmese430Xnuq2u/2rhOPY6ERq4rTqGb
tfCDvqUhSARreyYzEJSPMULagmv2m51JAkxwK3T0ISGigNpI5Pebs7sjEB4PXsJz6aZYvjIFXHZJ
taMDK1mjpjvybkcmB0cTJuO188QrhHjDZaPPBkNQuAGYQDKeRwBUKmA3yUq6ScxTUADKSD3igqzU
viHa3XDJLaIiEAnRMC77RkVzOV/h3ZTqVLVn3tPbYwrTpx73xus1GRVmzVBBTQSAn+X6qMh94rAI
4RAE6gHjeK6qOD6tNCZY5qT0a7D13/R6NsweL7sM6AVqxF1DMsJKsQvsVbb1dRI5x9jJLXOJQwCw
FYGKzWt2XALQDjJHWIGKXLrcYr0zCpL30JanpMypP/p6IbTzDH0fsSpbz5zN8lA/Iyw/buXy9y0l
ktbsxMesEYyO0bevbmGh/RHb0tgFU7H6s5fVC8T9WujSk9J2fDwBiE5F6QBYqwXxZpnPeV9TFfey
iwHRAhjkSxdrMfU3/ql3MpQKoqNMUSle8G1jtcVVhgRQ+ajPyjom7J/R5JULSBeK8tcBZ057FRoF
LQrskjWFIVjrV2YAhIiMEzKXl+uXZmqbUWXDDVa+W5CjEALm7C2jYDP8dF+M7CMez0N2W8Wd3hxw
MI60oTXTOuePVgHXvr0pM8EEMEglSgTs+tG7vWv43JI5ZerQazVtdqEnPalm8EiR5tZjETuxIj/j
etBvR92G5CfD75I5ZfiBU3VCgcwCIPYAL80A9JWptFPRQOk53xcQk2ORlL3uAhXAJW/WO9Qs6Zjd
jcvu5LrPN0DqfU+1/ntbTaTT7LpSQ7jVgSOAZf5mi394cIWOr1ZVAv0LbLdx79Z+PtU76i2L+Hp2
SD0QEUFVmEkUSZipooDUFD05XgMqQcIIO6O7GTSjC6M2TwzjuC9A+gbS767SJRFJbhnfyavKOLn1
ZTbHOsWx/NgdvgZzH9JdQrZmdDDCcWYtxrSUyjOhQLa8AU/ttg/iqgwh8EfMXYoywGWW46BXLJyy
YOQ4DwZD2nExvmVCSg+Gy1HQKlRjwZAsQullK9RFRKW8UqKx1aJPRi4vER2asb4e7RVBYCJU403i
nMeuer8JpghLix+XO8LT/jmUNn9nh+JGeNQponFV064ZcY8sZlfhH/1fBCXlO0CXqAiZQl0A6t0P
QW68MmT00pUZkwGnnRqlwtqFcePL7TVI/BTJZsJc88SXaOBWOcsvJu9sny0vuxDP7YIIMYqgRz3s
Q8On+slDkrjs4itmX7gPZsjmiOn3U4yFHK0ljPALR6bPiW5H0J4svu4DYCuj8XZguY6VgKnvujtM
Hzb1U9rdxIfhF+h0hOpKSZ+OqJOmP18L6EUd2TOBSUIcfos9lnJ0wZVHo/pKcNqsJacFTbqhUU7O
+iJQWf5cmmZwgHivnFvJxOtiiC7sDolbidD9cNoXbP2vTFJBIILmt/ZiomPDJ0cqLTE0RG7uBBHG
YKnguCMuce4GO41J5YhtDFGMoKQRw2gesNp4MJ0kDskIbzDu9XbPXweUUCCBCyOvnHMZJ8yBybM3
cyJz/BWeHPGfnuG0mAkKP2hoUCtNs5D1Wu4bbS8JuLuUwGkRl7yyAzdeSKWkOWySjF3j4ChbtQeC
POqJczUQuy/LcHQJJXSYxGJhp6Q6nVHS7kD8Z03gT0KBUkzkgm2/HprBDUdDyxoGLGi/cIEL5fgE
OjjE+42EsQnPBun/BTjqc1NqRwu9zUxbZK/osRka70EfOpP6WZ+bObOgACHqQwmoH6fOWFNyjTc3
fGWNQKX64HSByf/STRGRqzIaOvtamdnnqMpDVw/XMNjHK/V/xkeLPoUQKHD9AxmTPWhTUf/fkerZ
XMyBzohtQj2QDIViggI5bowWwyD+bSRUNfTZMHzF3JpM1spK+MFY9QmaPDhx6+vpV+IaK+XiR5u8
Tag24Mn4R4UA7ec4pbEj56lAtqujTbEzJkw38U524bHXM9nt2Zkm8diUkQ/Uod8L9wkrpvXzK96b
5qFvhk8yjydwPP3qNo7sK1pVFqr/MPXTVAAzoLkrP4+Muba6IQBvHqj6InkS8FiTArCR9cNHU2eB
+Mv50msuGc9TIJM1J8vgnXxnfVVEAr70Nrsxf92mkygb5DLW5Fqam4Ggerh/0JSpy5Yrt61rrBmJ
YbxHqnjVA/j6YFLZOPjWTmo4muZBHgw4BckCSZTa8fvJCiwbdzBDxiQ0LtO7x+GBJEda8Bd181MI
mBCK6caL4fkJUyasWgr17KpYfcZwwxbrGigl6M956V161xriE7Pf6AchNvClT5f3gyNH7wBsRTIi
6rym+EKj0XuXS3r+a3xOMv4RmY/EXg6nbv5YLqpabikAsAToco7PTfy4SBvglV3IEqu1F53gEJJC
i7zrslHyd2yK2CcT/De4HvtQmc9/r2duFUEZjerC7o5V7e+dioqrheLkpibMa4Vs3DdsT6ZjEDYn
HpN0UGvIie7t3SlXvGj6dhzfceYd9v5VCEqKmww/zV5cFLEmggKaNyKSKI7GU+TSg0Zyj3je7fTB
j1egj00ec7Dy/A+bMU32RMvV6z/QNGupNiZQURsEeoQ4dy4cxY1ld5AjzZBJFJ1IBapLerEoPSoH
Fatkh0ooEEl8VNSp9MkXe+lNn7frelJH8wii31GyWamb7CgjdyoFETvBLPb7g9bpFBQnFgjRP9jx
CZWmtYEy4nUGcT9+GCrPzG6uRzWS2MaZRJRYXF0dsVEdozgGTAFxUVyaGpNg85+N+VOtBEM0F5ba
roYh0r7QHnXn3CLk33a/KddArBfE66LIRI00kn+aprVqYl/bZVYHdHFpgN1cNFqmdAE99kbMlvYJ
n+OZUhURzHdU04tXjfHRFCXDr2YTvMoTTndlXiDr1aergGc1C4M06FLAl06HWmxOJd+l1aKpMN7x
3Q8siAaPCA/AJPyjSoIr/NbLWXxuI7M3nURby6HiitdrYhOJIAXBDc26KU92OsNeiDnlspuBxQ0x
l0uiEevNCkFx9T6MIHzFZMe5PpKOaPhgS+UHDGQA/OsPq0Q4GLYv/nXp/tk5ypT3DLa2ir2zVpBC
N5zuUoIWb+9YONf+Q2Fao6yH/LDll6IMQGnhowitvceSohP8o5oaTOlu404OiFob2ZihTBX0kXCH
7HWJpAJvZFK7uOXIc3fx5aoGxUWUTCVWBS3muESH04mh0gB2VBVdIa1skS1UfdEBO3xj38zV6rf2
NMseV1iik+uOUU1tOoJARd3JNXcSwRXZpB3qKDyw8iIu/C7/oHn8mj4KJn4apLkwvWfo92vdx3y0
ih9kwW5wK0QX7Oz5C0veZ1Ql4ELcAZq3hUXB4yxKfQiH7i04uya4zvHHCniX992pTp/Kn8Jorgl3
r73fS4Yg/2LmNIqEj465Et9rxa9+8MEIO+1/SeryN1UFuaWhWaErk4d2YFzeTcZHmV/k5DHt4Z21
96jynWFMCWM0grvkpsjjZG3ttMseTW5/+GdI9HQd21iULXyCtJNC7cfECZ7CI0uVj7h53A2BAyuJ
8YcQMXMNV0OVIXGijwo2EInYTbLjUGdQ5BJT2eYtw7pcLoaxVVyUlUOzyxKJoF+M2dvwb71Y+caf
2ziUbnG3ZE4ZElTR9wDcw0etxerntxgZxbyWyqhvuepMq4thOdW8fD7y92ysA2Jv27YulQ7Ruy7f
pD6BFqrg3Y58LybTUPMbsO7mG0v4n/LDUEaghtVD7QGNUlxXjS976VPjoNVI/TKRx1+qRVJK2Av5
rH35IzdQu+fGbs03UEaKZOC24L8st9FPwvi5xyJEwCeqpg0/3t0vuvAcCim/o65VDhOQ3LJo+rkd
+kJhRfou7UxT11TPBvL2oFsJQM+IZ7wFRdDI5YpMTv16A7D7xPVXl75F+eG0uobpR99m66GS9QY/
vFsajmQLNH+X1HbH4sSbhnATOiruOqZ7l/wYVypM8IcxDFMvEcddxrLFN1JYiz+vmeHm2Ons/n1B
sPchH5dpDTcRlH+rJ783jeHTTHXga85rXmnE0E8f9Xgh5IVy+eArBc30BJfa+bgxIj0EKuv94r3r
ioN410cqZrMIcdSixeq9l9yQsXcgIsT9Ld8hWyY+Pwb3XYonSo/zbYieOlR42AB/ycPzkXHbMqmn
nNHy5MTj2Ti44LdwvUb7NibXnfkWaGpE2OmHawVs9n9AYwk5vqkTFHRwt+3+ZT41G8umEE9+MGXq
ddtKr9lJbQbHF/OXHMwFsqv0Z2hYPNkdjWjzJIhjgeHqxtXEo7GwekgJrBNI7mICjLek1F5SKcxE
6SGE5JjVANFW8440pVsbGoI+e1CpB4LOxsTnSo3u9cjZogs1BWOS++BgWX3A0uSgm0kizTMPjSl2
UapMWQzCG/fYsddCeUg0uxhWlxrXyzLBc6cBM6DpXGnOfdSwcUI3e2we02v7HKVILPRtnx7pqCNA
Ol/uL4594l6bFBmACC5DDdpoZbRq4aVAR8r4rt+rJVw/GcaGFciZ7GLoE9sDUlKXcMB1lcS66tCv
Rn1zDGkBG6wYeXNoNBsivvcrlfYpm+R4zgUD8UAJE956g5dToudndB5gycmP06/TX+WspoHofe2Z
tdQkMIB5QKE/LVj5cJkK+nXP3TJpl5yCT+oYsppiA3kJ2iylahQtoJusKrdinJ9nZPxgeufPAfwc
/NkzB0uBz8NcUjHoau9EP5fDOTw/5KothdR2e7lAva7933/SzcJuLGn647OnYRzPlEb4auItNOOY
N79I9t1OLY5jC4o45h3r5SDdwXTbosJklx2YYyPH87+x5U2Q99kzDrR3SrqFx9F0QGvwgD7o2CS0
bLyi0oxZw2SwbGq974bdX1yHHX8n70lxopoxkQPbwW/cIO21RgcZP3/5z0uyQUzpqXD1NcIt4wDP
yIBu9lMPwk2SW8h9D1Z1pelyGVCpmLILMRkFxY3MnXIrWXBBhCInxQdCLDYXyImansXgWx5lKheM
iADPKV5Rl5vP1HY5woSNPKtVh91FKl4FqMIBF17si0p30C8uZn3h7rxhRv9aKxU04VzDhpSD7/A9
IiVdpwh0oeCpFrZStjBTQRQYRJHjkErL2rbdjU7W1iRkAEtjjt6RwgOQtIBoJP4guTw98q7RuSuO
rnsSWeAWatKjhSsyqpXUCBLtPyytCRkcZURptDVJSgErDks+YwMSUqdBBbIsjvmZs+99jXp59ePG
XqCxzuj6jiE6YaQkafzT3PiK6Y9TwRrVZCTBCpEfBmSrcMOleD0EqVr9FyNiA1TR1XyIjSHjJusu
NpXhtpgKjY1grHR7NWKQYbI3nBncKL26whKNywivUrvmazFvgzbqhIZDfDC5vZtjoPFeyMV40p8o
60nWRYt2Q8zwZEa2ONxKjB1TsdtTcBAC4morU5mPNDAiarIXVSbHN9+qlXWM2xxJAp8BLV+6wFfX
4lNOn/PH4jFlP/UEdzl6p4vuMpsCWS6BxyeR55UGUhtdU/pPCnRvmOSivQAaWIeeqNXxZHMoyD0+
ZLlGF3qyZh62Xv+CwVYpkSekQv67yjY/zUz2GpMWlspMj/KfUzlfQoHjddTIRV2VK6xLA8PRXTFL
1+jqx12zlqVkGnE7yWnf+o+IgrG6r9Xtt/vg66ZKAURBjLxWLIEP/KtzI3Ae1JMrSuLVBgLRyS56
VaY+138Bzo1uXREkzzZaG9BLPjLmV27KqZyHaaiDrSKaQsxy0vwaG6IxVA0T/0zGgFG0XiyGdr84
f2lueddk4YOfivVYDG9ecKzZSPs5sb+O/uVAel+Ax6y0AZ4V7HP1D6lA7WD463VgouPKTuR16naJ
zrKrY/myCwaPwhE38QWmg0zHyAVzmkMGgqwLAd017+EEadSaPt46gzYIcn5AUg+/e0al+Nyr5ZKj
nsPGmoTJpm9tVFeC1ZJrDANZ20GV1Kv1I8rBCAGU7eH8qC5fJf0RNm+Z74h3A7iduIjS+xodG3X4
5flOZIXj7BpwcQL2bilghpL/oyIYTp0xJUhy1es7TiziYAmFHhk0ykuLwC7z7Jtq63tDtE+Tuvpv
ZzOmz+/hGNck5k1lSXFTjWuTbvGxIS2MnFz0xUv19sx7PYYDjuyWRlinsabniZOgl9aOX2sIKKPH
h7jxynRxHMhTWGVnsztnFsFhZTe7Kc2zc8j3bfGRrkAdlU9XPUy8JeJmtf85pFpyC/lJ+877/0ws
tAAaAB/dgXUntGVrmkDSbI8NuQ3M7tDKhIfFzU8ObjoM8KAs7eaPPRR0L/rE5McrpPIgutPFv6f4
KHtK7522bzB/wBqaO1n848dLyxlYPRrf34Q41CEHvGKdcbooxR0ZQe4ccBMKxe/3PpovHpGz0KCB
HHWtJYG2UsJLWhFEuLrNxryRu851+gOSg/oZ0X0A2pZfwTUpjAvdTlG4sxSEVWR2Rzh6UgUvTC8O
Q2iEpPZZ7MXmrTSGvqkZShZBrgL2kqJKZtw/IWUCTYlwYCwWY9zfRFkFv8k5WjQ1AyoFIehdf3nc
LnE1RHBjIVlsSsut+ny9vrt6pQhCgWuRRJKz66rMCLY8rgF4B/IMzqYWu1Dz1MqEn6G72xrhOyrN
0UagWmg5E3B6eFG+AsPDDiJJzteoTDurj703QD2SR5XYaz2V94Ozs1WhSWVFwwST7NY2K7QYw3wd
iAkFLZwlboQzAf5loqtYrgCWoRVvqMwljhYsD0zssiiQef+Z00BMJGHmlmP+YwNZXF/f0NUyss7L
Za/fHCJYWBepx8+soDHcvOSF3qdgW8fsS8XQqGbxTO2RszoAehWH01TZDb0MKICYCVjTYvhm8Pi+
+3jAE8aN01qnoFmvzVlTcIVluWKg1cxkzr3b9BzvWpUlkrWnu9H8LrDl/SZAZMbY9y4bjhCqkU0Z
/zxiqpMrvo9w7MhEimRjwUzl2aEAMDa0sArWhmFoOOTSfi8IgkT44OiJ7qWv8mkG1sCQ3qFw1lVc
b8O05o56h3hj5ftP8+Nvmmp9Jw7Mh5+MFxEOUrtW8Y+vtpvg/EzHBD0pUA/VRQZOUf/2FzN+6/57
Luwxi0KtlaXXQp2DJeRHEiF2Svf1xzpLdAPStnScbGu4b9c9XyyO99ppsXwFR0CnBJk5LMg34xEP
mnh93Js7GpIK1CPaCXsfxuNHMHPKdogg8UEjztLr828RG47IwVbw/GH0Ahf0zYdXhqkH4FEoaAZA
Gh7ba1FDnTqB5y5SLiv3fBfAIMSEc1APFYjNCfWbhE7JZxEAq7v8pzRDKFgyPhuHxM1CtAI+SwMt
bAFE+Ba+oT6DAND/b/de3XsKm184RIfyuVeHIFxh8E7lLtmip8ManYlw1PoTrT2Lx34v2rvhcDlf
Boax1s7vhTGs37e0kWDMOH5CEVuxkA2x0u+IwLS/ovqml17UQjM4151kP7+Wjm0M2264CgatKvXU
zda9Csfp+du6Iz+16BEqNwVj6TylUV1V7YwFl99YakfNDpy7rLfCoZFgzEdLc+MRkLCwSLeerhgc
iW/EZ2unJL59txlpP7vAxrZd5y80MjrmF5yTGMZas11XR4r2PKJtbe1xdvoCevFABcKylxzwcP4S
kI1+ThnUdrtgwVBJ3rSdM2XXqoPg49+ZvWMQdud2AYeUAnLCeL5V7o16pMn0cIk1cUaBNlpzl92m
hz/uviXo9u8TAd9WKwM7n6ajd8mCFn1EGd2dx9Y0cHP5HzdI7Y9P4F4rzdCeckUEqpGWIxsxWmVW
alBVGyeC4DYthEgCCCJZun/lkaQqiGj6OHnJF5JnaOTt43SoRl8OMumbzYR2PTpw+3qVM7LYfWBf
qtCkUNzq9BrZ69nAGJyAJCSvR89GSGDnVyL6lfMv+Ddu6LEAo4Fuk/P2QZn8IIH2sVk//s8uBLL2
VUun20wmigjyrEkHFlcbN8c5w+7n4H1Tfuy4w+w5ZkWIs8f2tPFpRcbD7B1NgjSndYb6N7LwdWC7
Ko8aSV0l5NchsKIBRgcsy6zpI7EA4kPYxV/C7Q8nTVDB+DKzJGIuCbFt+tadIgsNnZ0Qh2VVNC4D
//b3UVCGx0nEl+MBoQrkVcH0WONfuVXTpCgo0BNHNbEQ8VfbxtjCVOT+7iW2QBENlPftQrfxInZE
nFxJez5ywiugpjQfRoHfMGDWii1sbIABZvqIQIeMlvYvG7IxZ7E/DkLl6Dy/PxYIfmUvGQECO5Q0
53E6sGrfc3afNT9pL1XUaiXtHUSP7Tf0hCPZN1+XGDQjUQfTVBiigbuehwR088qRU626oVXyS6fV
xoruoH7TwpLysIW8VcgindXCOotnDDOnH7pD8lon+WcuzZ7t9LWpyyr8UTsvc5Q5iu9VnGPfkUqu
tBJ4rmXaBrp/L67YjuE9E8fG72JBSYaiGP/s9FjVExj9YhTmWn8cMYuRxIhTKbjFVECazpc8xcTB
NyBOwF1A+nY+j5rnfcRX9l5hlV1jHkuvs25J9SDv+Kng5OXSZHDSCzuuimSdrrTZeTE63JW58QQY
xJyXTDMLRClb278HEeJ0DssolU3JXbdVfRWtiujqh1r98YfhyyTedcY3S1EWlHgwqWQ0OeB8cL4I
k0YNsgoMcAvY64KuoLD71fGbbiDO1BcTENxYX9bNxjjvv2EnSZyL/f46GKo2ek0ULRyRWVIyiLHO
ZIQdJq90n71ABytdHkCsnEP60OMWQ4rcOVpT/u01hEN+X6OFu/Dy62rpW6y7o8OxHhmjPrJFLub+
vGKn3yxRaKaXenI9SCsRsrrpfy8CK4WRTDVbODLwYCeUKTCBGHeZe9OIhqQ8d0iaww+XXXQK3F8d
GoRN7iUXk/ZssaNsvqsSNunsKNJJiT9T1tN2oHvE1Iz5R/KJKJ6lf4+cGKkcimrEovI9zt+hDUZa
eJPDWPVRQr9dcne40/ejoOG7ILiO2e2piwmMxfGMSQj35klDeeBX7Xsi9h+0m9g7GpIj+ARvkxZA
ALZk9gJ77hxxeTdxcKwXut1yDqD9NUFwOkF5kimiimCtzjuGz2PiHTPL52Mq/IW289WOv8qKANiK
CMO0j5ONUzZAhMUbpi59D89Ju33AvOnk7/j+zHUVo9zrx6eCzETpAEdXt+diT3HXOS580jm/6DDt
MciXuLa2wVzg4pHYaY997yY6yu96iovNPvrIz5LTL5dmKFr1tYmPXKtsbh3ArFvztnZrwxLiGrma
8Y2x92aNUSwxkvtAz6KI1PjMO/WXscauGlnveiLdLlzbNjqxVs1yGVdk82GEMVgO8ardBVF/TzcD
9laBTJDFxLGmPCuUcDxw0mtZabjRcPpsBu5nWNpV7ogfxAZwdy9FyvJW2/ugMzsq6LAyfutLO92f
6/Kub7zcWuaukDITBP1hQfEHs31Qo3ribhRt8S8e/h8WC/LA2wjOgDrBcUCX6hZVJUjX4q4tKFTS
2og+sPZ0Ny9yVreie0abBfYPRuqo8fY8QR3X598H3CyM4KuV6lYFkfoJauQfAWZKWvAIqs6Guwmx
Vj2fekaZ2oEyS4DSrUrCWhuoIP36h5rAcsySB3EucW8RlTsKdOJTvO0zT7O7ClPtbqzndifcASem
pMATXgZDWdAnT3B18+yYA2nM1guSc+Mu32yNLujP8/6Q90/HMD/j4RQDQ2kw98xDZFcisY4fJfez
LRQCm80T1RlHYbO3oUGTkGmR4Ys10EKtM9UFIqruF3DOBY11JtuE3TgAL2DqLtciUymqZKhOx+ql
cSB/rGA7Ev0jv1lr4RouRYVt/9LrmtC6BdCLTEBe/8uL19b7SlxexCWrYw2E6Q6EQwJZZBEeOd/5
CYbfNY8PMT2KbqCJsrplOc22Mo4nO50RfjD7f7bGxFzu8nP9+OQUJcfeICqIUoQBu1W0Dwqc9olE
5yKiOYks11dxZ39y46SS8YthASont5ko4kxOxbhO31f+wi2dlLqravaq7Ss/rFrV2WwbG2SzI2Pp
swdJ6OWagYUcnJ4kmdqegANIqJvsGNQlOCJ7UQLOHjJs2NjNXOmORO2Qdq6J8eBm8vOMsaDoVdpq
zC3XB842r9Ux377dpN9/dtpbiWxEcn8T6Gb51IBtp98y2jM5oGyGcavDlO/5aWAKm5uvb+2Fef2L
VfUWX1P0hlYw72cPn1aSJJs3k9VhlJPFxM7wFHvhMWbl3w2GqYmDgDWlVQALEhSFBgfQm7pTkA/4
nKzLXz3wycCiAsmQFsXSr6tyVZJMJLGlFt6U+K1GcOUjfV0Su7U65j6OhtlTcktidOQgOyAOpYyW
QOmWizIBc3UZdX6WisP3yle/uNHdyuebC71UZzckZWMSh6A5GcKIVkn1DvGMFf3W5KDIvi5PAYi2
ADAqStJVvb9HoIm2l8PUw3UBXe0we2equvUglgXkKfUzt19LVPdlqm2BtCrFZu9Y/plPrpA7+Qrl
NP6yo0rsg+4UkEO5UXqx6uMjOs3I86mDW+bLyCGU1raWNyPgb7K6bCZ9OPA/vy8toHD1Pygd6lh8
MQdD9GyJR8t2Jv1gyO9sbS4RfV109pBdcDfB5HGXd96VJo3MMOiMYSGQjs8jUbedi8z8DEWj3q8e
SSsvtyWyMcEVJn5PBPg7YSt22RQXWI9rdBUB/fN8WzLN+gPrXIkwtNxwyzjqT1nKT6SzU2fR8Cpf
UqsPgO7rmdQ42ghRKxvOfBkfC7H9ejCF5w519MvqYH/jJd5VsOJhOK97QZ3IPHS+mUQqR3ktjOdL
+l6OpisriI/WWNKMrOZEx0oofYNkO79clKCWY4VNe8BprNYA8MBQCwlzWCEJmwc8nNVMofsRn4vE
y1fUiJk1r6XNzGSPqMXU4qPBwVmwHLJ2yen6wYh9dMwwqDmyXGaMiGzmI94ewrH+jwp1jaTnevao
A/JJbDQesI2P2CjafkyOWjgJUMRSX3HSr7fK022x9UFlGeXQ4LSTgNvRyEWuZ7hJ6O4xrpAcUN/2
lxo/Hhqyec3IvoebL2s1uJ9QUD5d75c81C2rOb4oT2AaVYnwZOouIwh8JLODYIm8sY0scXTbhcvo
HjK6sGF/QL/Ih5jGvRUHMs5fSNIjkqy8HZMR7Xpj9oSMZRH8rA3SzGUesMaqRGxLkcP5z7V86erb
uJI4HBaOBiQdKrR6vONJr/zcLr2Okgtn9VsgfyYHbSABPiWYJEWtg4M62oCVE4urYqpcme5puKdJ
SHyArc1IWSB5YRGbffrhllYs/e/XpmhjF6ACfSQhP78m1Cg6Q5lSiqBORu9DeYasMQyir/ETYtih
sMaG3gBC0X7/B3mmGvQzXas/+5z+KDAxf6ZGbCctnGwWQh7gx4GN7+eA7uRSKrKq01u1ud58Rt+M
QHamyWypGr7MoDv1tgH8xaOv8iQ91jAul79rNxo5f4nfMuhfZDkj2cmlw1tmednPkWlszRu+RxGr
R6ztopMSEOm47SXMy2KzA018nrPEyh8mONfT6CbbMEevMfiKwlckFTIZcrSPrJq/6LWOT0C0sH65
4BgfopYXYlWEPr8xMTx703mYyUJY89pPnZDJ4cvJvcbfaSRiHZJXREag2+Ivv0CL8afpFCNRejI9
7Q3TNHXPaqFESAmHHRi2l1wE+AR/ZMuOx+OJgbu95ZfLQfeI9yai/Te4HkluAGFCY565Kw6bscjC
LlysXH4arjYAzNge0yI/lgGsNbv5SPqtjEQKOnuS6IDQjAetAUKGXT7fIBkDbmwn31x+CIT4SJzp
5RCg8D3ClBzp9QUEJ2I3LL1uppBfELa220L1FyKSoUxG3H0z+5PskZRsMRynVs8/uEsnTk/1A1E8
tWGW2CMcpn7coedCVJqfKrKqnSvSSoZBTnwIWu7beZFxSWAlMNuJRoaqFfZseLrNo+QzeqMvq/vd
Qtkv67ybYiu3tDW0NYFodQs/RDqvEurgKcKhwP0KyhWPf+EAYNNvZExjPlSB0dCLFJ4nCDDqZ7kf
cfEFb5lHBxqgoHdcU2bFGby8HMRfA4n0dr6yyW4HLxPsA4OIhzaapf6qGRaQC8o86HOHSTX8wlSo
TVc+3+dYLiAnkIJ1s8UsjHLZxngfyGHzOucVzK3kI2xrcH0esMhhut/PFoY+26Zn2BLyhEd0aEyi
PHdnOyJ0ARc8jyBRI2yjscN+fQaO9MOIzsdBUzFT26btw4V+o/Vg5aE7VKkN1mAr7q8ZiZMGYjc1
Xt1lIBR6B0UgKdQHnOeOZpQQnleV6xLmIxbWiqjnoHMHVmZr76IZ37NQ/VgHSs2NuHeWxryeXb2V
ZVNWINXVKcuXS4sXDHLhO+Sl+4sKxknyXwSQVL1+T+n9c4xqD6MPWzzpE3DHy0A3HO76B8HuuTNA
vhrcJly0BTpOk+qgKwmtIX3y3KJQc33rlnpDt74R5c9wou7WwOd7xA6XJUvdBd258PBRoYIQqrYZ
yP/Kwgki/dajtnlgWBnOhDP/A/1TTLmCi5SyH/BqPMR+Bbe+wHbqSnGIhJKjth5I1nnj0fCrYhdi
ytrl29nGcE9zqSh+2BQFnl4nbWDBHqQ5O85YkR+AMTFMhQj5uCfvrXIfOG3WTSYDPrrJpZBD91fb
ZNMpy8XgfqFdgO58KiQXz3SVtGpVbrkrqQuk+D37sp+oti+DPWyWf2PhyJPZBy96WnFX4oVEPqVz
MWmuV5ZTuWq2cawqUmXChApkrLjy+P+FRobvy2w34oTXa8riffJSDtRzYH4ZehhRpRV+/azo9Kw/
6Bq4XCp/6c7W4m9w+f8wjGnzmcfiOmeAylYZiCKtIl9jY4Qb3QB9pGdcYsQ7sCeyjmy7CiOJqxVt
h8kE5uBUQvTHz3o1d/YF3QvJmX6HXvhXfkthObmLreA94qHfuUi3XNHSdvB5bx8keyw1rx0spVJU
oQxP41rs5EVbZhUZL12LYon3B0+eqwf/4uymbZhyPpf5qpNarJ/iwSa8Og4vDl3n2dTPGdTwPUft
hs+Pbbbb/nLb8+fcCAaAycWFoAjuDE9REG56vcUda/iQiG+Za+fokAq4b9Bql5YXIQ/N9aIY6hNt
CbTY3q7XBCWPeJV7P0mRbDoB5PhRaGCCBXKvpKiDhMdfoeEbLofDz7xwhYVXW/IehQ/d3x3Ki1Dn
62np6iyG8xOJyblvUGsnCxP3E1daFHyPO+3kSrEtukGecfNh5RO+V9437Seai4Ou2g0OULSdCzW7
Ak/GwTG1I0vILqH4vjZdiaYq/txnnqkNUlOo2mE2xClhd7TLYwXnt41W5e1/miAM/PONN2viKNz2
cLTEw208p8tMt0z0W6ej1TjGuY8j+PpA3q8hAOkijad2gQ9Bv05VNl2o0hIcSvSpPjQo864h+/YP
mYincKgVOQnFKW2mvnTchoEvRcZ0NuS787hANAYEXalxmbzEINtmy1VtsBUFLNc1lPxaUKpVMu9G
g1z2STy+LqOtyBS9XxFrAssV4NBVBq2V3jN4XvleSVZUM1hLaojIAxAtrSSqpuRJJmIQSsM5TVIR
AR9wkEStQm58sP29C+ERha9B9fF+z3/QfJuVMu4+cdbqf/Mh9+wXA4QYpIkGRdJO/i3rrKDp/5In
5Q2xXiw2X0+PjTtMtUPFLczaXGLk367HizFE+axGVXxP7ujf5N6zIm3f+fRupgNz0Qo2UyskG//f
GiXxe0dii/X+k1Zlp3OQgNLxuRsfCwZM+8sbcXvjdK6PDdGs3SXyuSy1J84dEqfieLYXok/1hWC+
Lt5qHhl7lfqOGS4mkCX6XuZ3dWumIPYzF1GggIfgQ89qEt3btC4Ox1xeL37KT4VZBZfpQpXEscpQ
4te0ovc6CLwJVug7ZKiSot9uJAGGBNtSuUL+icZ6Mu08c46umen3dYERK1u+Tz6OnIYWs/KOJG3M
DpepWDbCVVZZtHCW4J7WMiKD43HQAP1sr3lw/FFFYcXpOHbWEVAfjNwLNO7NQg32poNqImovT2to
LzBpJsYi7DMEgWRkwm4/1qu98oKB8m0Lwqo4Oz17ujx3QhZIe38SYXkfQ//HYgqIkWMubdFNN5jX
6ZI/5s7vTbFuNSMALXnmB16ToRn8Fh/9G76oFTVsjc2EUbSopYw7JNLUb9Pgup9ExFXwI+MGgWAk
pImyEyicUptFx8AGwDy0VRdQOvxPTFnhMLXTCYq6vic6ACNUQ16AQHkB8rlnpFi2q0OizDB+mgX5
mUWOEkw6tZQBwc8uD1iLGBJkQWDIhyHFYc5uK8nVOhL6O/NqRggUdfPp6eY35QNwSpcErWvZ0QQU
uFCiVg+4ijRKqQgz8YafzFpcG6rYLYs/Q4C3KaP8pm9D2xB/giRW2+w8NaUpHdurx2lnJwPZ+pws
gMzucvi/Tp79YIieJt9oN9OFqc02duj/oK7e16EWG3X8NVvxyE0lwAm64UloHmw2kuZZNDuLhYZV
QgmhAIXPZWMRWY1vFDqbPBQJ3hs+599gRze5gD7Ux6LAA+y3OKrQhViCU4UcLJbdTzqDHYvxilxM
3oJle9pjz6h0K/BxJ8d1maB7I+Kvi2WvPvg3hLESUfHixKZ5DzfgeNZqNJxeaGOVnZenAxvQ8GGl
vJsFo7ChqKrHNnqQ68AbcAuVLaxEuQLl1OoaxaiB8pgp92zYzWc1VkonQuYlalT3UKCTzDqLMIWe
DzFB6/fmlRqOhxn6WklLhpE3bs4s6Rdf3J8hHFcx981s31ZU8we8AEbotCxKMCnnl8V84CstJ9CR
ZB5EGrvfpL30sKPACpphJti9P8SEzJ4JurgMFYIxCgAUe54HnALAWjuyRyJ0U/6xnXtT4x9pPM7K
BkjyHZLRz1+9rxHwuzh9EFoYKbWTp6P7afxbrGbaW97qpTGSItsgWU09BweJJjU8aQRHGOpuAopk
nDKz7qXdaeaZFtb1p1KJ5rk3+pjH4ufXrRlY/H9w9DxRkdD7iZIDXa2HPI/fW9p3M/riwGnFU4Mv
LvlEHD52dVhpAK4a3bVpIztExI7CqqEuyXYsKB8JfoDGI4/uCpVDf1flC6grg9nTtpM9J9XDJGnV
MFSVkgYx2BiD6kkGOP3QKIufOVAAP/L4KDI72MBah+NCTxi2RERO2P4LIqxeYROCgGNyOD7oZDIi
kCIk2nA1LRvLSaoUt/thieIT30mbpj0av4tc/Lx/Ysgcr+PqTirIkyp8Vt/fMAd/42zaQsQ1CuiI
Q74SxWTb+SpgZ9yG8Nq9uONBBhdd3sRQ5yzGpKOJ5K8WULiay44BEd11Rqz98jR+fZnMUml3j+zt
NUt33E0vEAr0lQapWF5M9kXUscnFq1pCNQ5TFPcwfntOA5WwfOvEoy2U9c9KH41mRfGrkbDEsW8c
iAFL95wnczd4L9Mg18/9n1Z0WNxbfc+oDThtzmVrGFYPVVWmrNfe7HVbzHEVO0zsy9+ZEZ0EvPfQ
qSLYk6JqYBWKtShBb22ZDaUP9Av19PG/LDMZPcP12UW+M2RCNEAuXWUIu2G+2bOlvuc4Ige2F6eL
5cOa2HuCY+fjPCDAGiUscxeuX86oHrt/xsLWkzh9yLmn5n4mANgyfvNVrq/Kg4P1AfuHzw6drUqP
0ilnvCUxLu/5iZp6CZ/MoO+YGBJxB56m/2QSmRpw9BohEfdPwxgggXlrpVIGTOG7A13963K56sZJ
SRc1jMqzoUtbHriMQUn/17oa7IdnyeA5ojieawXpJ0HaCgmXN4rM+PniuhJ3/JCzVVpXaqx2GmAV
CO36R4zupZFfQko9n2vmoMQgyirzY5db0NJXG+IVPXnXhX6YuynVW8KDuFrfXRNL5ItN9YV55USc
vDttCUC2D5ZI7odwyt42o1e4GfBomhx9TvMLH/noWjMB1aYPq3YU73HsVgrC1eIs0JAbXCjxLWt8
cegigCgtXzSFNIMBv9+7qkaAXv0rz/kVHZYYzkbn/33uqYW2poZ3ODawz2OFZ2xi0RiF9jRV0wYy
FuP5iXWR5q8AoSK2X8JuMtUU2NFLerKXbkXupB87cOcXSrF860XUA8MnoLiXwear1xx8klfHYwRO
LOOCwmXexsAEymJocDelYeg+jU/fRp80hyZqdPyj/lftq9q83wS0rm3e2L3gXP7gjGjWUjCbuPDZ
jc8QKaTpDyM6muBexKZVx7CY9OGA20EkgENQutbJ1Ds68vt4zAPM9aYvXv+5DGUXsHe/jwilYWfx
DPcNTlKD6FgHBqHtteH0OquDsn3JGbjpKuscH6eVCpjm/RZMxtLdC1kwPzHfGqNlXXQt/jlS29zO
mer3Y7X1LOaUS/VPZZgGBsoFJtlkhJ+xdZagVf/B4ewtQ/8RppFu+eE4ajyeRR9tS6xGwLAV+ofU
twhC+mgvcQoIjAIgpEO1IUl1Ogc2MCzA2b80s4LA5QzhZe0iyMdoQz/NxF1V5Eb2gIORcvp6pg7L
PtIPi57dBU8ba1aY+kO6FBkZ/DD6qQ4b+0iwb38sEMeW/aMTLNZhtH0YRP8/4o2eYyjj5dpcA03/
WTTxwNCYt812p3LOPXaM7yy75SbwV9/2HnoxfwAeeiYTq3rJnZjFIqjx+usHV3MgSnOski4nHvL9
t3Ix3mTdvse3GJjX5NcZEpJ/MW9P4AAPOWDfQecRxsepmjqIXj2PoEIsmRNoTppNRr6fCSIk4Yfn
W85vERnaofCszh+S392sL85MGxSELVLBScEI+0aGEAAb2Yd1l6iyfBR8yoo3/0B/FiEAk0SopMu8
+oMnZ6ncQdQjYjzkxucK7jGOIgTf+QwGSD+W4/8ioxP4kYoqkH2bMnl9PH67aq3OZqAuEDbolO0n
IibW2PWe/tZme7V1GDNWJrLjIZwSSgCjFpYWu+7ThDP9wVKq++aVzejCJswh2Og2RfdIlVgKZCH5
1k19SzfVSUsmUjQ9F3ibpM5yKRwoub0GF59iuL0xKcr0bl6U8VTX6ICUV++3MuAELhdq+H+r1CZ1
ny2G0U5Xpy3AuLB/6lEcosofmJ0AUt7exFg/+uqbd+0ZR8+1O4E6j7X0teSYdLv60PpNT4Klcg48
OnRve6ivixo/oSM4DqFBn8OYIJ7aPqMbBjc/0VyRZdCeWe92z8JF0KI4XeZ8GjvJZ7nUHSFyA3H2
IT6LRZMPwd4NQxs+LlkkVzdaVYQZPmpt0JliAjCRJJp+zPfXojc8ew/7Kky0i/nOLp1wA0l/Rz0o
qVY7oUCH+cdybgSxqTD7DU5NFHGIktRhwmkQAW4f+ppmkKshCxotgFkybGxObV5XupVwtwI5kesJ
si4mcQGK7TwBzhuQe4VuOCqg0wXOi6/8etmZSMFo8YwEpqNCiRnt/ZLdJtUwh9VER5y+ver8LFoc
lgD47RzEWZgXAKypdQDfXQ6raQfttD71CUkhKJYi275XRHtV/qXdJHJjMlE/jE3AlAxztuBn+PcI
+3nxLpzlHb3U8erJvOvvDfZql30c+p3vyLT7XMUi844/3TkUOa38vRRJogdXsG1BoYjPqbkKqjxn
40C12OMNcHgGdG5SmmZYmtXaRz1ZL1DoyDOn5zqHkpYNQt8ECj60Hs6mHxC3YdeGbFutGEi92+ay
UIHJVZrOtpmQr1w5bmKExX7WLiLLnTiOBrhnZb2tXs8o8bZBUGp0RSUeO2A3AXRGLx5g58K/7xKJ
Z8Suyqmsisjm7HOwfbAUzm79qxm6Za8ziQsWyRlEG65Nb8T5xhkWKPlXI/CYuWenO5A9M9A9eWl9
IODXqBeQn2M+tcwYluCKvvIz2tzC1c3Xp0oeqchjhy3bmVjh9tAmwCTk/l876lZsO59kY5sS5mM8
iowa6ArNbrcKLPuYQ89Vi9wFeHFT4pExIXAZbG/+NEBcz1mOEoAJdBi5vtqXe5imgA/oUlg3heGT
YmFIEw2VWI3/KN7bn16OiEx8Y0PqYNDwkV2WuLuHezUtTjbaK7MLiTIKeUsUW/DTT9NpzgVZ3iKE
TEFb1hg9eBdvLOgyUIgpkkBPJYEttEg/AKjAmKsIn6QBOr3tCKoWoIkip84OGyUdZdyJsu8smJgV
Qbj3wPhis9YJw9DfufjtX/fxpp9DOnRt6xYcr7V97HiPtEUofZDVfbjD05N9ykdx0taPLAy9m8HL
MeGbvq4MtVG94BEgxHzGLdkWEXBvVMsOmmw36UR0255jui6SYm7HTGfecg3kUo907pvd+uqgm+Lm
ynlsYF4/fAtnbaSmJOJKnqJv7byHrEwrWyhhbQXyRdSrKo2I10S8KlygiuMGzi3TD2n3Z+u89/hK
Z6VN4ZdcCSnjl2qqYg4huECo6yCfYiFuPwFIuF8HqstrH9oddacEx50ugp1Q72uPOyKttv6/T+gV
NcDqq9gmYVIgG7fNk/cwPIO23vC3ySSFhMg68rxb0G7IAzsGW8PywqFpaReDmJ0uGMCnfL6xipWh
fOusmGIMxuvelsmb8PPmxO5aWAaikcdcZj8/+9SrCQhlNnrIN+/Q4WEfSNimVJu+nfdOrMiY1KMa
kwENL05Uz4Y9fkv6YlgtzM5IM3vafUADlNH4F+iMsJ+cB6m2xQF4NNxnk67+SSFk93CysywUfwIj
VPnvhmPZHA5OKNUR8K7F20oS387G5bowXf1zDSBu8JwbFa+3N7eVWjLXxPs+8owH5x/2ektsWqsn
BLodz9mfYl1nJ6TIRWVB1aBrja0kNffxEsf+BP5TtBRq+4r91lEDSP4jt1HdWIDutP9Wt1xMKAJU
PHDfm+yPNnelG94PPxuYoIeEt3A9nWjY4AUN74pcEW6C9zfLCq3Elt6r+3oEPuar2FGw/UIAq92x
BFdod8rYCdHT/TvGS9O8qW7ocOPVIuYcPwP0G/7NQv5GHkgm9F6mHmcZmIq/A8SnCNmg6KqBEV3p
Yhf0iUqz02OAXHI4LzFeRXLIdltdyviQkywFTmWejHAQgbVgKxjQeNAod+oZ5/SZefL2d3XI1OOW
9yJUnRAWA3/xMfet8JPnn2nRj9InPYXZXOgFBo6FHaxNKvPO5mxFwEJWLTC26IpDZ9Kk4WrbrjKs
cRzdbqTRlKtlyRgh8j5KGmmII/nHiuIbKnIpQRUnFvX9OcrP0dQ1ARg0L81bZUhfUBr3zVE0OBd+
H+FB0SonbVG2Rv8/I1zjDnYHyYFQHHEp3ScRAhtvPdXoEmajo/kankBu2pxWQtPEo9ZNs8qLtkn8
HJpvevEKs6yCncoX8ZZ275AO2L9g8RRXzIM/kxO/tqvnYRU30hkSJlGBNWOzQ0xkmEnHJhlXyfHL
6ancL8XILqQSFRq24mc8u5PFehfwltMG+5I9bkOAoaDuCt/jQgZwBWbNxhs0rqHPcsb8FhGcn0en
uMEJy+QwCOQXmH88pwpRNRmuydmaslzubI2FM7C1v7ui1nCHwMTxREYhq7S+jnGvPwNGME8n5bBi
iNitMyex9MOLj0kLL7aOTORwqe/kMMKuYUnmbpuRMDo5xwOahTqjB59+YVW2NHjQcfPWxFCtpn4f
EO+w/TowSO5EHWGyqAPwQbsxa5vVzlStoJIWAp5XwEAvIJTdkIpirsnWwrVSFIb/wl8KKU1ljewp
53UaGeV0vLBgDY5iD4oor7l+zDZ0pw1tdpcwdnvsoh31VnhswJHmcIvommtI7D2XTUvptOgInQIQ
P0QK15pVHIXttRdMKN6NEY6jySamu06Cy2o4pVjHJAQP2dWTmInzSKPUkNOogd7ltjKq4JN1wMLO
eWftuiCdigc2tBWx4C9Dk/zlhMcsJSe0SiwEiCCFhAQe7i/VnmM0Ykjff07R77aqqdeRTFlvS4PK
fxA2iR3ovcuZXvkE7WEuM3T2BTI7hCqRDrZkAWf93ZwsgkjRVJIYyHu1GOtzHaWWON/WoFZlI+GP
2XdHp6rsxgF9cZx7n39KGGPxG2SkTLY+LoN6KLQ1FGJIX9FSFm5MPda9gS3SI7tBOSKS/pC7AAD1
HXPjMtgFr5J6LcOhvRl7IWjowYl7tFSV/t0FdAQQc0eFFsGG5l7BfdIryuJ7VMkQuAZcJb9t1pKo
Xoz1mDp9aotD6h00o32vTQa7M/nqguveNrKyZCQecyBrSUFUJH4rEl9l10E3d+OzNOaCKbI70UGO
XHLBKQyuc0ZJJjY3T1hw/txPGE0zA0hCKP9yAbvrcInDEGFvAQYwPYvLcNqBG4OsQjuMsqmBie4T
4WnnPxj6zTH5iw9U2YTbGalIPPoVU+0t3mprfmUo+koQIbbDKiD6zlnrxJChsJeCAYyUCK6W/2fl
zirFs5ddYD6aEkPqbcbj8erxFTdADpAQ3sWYHglJUb5YOaqotAKnGPPby/P5vDX5uxmLm03SBksn
CcePZxB5piNkrctgMfH/KY+CzKn6G0FGW8nMcFmlpv/RC5v2R47s9owN9joNr0spOM/CXgO63yif
nXxU39iqeJzXKqqX9V96htmnamyIr/0zfN9gf0Sp6VR9c5G3IAYOKZnnEyI4TPWWDJDyErJiwfDd
fWymi73qd1M3sUWPFztVSmcq+zEUyNyk4ZPAWagjlaWH6kqU5tKfhTx6g6huvKpdJTiPSIUVbaUv
FRsqbJEmZygVsY9OHoHKzQ59WUC+d6vfxs4GdUiNGRiYvCHNhtd/1Z+Ydxw421DkJCILBlqhDsqy
Ljij9Q+03or+L+uKpmEZP3+U9dm3+/Jp0+krcar19yzv8PTJ8UdfxwTKOaauGtXSbnc6lxBtXcYo
QRLsOEjA13ngJWQfwomg2edk6ea6VhG3A3TAFqD1ChfbRe/Qn9em7PA2HxHtRMj1VwGr6CGg28nq
iZaewkfxpmdOhlITmkUohxESBRtYERVpU7Ij/3Al/bL98hFOxH5ZqZuI21tuNcElx2oOb0nMohD0
hmfW2884PA3Eor18EY8lTr9rF5AMMQVwvVzcum7HASAW5+JUjxKCxpf2N6EtaoGiwwuBdd0SdYiK
oWd+4xYZibSVuCiV6jm9g2wJ5hZuZsM31BepRK8/wUxsHr1GsU79Fmi9c4U4sZ0E3NsH0lLS6wu9
f3mJe9+HV/w75XIiYlSJzbn1fMboxgzkkF1Skity6fDwEe+hkkyBsRGBg1YZ4IVhr6ppuXaCLcAG
QbsGDrmsm4vCOEfkRZ0/8/HDPAk/NHLZc63YJKRw59VirYHJUDLDDz3ChwRN1KLYVloGwX8H72Dc
zPqYV1W87FbaucejJIeQaR/Yc8U1x4CR5Y2aaahKVX8gOEPO+gjy6h4c8Zd8pjNE16cnw7WSQUgt
PfW+hhal7+Jc/1vDdklI7i2CCjhYNH9bONkYSNkRArm3WjNPiTHa12NDQ7vhUonfufStfJn5GaUf
2tAkhPGWc9lFGLaGSc00f7EhTylNfpBiDmMWeTPowJNuYf/MF2YThJnTnVMFvxEUFSWcKb8m9YIP
LjlnEoYuomkxGDOXnplqkNoyKu51EowULfqEtr7bzuz2gs+mA6IEA0tajHeBNnWJtXghKZGZ86Y5
KgXPVtfa5JMsTp8/ga0iQ8o62/GyjPztrCkyR+xER4wLD0HvtBu2FZ2B4RJOVgNYFz58zRH/dt54
YqpJa+j9FMX05Ys6/RIREGNIoorIO3RszdhtONgaJ8pfcMhqGeTiWUjFwALIETBALzyJnWf8XOiW
aVNbHq9dJR4wP5TrfWsErEzXswpAjUOJ4020cdo7AgGoJWQmBoNHiBQIAFhMdOL8mlitaA226WWm
Ud/CICfHmEXHxCABFcFC1Ia+OxGmblWtZA29ae9t6xKOcoNHovaNMB+/gVpDEB/3zKzdvrRSavEa
p66mc6+22rkgkXet/3AhmgNiFmv3hgfB0oE27OoL4Y3VmpTCzxdDy30DtZ+RjOBbq5IFy8j+ppAx
lSgbA5KmfXbcEug49giQI6b9uBZd2VKbsTTH5q43aIIAh46JyNMFafiKSU+MxSVwb/6GKiB/3sqD
kfT4hF3IzfLgPCDeVy4+qMRNJemTg4ikpeMqZ9hc0I68/TTeGqdZlfyJuNNfnUUynJIDjRCdSXqM
Z1n3cq5+Fj73zKzwLKLu6t1xAqRbe3J6nK80KuC8J22KdkswL4PrBgPtBeN9u5lrnEPzBJjeb6NW
xS+Piz/1szjwGf/z+rTPDft/oVdIRAEFuk+8BC3myVwTRbDnczackK0vljk2bCGthV3cREtZIYwL
kVemOJYcmu2bgnEGqr1V32aH8bCdCYT0G156hpl8lYorxGR6Bal4i7Qe4BtmpHtpsY8IvreTrjAp
AFEfLyuqsuOm8XkZjmDqVGAgfrAT4sdFqJ76aIQayTA5GkgWmNNtjPQGteuM4u9q/BWJceX/Bcpx
7gUqf0r7nFY6/y6zhuwU6Uoxww0lxc+F7aTq4t4COP59SjbCYg7EAIpbj3J99aY/K5di0GywYR7F
oAx+0ebMDor/ySVPVWebO8mwGyopxnI23hMewx2JbYXaHGxoY+JFTvxKoLTEJJErnlbyJe6o2q8t
3Y9Y1+ujpMUHfCErFyy1qbqcZzOOlPVHTY7JhyesT1fbZ5DmNBp6usX80s/0hdOXMcVP/h65PO/t
KKad4H0LjOWcVJzESHmUHZjwBzV7vT8L/USolu1qwOakoBTBzl2irS3g5FFfenInRMf/5HKpLH5Z
0B0HAO+XGueIUs2GZ69JK5dfj2jY49xRk+ETn+ydiOpArQT0+uQeX9iZj5IU1Jp9u2UUx267egg3
7HwBUCZRWI9TVI6bZsYpfbcPml00xNoadA96mNlbz6+1IvsE73R8PGW3OI49lVnOAQ6KyU/EAYta
Zq03LFMeD9p7w4f/beeJdQqQMEUwk3sVHAIFZ+zKjavbEsW1C3SqmUlC+81QKPpB7Cc/px19YajY
IJwgbqwvyEJhStuTph1ZGl1u5zqITm85oJO1ZJllpJfFgT0mKc3Wls70Z66A5y9yP+3VRBlROapS
JGN4fGBgU5pR2bjNH+3LhW4ChL79vbd6tSc61O28ZrpWCHxp9DkvhEQZ/dgSf4FSjseXF/Ib280h
Bhzofpgv8hU731HzV5mnRl9oXZqhB4lByaKoD71lTC9v39Mj7AwDBwTQ0/dfkHUCwEidUsd5u+uc
E6MWoKjdOS5Z9ivu5K/lJA7660G/VNy+YYavW3SlBFvSxrILdyImnEwZPjfdAKaUw1/IKFDJNfha
sZziqFzAfbGS3jquoSl4eqBi0pKKGvp7YgpFzrCZJrAgeH4XegqgTxpw+WvA4+gRbVnKQJuMRnHr
K0tIyD3vmD5yLN+oQk2EYixvvUEyF22Uwjtm1dpzLo5AI9J7e8uWih1KKdcZEPjtbhhT9JAMIMH8
uqO+L7+775YE0kbDw48BcRteoX9EBht3OGanfAbIGiu8/DFDa4HeZxgI07D3A3Ok7H/2lPs8A0KK
fB5HPESxMVFdcCFFr1l4Srj6CXhcGvX/joXBK26yQPZPIjLpAcQ5tj0IVCBuBH7SIp1BIV+q5Ql5
KWFpw4AfFcxcKKkGtIM6HJFeulXv8ccRSnOX5Mm/N2Wk6wazqpqHnrbIfpE4SmNf1mJ9W0Hbxy3T
HGrxwYFB/oLED/2LXxh0KMQERRGO37jaFHFcPuZVKldtk00XRSDHOFXTdMb6Aj6fUL1ZhratAkLX
H55llzwcrgBO+TRS1lWFD3dqAK3vU8/fz6jnwRCOQidTs06s8DazAv35JnBvJHVtk4aNRM1s8PGi
XUULIhWfPOB8UB0BiRomRoa49gkxfuPVwPCfyE2AKbaZ/0RNnP8cwIPJ8IPwGDycJzkC1o0dTeJx
+3KW8vugWulRkTPy7Ri0IN6KbVW3dSWFxGlhmuJEubq9FgapuZASm5rsI+Xifn5SSyzccc/s4P3t
tzSNx/nLYiM5k6qVDCLx6t3bpNmuyKAUP7590q+WILgeX+E9uZFQcBO8aw0vGuX+sHQ+ri9btA1+
CbAJFX9gYsOiIjqRkaYKObys6nGdTZSeaVn9NEbwmChTTScXkx+22IPrIcVTf4nlee0tbbuMHAY2
zR1UvkARFENGYR2ilarfKKHQCV01WXYSxoud1cn2y3l78yVPwg6Mi3wzTlb7FWT+UeNxBgcVEyj1
7xVawPAeNUPwB8xPjqE5wtQhv1KRQ2WxLrOlIYJ9Bu74yjx62JGP5q2BjIsA5WOYw/xDsAK/NvBm
mQ7vFgzCuhb/t1a0xBhK5vGq2HpEvOu0abS6rKI0FIDtUvbtPbNlrC6YDBrrz02SZcKC5w3t7v3f
a0GD1rGuSQJ882ovX47uslTQoKL1ADl+R69xiMsBjjdcIMJo5ilGr0IooqiGkzLVHu3RaCFNdIXT
OBi97e6MUozMQE82GdpO+agtTJ+1snhU6Rxvs5o95nDRaKgGFL6ZCUk5rgoOuboV47KQSx8/DAxi
hiGbttYd0WlIz68fRobcBUQ6OWFqZ3ZSc0RtxTYUN9BMHv/YDcGHtk0iP9Vgwqm7zH5Qt9bwmj/c
Xe3t1MYcekchUqWWgQMnPJmp1re/R+RbE3mXwuMsjrtwEXZC2Igc4Zp/0HjTMzIN1HWDyMXOPuzO
Sn8nYnPsteQUUV1DHHu7ZxH8Uc5MvFUeWM31aTunhe5/VaBzp7MJaiYwVjMo7JylJ0i2XNILBgYn
YFR42C8cO0czCvFe+eYn+cNWvycJ9yYstsVftcRExdNckeQ3/+CbvkLM8SD403I/e0Xf/If1wt99
EKhQJZO5lRuSnDDb1u2W1/IDscUMmax23fTgqkVOed8QgCzT+e8i7LNy0k5FZgDlXaJLpO0xQ0fI
+ldnOrDmer9K9/fj/4USNdCFZxjZLvqTEcZvqz/IKb+Xd+iJyFXSAp6xnGd5uSlB5+Fa/QEuySYG
fuEv7uS4HEVMgnwRTMwkmqdvliIGUDf6Qkf0auJIk/BwmRBRRDLQ4lgD3ExnQSro63//num113kg
z3vOBfU/7fVx0krEh/4y1gmsAEj897YKMW2e8rp+CVNO/xWxjbUHpVgyPkul3ZPHSZxyQIFUIQJK
7UbUc02Bp+BaNfzgeMVDR1xORgQQctd2LPHwZfWrMdv5XsPKMRfIShHk28qYpqeKOjxvoZHRy85a
VEjxNfmRDbg4evVYmePlRueYY9Mt08+Ljm6I81fMXPm8rsAUK/b//K4SMtmLgUsqEv05dKI3dKlU
jplL7qeZJ0onVC3i+gLOQRbfRDESDJ8/znU1bR4Xr2ZAWK1BdxdZRkWCdeneRiwPSiXv+8+XZrP2
b7+ugKA/MVLYrPp29XC/KzuS1MJbH3oK8Hm08/d9pAo0Isw+ZFOvdhvnqh0EWICy8oDJBvGRoqiL
ZaduOawZnswyQCRquLywAeV5sRzEW/IOEp+OKTqPS+Cvx7A6egXdO33aJ7ROkln2q60ZUWaeuayC
xYnJ0EvWEgwaQa5ZBQFVRcOSCZYHRuU0ijscFZEk69ApHZHdw9vz7+2svf//uWnQpjfpXHF0qqbj
Bc/LdGxDsyXg9xM5M20fYTqBycoTLkDQQ6KYg51jcqT5cC3Y+5kmWMfaNjJ2pFr4DViKk2N4Ioe/
buzkx0H8THjlS1U66Mm8IkmeDvmSs6g5V0oY8KQXk6GjrX7jcj65LxTA0vdBdb0mqgWE104b6Jr0
Z7z/9dmDNIGR3nA5zmUrB++aCS1lt/q28KNVcEOPEOE/86UxXEf+YWRhee5iUO2fysJo4ZEZ7sk4
5JU38eCnXODmwrBNPQwu/v3ETk7x3SXJrENgmkxhyvBWTXE3b6TeNmlI3kRxn3k3jAYgcAVEKymN
WnRx93LPUSRRJs48SjLXsDJA8PZMiA5yaQHPJvcMATP/oIiCtULCQ/0iCJ/l85XLkdX+ev1BFktG
xERINDXNnTgLxRyoJ3483G3Oay8sNKTnkQiuFAokfkYt6pTeutDgnaBs21rVOByUZ61XLIv4eas4
adnjHbJWVv2MFpugg94AYc0kkw7bgIm3g7+aAyZNOvWC5RammtppBEybQXrf1Nhx8noKrBsXUTXz
P3jB/DuvTUdYBb+uQ/j10Rf85XPHCa9AUrzG6DsjSz6y0NNyafGsPYFykIN0b4Av5xXjLZxptrxH
Q+N+LMRPiyJYSaPhSqhbRYxbUDCh/9Lkvz+tSjqTMbOa76rTsJe7C/mfI1ALLj/Ut5DTtmb1OlLC
0oRgHpuIvHBRXYpZZw0N/94De4QUsVe0sg929v7K4eEAE2QWHncil+Vt05scurr7MG0lpRXn21JZ
0WiJGuxLLpcihDQXUmVRuXO0UMhVFaHoqKPAoWIeeCeVq2GWmX8mxySUWVoA77yDSnu8ZMSB6y3+
m5J3PdZpB7XheeX+jYRrzXB9Gd98KDrfdIACLu8x1e7YC9nGJQg/HDwbgdnGxEQKCqrrmbxBLrQe
kLR7siLMl5Ra0OUtod2rA174xj7U2ybfMNwha6iuKP4HQPhzP9O+1ikhYbwLH4cAG9yb9wAzgVV2
Ct8sAVGNc0+IKyG3srDlO3OMYtym/n73iD6MG2sVrbqzQZt3AXB9ZM9pV7vr50w5Nv9/A6QW3zBv
SgUtsjpNCdfAWg3wbQ5ztMXsPiDtowgnWkJwH035ksiQkHRW2CbTvtO9L3LtLzhuuOG5i1z227xJ
FZpiuDtNneeM/hqdo7TAKMsUDy3CKvuFM/M6erq4fjjEBebU2fsK93b9a5PGx5wLaBcMVWiwdttm
+8SKOqZhiPbaz9x8wTs3QDEDz90IhUHpRsXu9rvFS3yDnSIMKPAg/5zLNH0ULpaIBxOeitAyvhx7
PflTX2zNye0IAoQPDGFmHhxdyw2/hw6Z3ARYw6yw5nkwwJsxIfv0XaCZrLRe2nA146mT1tZU4aUh
ZcE+yW3BQY3dVBqyeLLRy2bhg1W2cw4ebpgIpMYXWOpepzzScxqjiqQ8XAem3Bp3u66wnFVEvokq
zHBB413G96xJCQBKu7BBrIgoVgiDaXG0FznBI4vohBMN3U+PTiL+6M6o8NXOjiU6DWMqAjjdErZh
MJfFCx5xAzqoaOTh1pajiYRXY5aujesrx6zjtDAiwA+kJUVIhSF7rfKwrkDR731X8z0SdPcrIQoz
xZHAkPkSoMdUQJpPGboMQfdJLMUAx/IORoltT32LoRJ3IoM4gX37/XsLGGjPjAOucL1xoDE1cXvy
TbwRkmKWhM69VDOsm5ihdYL/QrDoEIf7XQ/xGvKgXWET22Mn0eV+TXByvfquu3RZHmUKflMLM5Ab
MW7Lbgo2Dx8LV4gweCTMTGu6JuoZkJnNZT/iLrwTOZeE+Vx62UAiGyiO/eh2lCNyET3KzTWmGMF/
GEJsDzMeFsG/7+0Fwq3xgffUVgqm07OFKi+qqTVo0iImnqcS47PGHh25YZjRDOqb8BbSe6e97IvI
Mhm2oaEu9puN4uJAZVOWmWsC4csraQvs158h0xW+7qWUNt/WA9HBx/Pdev3lk9frnu/0gMw5lwSa
JjSvu+PcKmgAWAS5ItqzcTGxM02J03ES092GuVdpX+ibw2OMFDMH/cH5HuCN/zEIzLQZreaBdn0w
heJvqniqJKXK37vy9VIyG+RKF+z9iZDnKu6M3OPtBY4hiYAE0AXdY6XXTKlKWO9HGyBNFhKUYWQe
E5lUG8sn5H4DdWcj2YbSmP7ebWz4209uaqgouFJNGcEHbS+dEM/yhzzrgOZ8/eLSgu4k80NwAt3m
v7vpRUWmagZ4D6ucFJkgjoo+jJV7pD9CTn4/wjhNUYMa5hxB20u9ZFtXV0N5/IZUWnrdW1K8ZtsD
Q3kQoDwvFo53gwAYAWTXleACyVGuUu54qEbHplIWHMwILA83FJiGHDYbC6jf53KorFOVmsO8nkVm
F3R1Cev1k00m6/Ft3upg/tf9lyT/3jfUoCOVgAmjqoH61XD5OwCOlVdg5Jfx5PXtJmdcgfqwWORp
puczOgClFY98ia40T/67yyyhYZFwH34PrlXwqIavriZILpNGLxGISdMIGIFsN2zYZbzc9ZKopqh9
E93aXlRPctyGyQ5sLjrXwIkucSWrTl49P4M9rvkklrjdgzBC6CVlmxURbKiXlONj6KtWibXp8Qqq
ttNK15+gPzlX1riLRmLrQd4JEJDsZmh2Yq87rGnMvUTB+6Nf3HALVKbevtLsJccV//LnkHzTUhIk
Cy5WF29frZajseULQgraccAQrz+NtfJWvUl0Ut4X3tsSX+IiJaU/0chB+ZTzjXXjoIPezVgT43S4
oHn350oyqO61Xinrcb5aQYthL3rxZhuv/h+JcsihxDkUmhGDNYXv/Mie68qa4kKMjHJt4VcPBV7Q
zVhcP1ofx1HontNiC8UT0ZTkjt4iSwjSEYT87N1z+lH0f7dIfk2ZiOm3OllmOFcoBTokW2i9lHWi
WwWak77a1npYAlaIATglnQ/BBOsX30b/WCxaAayljpq5mvxI/eiuXkdI5qGkmxpCFKs9EGMmC9Ro
IXMjltVVgOH7DmRrBpH+abhqu1lb/6kEaftCLKk+sXZXkKM8snOuISMB5ZBT392MWjMOXRcQ1+jV
ib9PDIvCHz9HpGD2pACc5FCrCCops+7EFevpkXLI3y9eRGBMJxvo7H1w854hAKoehec5xT9TYXlH
AoCXFtpliHypH3e897kEzpbQSZbHhObVgnTxNBJfMabUUHgsv17+6mHecz2f/erHYHhJcCPeBzms
4EvpZlUPyffIuDMxm8GS7WOBTOW9JcCwHLRN6FLGME2B0XbkQ6j1nwG4U3qdToX6hDjoiWdAkVGm
EO6pcJ7m3igwDvN2E1SfixuoA6PmUHLG02ZIYcteSij3xOciDfDKCkg7fH42qAyJ7vbLr7dsX2j7
tSZslcI76t8jihFgsgG4p+Pe6HuofzAnjU5qujsIaWvrc4/2452EJOnL94GCHZUUW1AktYW0/6hY
phnmoFPwPTBVEp+xvrHsy7KJABq0QQ93kGylJpYtskGATR3Ruk2zrrOp54+dIdks/BzEuKvlfiw8
W+YqA50ixFqqCisSJX+gNUd2OWc6KEDUExsz6aDVIJRhUJIelZOn8CuNA41tuijPAMpQQUqVRPrx
VUCDXEDneEeiD1GxRwMxjdiX2QwXpqHlu+IEy3xXuJgTRZjeOViCstVP1oZ27n5wWJL9T6xVCRlk
GUwWej186zsYn9wUYcxTKta2OqFHMCHPt/d5N7QQdSs3CfjK51IywEq5p1cg3QAbufvPzilkDQcT
nyLkca0Ln1jb4a+65l8FXmHMTj5u9k8yLvQA3q/fB9MJ3RiwfAN+PxaXCD9zvsRDZE/4VWRk9BHh
JihWPOKP9fZdT7a9vwAQ2UhzHKeEqdbnvkjRtpz50MykzWeClwRUI6CPD07euwhl8Z+ELYobkPDj
Bd5spy3iGi5K7BD007AcdskRJslQS8X5zRXrnnQ+0z8s1sjHOEGGLxl/vTrdOSnvqZOWpmNAUaO+
4+2wgMlEkoSJL36/Xw7qlxe2jAkr5DXsqwPl4NmVJxKE0V39JWJnSbyx0hY6uWtzwPdCCRxCsbdX
uz3o9YI02o3aONzViirgwwVVztKJ9HhGpkeHX2BuGDWIh51GQ9C2HXMF50VZdTxPUw2sFC17PCST
FrlVNbqh0+W+sgw7qCHW4eLtpGJrU7up6Jz/kd7VNiHQW1DVGgufsXHPO3tcKiyl/CK1em7Jop2J
JBbhJI0SyjP8/Le512KDlxJU46Lt49XOGm8LdAsg8r/qQZXxtediQWHGNbxuVFt6pfhuIbasP2Jt
aT84mThzSUQw+9Och32ePS+Uo5R8n5k3LXps9HOqnmhtUIw8MeCMLJdRZeCVcyJsgt6X81S+SbZS
RMdvHuCB50mO68c7gewWN7oxAZPCe531x0Thm7/0gjTrotSkIatMugWmwz0gC7kXG/R4J5p51GSU
ILMd6s9iGQFswnmlAHtAvWvrW2WPwk9oRyPr6RZHm2P519TmSpNYk3injNQeiAteZqWl14LdmwYe
uFtovY0HfMJQw4K2PpqVjDX65+ZenW+Rw/+DPT4RXrXTzpxggnq77rEeWdxLSc08vJ47LOYR0pf4
YE1G94JiE+BbzX6BI9b6uRu3CxUhQA8XHpMu2g48z4nXfO5X/rYkNYxRgF91PZlBGLIlTYuJh+d4
rbSGeD/gIDSVciwrXuqm92bZSSUxRB4SL3mfokcE8M+7plqw93Ujn6bFnPzICzHamsGdjYXvyVWq
TpnyMfQ6bIHlL9Sf6DKwFpBYNWsAB/H/ImhdDbTujDV57zWz8E+DraGRtwH5pXOrkoRk2l5XFSSN
oLGcw5uHoLH3+onMjpbfGMe2q0wBC2ysusNJyMERTHxiWqgrD7GuQNq9mEa2WH2RO5VymnE+utAk
QzEuZ/6M4kmfug4Cs7w5E6c/Db0uwyvwrn9Pot9ei+zJOY+bRShFG6Pr9HaLPn4grf9d359GGSni
oO0VAnrin5K5C3OxJi7eXqiYhIpGmqACCrOwSr/OhJuBWwIWlRhNzibkS1AXZpSfFlWvfjKrccyr
eN05fAuj0VuIjqZr6m2NutuNOb+lB3t4wTtz0wgS9BT+YKNaiCttCjF5UzGURuNbBtMB/XDidmpV
fJ0kfrmaPWym9Df0T9mWPFOBACCch1soKxNpc4gglyqfet22CnZJ7/50BZVSb8hRmS971R0rF1BD
VbLHz8t1Koy6KyrzqSuk+90/QOCUTDgmDyYu114Pp3AAxtVBccLBpVsyAKgLaCSZ2COswylGnwmk
o5a7VCogd2taoLNMAPsuqWaluMi2KFgRCbkZTaARwxz5LqCWBGgtFVkKFKdL7cBCVCX6cGCB/u6c
yW9KPV9BrszQfq4DV0wVMDFxWOcHHUVP77FCyLrUg6ck34UyJPyxCeinyQBNCKl2omVzkolWLzDJ
1zsl349zfwoaj2ufGzTH/P05COMAPo9VN4jeWTgjLTqL8hDLn3njiGuxu9D7Ekd1DRA4jWUo4bSN
zh3HAdMGCrym/o9sZuYRyJyIBPAGpUbciG0XHCXW72aM3hcWQ60Urhmb9uuHQ9Zgm5h2YtWcx8Ll
jQ5onp4qSTP0j4eoTzixH6ouajVavnAmhwEIhFxKeIX3ZV9Bo8Ih9r+aVctk+okV+ej0DvNz78ku
0gXmi5yzo1cUVyajBIJqlSQwDe3RIYKFhpMCYtXZnzl69BISsBlBAyZPTRpnk/O6Oi/rj6LkbiJz
wOUYxYarZjEUgKbJ7m4/Rc3YEQjRsWB8kJ3OUmDjYPgCb2nEPdOgnVlNGwihLUhsY74UpPb05J2w
ldMm9oXadCOJmUsXt4vci8Kd1g3pwl8X+Aj01pMhJVLkKKcMi4eJhzROYe0PBc6yDSJ4a3GFSg97
BLMw2gY7txYhHHnJVjAtAFhqn6EJWkPniEdVgBpDCVI7Du2UjGIXkd9D8AyX/hcID4oz6SPhN68b
2PhClq8YO1Tzz8neDupUX3Igb5WUmGHPObld78OHphxUUEr2MVSnUSPyP4XgvT5jnS4xR0ljTm9b
t2RattW60Das56UCb5EYxo3gikorG9tdSk8pDSJK2+pFAjRugGT+mzIG9RLxMipYeHIFxONpjI3A
v7iKzy/N5QqhMwCfcEbqyHTAj5956jYQZ9To2nVL4/6nVs6raKKFu9B8wYD/c6VGKdftL6n8W57D
Qvv2KNvArxp7TQ+OjAuVohTIgGk3q/JbwQNR1KdryywfPDU6sncWp6oiqR4O7GtbU3k3y0/sRya0
BL6lvK38QfENQ5Ip7cx7gjxevDuVMiO77GMD0L2cw+TkzF0CSl2wzcXk6EKeXLjYHB5yn7KbSaHR
6VPlrqPUre6sR/iLB24De3/fsqJVE43ROmmDgDF5/ocjGW7ffayqQUnf2yErbGyfS/vXPI/O3zkt
ZKfmn0zcD0Y/SR+IaJhmvMRjc/RvDhVBKMVhA7YdmvwrnsXMWkA1z/1qLaDAiXLetedtvPqE2kz2
wRnt28xdYmvrPsfpAp++5O0JeIJSKX0m2wtwxTmsIU6GlwekF7JEhiqKJ1TgbMSChgpBjY9FDJog
5iy2okzzJGhNMqgspZ/DC9G3lnCxF3GaFBV8NVyul9UXhBIH/5DHTwVKEd5E1kP+AobB5mPDo1uR
RkV12m80yPozadXr/ffj797YulX05aBuDUXvJal+Uz0mUWw9JrE3/6TExAZIsDFrP6JeX7rrNuLa
WlV/6CCvK0CQOeyk/glu/EEz/4bqhvpTtrdGJatvdg3pJL3500hMFlvljWHlcWA4PaWvdDqH/OD8
bCpBY8P9GuGNg3zd9yxNmImNFbrAzsUz6GUo+5fpS05wmT4KcX0CFe423YuiGDJ1U3TPPSsHQn3Q
pfOPmrAS0jBtCE8Y9Y2sXrpylsQNi85OZO1juNuxtz70t1PqlEPlv/7LLAlZ+65mSkP/b92ZK9e9
CzUEl3gKiAdIe4BlfsdBpxZ4XaKS4yhDJvtIZqgCjf9sbktnxJWigie4oue94PDgDs3ao28FLYts
fHwxlflRR/1d0bOr2l9Ev0oUG1fsBMl6H0acFQgqhSPlCCVvXa53VRyyKdG4QhzOPtwqWJl0V8Ew
jo3P0wdPAhoH2yEUEvUC9Vgk62cFHup62oNPAXbIjoCzocPXCsh4prdKhjqHoEUDQThvWxE7Oimk
p2RAJi2Gm87aioSQyIT9kLu7CmWr48y/jnhza8tRKY8tI5AR/xwidpud0mZM8xn5ePQ+BmDDL/0o
jU45j+Dz6jt/7k5plx+WMiu7Ix2cPV+qsClohUm6S589Pe2gUpCfGDCEmO7ujdoTkakvoKG/3jhB
0zGpo6HU69Q7uaK6PlWqn79vlhZnwV3tr7GzbAP5NDILMWjXt6PRUS0FiZGUImshlkUZckHlp2Om
xY9r84RKP5ySEugyIuEgn8/goJ3hfUOhp6cyxBQtO8U/Q7QDewHhHrWzEnH9p5Nfx9jaTDlz1Aym
DnHEQxy1vChYe1j0mYiCoMxfYBk9pmd0LVh5m1ISYG9GzkAOkZQGkeElYBykJqOR0RchzT3gO0+H
YZkVf1infVztYGglzpyTJvbV2wWKXfCzo/3P7sGKIYt9bTtDeVXVgMgDSewYyp+Dg6uFf0NffjmU
jijO4ZIBeDIv4AJ9jQZ9v9ypdezY4G+l9RHNdPoFZqABTuLTkv3pxrsaOWhtZG2G6fNu00UL5H5Z
ZL8haWLSsrn5nxhwxIcUp77vkqiTVUyrhfZNb8Vj8axb1+qOSgpCM3Y0G2Iat3S+4EAPeuLNhNWC
G3CNFmGtGBMIXzSfE5HTI+axALrAM7l1A8mfsV0ygN/nSsn+p3Ew+yJ280X43ncS/ZM9bQAu9jEk
gc+IfwmlLaDYq8nUmt9pgszEll3eKEcj78LHTFu9VV0DIoODmX7wlytqzWBm7MyHp4NzhItVFOZp
i0QeKpZ9ndR0FLHAOXJNcs9/mThB/+mXXWxR+PlTRzut2HysTMMfyaIg4AJ9ZbTURjkKd43Td5L1
fw1bGjyWWkhlFOPbHT7xbsfs/WG3noJ/OBNifQiIqpsSBW8+w3R05vQzVd6LBn5pPPRQ+ov192+0
VasEvkNsj5HZp+IQmnZmkp/gFFttxaoibG+DgHFwYo+oxW48/bC+94UguKLF5i2JoVZbindcZ6F1
ej0Cu07cKzV6wXMPFmGIB28tR7SbcsvHyk14ifwa/I5XXe+e3l1RLp9QLkR77wSI7HJNgyQNBmuz
MI+GYwxGkI0MImH+t9fSji+Y7GvG6RihK8XUvRUv/o4FNi7lAu7UCAHIUuW+Kzclicogqs20qE/J
3/4lfEdcO1KhmMjBU1L0kk8zbjYoFJK7xz6fTCcaJdi0mV3rS2Wl/G0wMA3lgHVWLSHx5YK3gFkz
su9E3J3EB68XIpaCKc3gvQmNyshlHPTWoD8jGDtxSwLNmnE9dP1Wi+bqrVHL2lE//ggx8l7VfGKs
EaXu5jsdJzQ7dkdsmPMblObKb0VCZXOMYZXgRCsx3xZSqqQtIFAYmPtlnUtQ9DvL1CQF/HO7TFM2
5Ew82zbIcgBsvceOBV2BRbEQlTIuVKUFbGAMIi5Bx7joyxky2WzGCknwE2svur+tdmQRtZgRt6V9
ytxLg6G8GWxzn6H9yeynkpJJPtD8f35WJ6jcifQKMijJbZhbJgSVI11tOzgq3pr7tQ0LDv14mEMm
3tEIHR1q51EIEM5x2G38LC5XMeSxQZxRwlf/1z6zFw0b2m8ltCYpLzA4pVpcGlkkhdYm0sqykCqU
2Brny4jbp67BZgRwLjGCPkRmRoszp4M96WihgfeHRWuw5E+X4Z12eLuz3SfQjbar8cTEi7fW64y/
U23C1gQkFeJymOagrVqG2tOIXSoeYYkq/nceHBC0UswIexAUoVsL0zOIfztXlPMbUHffASfu4LLH
YZ9djjtyz02CbUlPSSZX25aaR9H7CQ3TSAOto4WyA53+X8KLtjp7eacitXIoHfnMqqhqAsB5KHJ+
OX4rmNadfbCn8xFIDF6k42cThkzXh6HlMBRiaVMW9goPCQ6Kk7pC+j233t3TnmHZX5Ay99n+iFJb
g31C5EcR0e1Bh6wwDp5d4ZqoY1NlEcw+a0EOG9HvWkuRElyRhjB34TxAMw0jbT4rco1dP9P+rgdp
PERAsgDx/YYtI5TDBBEP2TD4LEAm+I3XNt0kpZRYwtgSGQuhE4VJZdU/DX7TRCiBXCU6uAeBUdk7
UtVFomWdU5AP7iaBz1e39Z6IIIv9V3qRXMSJeDogCoKOEZPUU8sGLNfyNtH3riLFvw/X+r1K/K43
Ap2+A26dgj2vQVw+Yj6lZDWqo6DPf1iAkaBOPRyhZmFhsdE5BD1E2pM9yI8NJHTg1ySEXBrVWNSp
UUnvC1goerHDv+jzQVP5Zz+4JaenRkvwY9OPLJx4t50lBruIYGgQYnrTh8JU+eISiexDTH3TI5Bq
OkTB6o1U3VulYzhChu5ayDhDVrnRKEsApQ7F4dPgnu0jSa29X5FgBFGnqghcSbEaHin0GS3pxqvc
jFhaRSVRQuD9Ml/FKAOgK8wTNoss1NGxzEBf5S+C9Pl2L+7tt2Nrl5BvSi3gq4nvT6K65bOsAU50
PQjWVzJci5V93YFP0XYuXN/89cz3JcGIJNhpHuURUdWObQCIB4LIiuNZpAurlBwQG+JuBYQjVOoC
wnml1iyXnQxN/1XDXgJyEaoF8xBVW62lwBQ4qrWOYfMlSkHgcrqJqO5TFld96VC7Y4m+NYngiMHd
AAQb725wS78jN4puJgIPoFv2JNIeJr2OqqzWFLppCMcMy/TL78OMHIxH7qwiv4POPe+XWnAMRdCH
zg/NOXcxlSUWqJQvyZVDBy5ummIKz786nFpV26tUw5AgYSCy90aDKfIXQTybRIpUtDNxe8ENkhk1
1qjr3ILZpG25n3uWe0N90V1oDrw3LubAA8mljEmaGVIXSd/TiPsf4nTjKMseF5v56PKZvgDj8Cu/
gzHRWO21wIOgX4xb64+ae4ja1wWGTHDHqg01a79Vorr6Vlqyw9hGzxe5K2YcV3y57j12oIrL5ICk
Ybp2Jvs1NRSjLS/4QSzuPu/T3RGtz1I7PhCQ0rrgeLjifDO9ayd2ZfG3CEC9mOhddj+bbMoQtLaY
TcQhv4VEVn9ufOvxCIBl5G356YkwJ23mcwm2YXgfojJLq+1oAeA3//DNBwv62ypYipiYCSUjRnQd
RcGCFl69GgSux6WzlhHv8lnDgp5grbdpmLdfv1JSY400Jbi3zVocfl4VWIKKNOr4K2K07A2B1KxJ
Ek7JaRjAga+1lpfWvJx0xxp+RFN+45AfDnfoJ1HF7wHJnxci7eGKJzFPev5Hiduee0Q10luDnAF6
xFZrlBOs/ywHRNYWbeKMtKlFv4pv5oH/XfnPuONJ3tnYXiGgU3ypx/GqTPQKkmwTSTuV80EE6c1k
0XJI/HnDsA0OQQeBR2xwcb+mXsMjsOj4n6DExEzrnmhQNptFlhZZs61Q2okblb+8y2NHO26+QBpc
4M5hMCHeu9+74IzvyL38u0EWL9iC355EWD7zoTX68gN2/FT8fWLgt5x7UhkJzp2J7ZzyRzAJcgtm
Uf1E5FCNOG2Ta26syoyspXFuInzyZLwTpVnYu/f/FHP2LPAkVvyMaN6znhd4d2VKZt6Qe4mhsDHJ
NrUlX3jCQg+wHDZaMYVhS9WYADDP+7GzDaIR3NHwXUzoFc9ZMg/G0UwN1IoZrLExHsbZrSZhTPDa
sZJDGQywWqAM/P0cVg1lMenqrRcAILtH33cmwQwypM1DQfhGtsZeHtcRs3Fe48aIa3LQn9xzvT46
t57DojW1er20j0WuT0vAej1lpQcXj6KO0hcQRpoDzL1XuIuFAEnQbzucVhH+cfgaPVLvFSL6A2me
27S6xj6/50aVzYVX4YeDK4zfKZgV8HeGPqmBuX8FqC2aaTwXmP54ysoCFWlVeNH1kJ6K+KSVYr1D
lE78Hiaclmno8jdQegEXJEKxYaWZg4FtODOe2GlJ80shLC4THEvUmzPwZL7pm50Mtbv0C87SWPh/
dmKh/76Hmylk+8+dmME64+uP3aGt4Dtmv/Jxh9CYyRy4Z95TrQhnbn9ipsHDvc6yi84ViiSV/kuG
3hR/w4MeLR+eO77M8shGd4Hd7/BMFk7zt6KKKRetWZJjEJcSxxMhm9Y0zEicZ3lR1meBz2jZiK81
EXNOIlzgSCu6GYdJMVtHzmqNhb3bj+qXr9AdZx71/iBnxsthS28AfELyX+yHjuC2A16UonRgM2JM
i/6h46Zi6QpS2iiSsop9TF22TwzjYnX+PP9yw+djhm4MYloyq1fMHqVW3oleqE52KXI79xNtPcHJ
bx6Ep6KteSxerO0oWmo46BlSud2SeYbZ1Af4GGScpRfQrropjssmlb/lLSnSgkB2i3/7afCl5el7
0dMheux4lj/cyNbKp45e6ZWODqs+PF/J01SXyKcFy3hXNQ1f5mKHGHzE9A4wt6XR2OLjfcY1NdvI
/zVMIgdQxMUdufRS1Wu7lg2CxA2BWgSXzeq3d1G6SMZ/fYM1gOSzy0AUhxYn/gTCMz16o2wGkeMv
0VfBkgx3nVEYu0sYaGoJLFLMCyXKDVSgVopNatvSs9umQoJoAQxpcy6uEf/ifgpjwo0dr/pTGRnA
1nFBEJyccqrt4hX6ejVWUxZS/VnrCCRFUtnLiEAwUCqGKdQNfyNhhASxqeTOG3tUlwsgwMA/ytPl
s10/Y8DL0S4+PnI85mKy9McnrpX2BIGXJkY5WVZ5zjIo7xtx80s/oeUUCwxDrh2harvoJ+WMclUP
zZfTfkhPge3W+MIHp07YhmGZn43U+gthlCWiS9GrqSupJt6cuOJDxIU2/YtniyyQnecWWU8lKNdB
C00og2lwlqCyPIb7RR5dmxAbgvw1lxPD3GkqSPDNjNIWmNdD6p9D3mKs46kat+/XwHPiFn4s8zq1
hIc/493tinZZcUQ7rzaFOGIURuhYgmaLm+22Ekj6Lm+wZL3diuTbE13Q5Ce5ldpsM3tBFOwUPzL2
EpTFNvgkpiqilCrivp4iJkKc1lYXTQ8dzpwVd0g4loOABYTZ4iZlFk72jolvaItO7zU4/Ias1OIv
G+bMKAHILjurq1m/6IIFrwE1m42rGKrG/xHOAKVb2nWLFfOcpOybyLRN//twCspAAox0A/sGz+iu
gPqpBAMN3noxqL/lksgAERreu7n3okj+2Dw58M1QLW5HSNLMw5FLMRKuDkVrHWKlDAkkaabP3X8+
sv39cNgRb2w/Dl2hn0MGCTqHImHJSKyecxYFSNrfAEuhrJqF4TAuANfZYRC+SCZunuj0bHiHEhJy
COoGC5Kwx2BN/peSRStWg9BInFJgECczUw/PVChlEiCV/yH+jJA+n34rTbrTlUlP7I+77kWMahuF
ixjjwMBigKk62CXdvCB4RZ4T/RZIOtLRB7wlNlqFf19vI09o0MZqyaI0Vevx4EFPyVS3rQvbZ/8s
wEh3tXqDv5RNQ3qpH6bNtiGRcCQYP+Q9995ZatxMmGKET1AEv3R7Rgx9tt9gPpSvuwLqWWLKoM56
zCkkKOkp7Vi0CTvNBp6ncmEw8MzgTjlxtgFwoxbY+aZoZTJzjqwWJC/YBMyL20Jg95Bgfor/le/n
NcmAX7Ve5VOExjSW/UvexQJC4ebjuvfigE4dz8450iBD5f3fV0zdJdHMplfvv4uYRbqPwjQLNKLU
1UlKENRuEtiFay6KG1qi9AjDhytO5lPvbhSLPo3ghmmsveUTCnRrlYarOVWiDYdbEYL+nX9tgefj
HQgDPiJE1j/pZFEr2nOOfzoEVxE7C8bZhq0uIptgAEHHu2S6BJga6KCVJduMW9/Q+F6+UFEPBSXk
4onJs81UeVzPUUGc/hUjkDl7RiKPVripCYvaOkEahWXGdvCu1lv9HbC2W9UQRoBV1gqzs4Xk+TUw
fYi0+Bcpuks78ha6FW0GJOYsD54yinUC+j46o9vJev4OItK2us6ag3+hfe40tEwVSzP/MgQKaxFt
Xab+FzWpIOnOyvkNiUPL/h3re6/SgfYw8LANgDs+DJxQu3+EbFy50+yoFwrISOUlFKEZBmyF9f1K
jeLQ+R8OlLojbXHPFAs4H4k0AHC50c57PbwfzBTXRXf3OGZJEYdK98DmrXH6utdkoApIOxQyzkRa
kiLu/n/RO1jD+KBdo8SxqXrpffC64ZsU7jFDhWpBqjTR4yl9xC4WI1UzuokktVT+mDIAQZTArgwb
UF1AwokZW1ht3bu+BIZHA0uYsmf5EH1NIZj1QiGYbY1B7+mAvADA42oQTTzPtzuzlGuuGF8yubcg
FyVO8PqBCjkdUpQfVfJDMfz8pn2/PwqL963n2gAvWdBLhrEFpovhHYiQmhNJ7F7G/rXwtYX1brFm
ImqHbtcX4/Era5OabUpFlk6bF4vbrPf0prDnw9pXIIXAhg5fpweUtjRnWUpz94TAaVvIiLYVV8vb
hnBudK/1WPK01PCoK7POw1G1QS9WR+C/Nb6XHHMSNm6DiRyqUbX21j8j7fuV9tMrSqmKGXlMwMUl
SH6EOiLagMDaUzD1yrPxwMGVDhchrsVDcJwvMYpetYRG+4VzIyWgqb3Yp4q27VTjtVFnA5zpbMWn
8ihQzePfcitGuIYWOEun5JiMdCm4kXptA2OJX3WbGfjkuD/zpEXOtGonF8wrrG+0v9pterZC2tXZ
Qt6CN/fk29lBJiA81r2nzvueuoTiyxnRCQDPgDdY5t0tMGe06CbhAQmav3P2LXH38mShxwPhd147
IuvsGPOBFeSE7XBNQdGi+a1/jmByLmVPBYqeZKOim2NzdoaeVcxnlSL0SP97fO4U6a0F7+/FBvpv
Np86Wjzrcf5ZevvtRea84evTIFmCJJUcJm/G96SLFf3lPnI6iH5qQbeIU7wsqaKN3fv5k2U9bUMf
pcvEMlVxMOQ1sPXGKE3gcus1NXZUnvsD0ubKyjqMzQ6wdXMcsaoV2XnMn2iQqZ72GcmFJLBOtUw+
g/bpFRyB6PFZFDo7Eaz2JAfGjI/rj/l9QvGeZQDw299DMdzAECeiI/Y0mZyqNDR07NLGE0U1rGXH
kiVFTrm8ZpTLPPE5xLuJEIa1YWCv3LKRl+IPxPxskN/Nxq2rKwMmOJdSGO4w/FzI19O5AbGLaaJ1
Rc6+dCe398PHx9Df1OD6TxUhwuscwQn9xO2VUpT4tpB7xoSJM5IJCBEj+gUK9gnFgKrbKwSdO5ld
lf+csn4oF6Hdp1x1yCBO1T0+ZsHiB+/k64eJ/Qg37P7o/0yW9EWNs5qf1E59iNGJkZgvavvExxuD
jZbMl1aAK1dkz61eDTeHPlEf96PG3SwTigVmlHzmi0hvZ7smDhIKU9mRgd7YS61bsK2WbUg3L6nA
cE1dvrNG/OlspFHi/LBLeadNbmHka41zVd5yoXmUObOxFPNrED80JCefwf5rjQ8K4OJSys0yb404
x+eLejAEkBxH2SItjnByXZItRpDqP6J3MwFy5FdmfT2W1xgiwY1E46H8pa1YgWLQVWPEW1c22biO
9V4Jqih5ElMQm1tG0thxIBUTm25/Axe8sPOt+YLUtYQpnbuVpk6gIxYS80Bq8T5rbH+zR2VzPq/X
zVkVyxzFdAy+PdZo3Hu8u5Kl3YQfLTtw+TqrCi6To/TF+eLdQeqLzmrqNjy/sYCdjRXH0w0voKR8
6TvXAhcgCsOq65bW5ZhAQ9tshqKin/xSSIiGEtf4MDmTKzbw0IUrldKlZdxnmjHC1V4DjNaSk+VK
dLzakmD08kOs6GzxXpBGI+hpOO4G1LaBtuCBg2VkzCWWvkV2M9lq3C3qBr9iqBxGSFg4swrXRPJl
Cgkd6VqbziaDqiATuhc87uv8xBS4BeX9MyivYX/qXha5WUxFc+Zl2iMRa9CcK9e2bwozf8NFcHmJ
TusZEsBQ6L7vNMaykzGEx495+r8GQ2ZLgGMgTtSrHWXiwMR0UjX5Id3T21tptkTDQVNED0ZiASdD
Pm2cO1rrX2oo17q41bQQ5RHrEIuRn5zynv/4YWkufONSRLZ1rS8+7mBBcO01sH0rEM8XhiJ1hWuB
EIpStR8usLK9TfgChLdvy6TyT5p0WBt/jb1M6uq1JiYyKNlD0uu19FYjzL5u7tBABig96wddxwxj
d78inwdegiwGYPxI+r8qx7Seu3nP8GTlXQmdgAPoaT3QzXl8nZhKcSmnVpV0FZ83Zqu08hAOd/oQ
iPiWDQhluBd/6QJn2Btn7TvK1/hzgTR+yq5PmUnJcmiRnMFscbjDlBjftfBLIsPUpU9qsyHhxG6/
3baqQgRQDMmjG427eTosw383gMrgRUtD1bfYpZ0+akxxEgBwpZOXoBWjT5mL25mSPCPOYVZs5M3A
/8JWbHSEvMesKimO6tAq6YhDyYMI2dpjyCNNm2kNgHS//H+YUwvMZKpyWX9yGwhfMM5Jmn+nNH02
DuParsRsr+X1I5IzWgOfdYfilMLJr/6U4rb66D3FRCS+a6LikZa0XH4EKER1IToGng9MGXFwI2Td
ov1NV9J5gfysmN+d4JsRqej0PpwneSYtAI2HId4H4n15Auph+6r4vOUSROPMwj+sXMBA65VGvELE
aA5PFxYtQNOATifb8dxNkMo3pDD2PvH2T//PDOFR55WXqt1MGklopDy7pA3qNHk0TsplMFZ75o1M
68xfaGun1eKWIwPxbvSeXyO7P5RV5y5bGPGE8dhOacUmmb6n5XBnYl3GEFR+9+9GECXZdXFiL7SX
A/dcyJdzTqnAfED+Zge3JaLEI55TzV1Gij7vSIl6Gy1aiIRC516cdROHqmd/Vl5m9yEuEfRUDYmy
NUEV/CqiWLnN3nKoKIQa5gjS9vq8A2eBvkbX4AcMLciweLTwqptfp4URK6UZvD3W1cKPt0lOsE3G
3CPEVN2yYIYB63eZMmArHPmRgmlwTjCgn4e8lVjuhS+4hwgw1SDKjbOCNlWb11awR9r7Id0Lm4/r
zrS0sawzAh/UZcMhJtb4aiWbsAFGm34KO3GVHkBJv2duZ8mZvxfUu3bAS15gHr/E5xvexJAXIqZp
PZfvRoU35czCIFhZoelj1qGGa/h0EkAnVuGhp6pPpk1Vr41nSCCl+8dn0ES9C2MO3JGtGTUlsWL5
f7Z0si7kamJQNqrAyKSd58P/Uic5FrEVZDw3TYZgve+BAhsN14wxVGRNNqPzh0z2iI11akpV/jil
QeNqMpPULL9+oe9crH+rDJK2dGu9I9ZGEuZC6lgr0jA99SAWTf3n7Pz7DHUQWDlrShMQGjhSYMAk
Or3ANZ0DcefsgHgRhY/Rvr4z7BeVEOkzpfz97bn35bLjyXKTAKvyy3P/NsHTkIcKExJBw210jqc7
oTh8bWz4MXIuSnx/9gsiQ7iT5NEIYLVlrdNMzs+qUM5DpaeaSW5ATEwBtTyvhW7IMIpFgRnA/JfZ
eC+LTQMgHnHHVcjOicw66gDSxgKz0qQDJUNIfGFHD8bi3KJzboQabu3vZSAhRmE3XAEArsaZV9a/
R1F05yN9epTwvjmyyIrP/Em9+obyt82cFH0hMAKQKZKwnTX2DKrGQLvxzQOF3pvvgGTpHY5cO0A5
sHAjEeaqmw7/7OQNIytoLT4a1QFZjz0TY+z15c5eO2lsB5sUdPQ6oMkWRi97T5ccc9mZe8PfJxYY
ZBchNzRurQDTTXH/FTKxkYCW0vqCQIrjEPhRNunRuhOCAc5e9/5M/+7qxyGEh+WbjK6rTUzPcQ8W
s4owFCIPs80syUHZF5bHprSIN6/grg6175+wE2KzQHvEk6NSJ8fw5k0yUWDgZ1/T3wD3F5tYjQ0U
DhF26AWu1OPAxymkt/W/VXIr07ph/fRFhwWQnKMDjNr/J8je/GcDQP6pDd85/D313IdHKHaonZ8i
vBdbPTrJMg3cqeegG5DDAtm2jZatuCUBL9l0sp20GGeoaoSnBVVStm2aSMed7gX7UnD7fFbAQZR7
/e6rZVPnCKE2oCLmL+TSILwCLkbvYXuyX2SPRqM3FBvqRI+K4TtGICvr5Ls1cLQKNMTlDFzuUJhy
q5rJv2GoNTtCbFewaXP4xuROU9pAahfNoLCRXIO9k67OgBy8EF6mPTuGiJFyfOxHAnTfOHHnF1T9
aurZe1XMtvIfEuXWykBY3ZKN7YyQLNkXKrDgD8rsE1NGqOcluudGioozKbZ19/AUj6VjiOG12B2q
+Gsfm4OCz28zJubDXpvjpddUyAbsGbhPyMOJ88z5ZdPmY9gf9SlMl2k54aDPX0O4MKGyLaISb6vj
6IK/oF84pkMNkmsSyIpSsEEuNMmOCcw05owBAy3uX5isiZlivqik/bOeSzFjlD2xjCpyWJESCmfi
hbtmnv1+Wp1h9gM011OMkFEP6cI3gr1BLx+O+Jp7votyrK4M0qI4MZO9tHKcKlnbEL7iL9SNLjdP
nNt3zG8tH6EVI9vm3sJN1QI2bw8mKQOuvc8EUqwgVkgwuU42X7fBVqW8bf7p6/Dq7HBI+EKiLF1q
I10KmmNBZDY5l5ewjG5rQaT/CKHvHv7P3bALfVBtlA4ZDrhtGIaaQ/UvxsNrrzG1YxFNtc24ov9G
ooU4JXi39tthQ2ie+pbc6/OeL0wviZLEMU8WFX3MxcxEPFEcuWwD+keldfYA5CW9ymPAjwHk2niZ
dtnnyrk+ecwLDphbYk6CXKf8DWEllE8crY4shXLgLsvv52HbBtQNUzCCmvBxwFWQ6IvrfVpXZmbI
Ot5j9Eokv7HLXI2CQIjLxoBRAVS3xSNyDCXXxnqugqF1Y3PxHhSs+3Uf/r5bFUPAzC5wtemkiLZD
tya3zotToOmEPVQPBkVRYXknHpkpOYNvcAUfsVv+8WXkKxa6xpplx3qIBeP4kYTprt2u5SuYKbW4
MOdlmFYHrbqcN1o2JXKwX0mM8UWqCUxW/KWVXNva6r2JuVLBKul6glXOjk0xE4RmMoAKHgRnvn8D
3pJyANRj1uaeX2BxpyAPdb9a0iNQUEoLEZQMtsbXaVwVucL3ty/gEsPGeJ1G6Sg+i3jfqFTAZluW
0ctNFtVKVM97YYtOXMUS83AILf65L1o8FEbWC6ZpqZox6pU9qjazktgvMW6rTr6hB10fXzsQWoxS
EPIpgzMKWHUBocvbVMCHzSpUzYigV71q8UvqjrG/xUeky6VQTL5G4qmfarlH1ZSiFkTLw+/4588s
Vv0W6l0+73QdQ0BreFhMJUx72xp6W57Ph1/VfN1f/YxrYSZQ1SlFGW/CDD1QyQtIZe7Tsxbf0n2M
Suow5cHxPhc8YQq7Ua9zWxOoyTZtdBpX+2Ili3cmXnOhAg3zFgorIPumyv91Fq/H8o13xkjludNi
D4BwjYTal1UKBjT/NZkz1wJf0LqUMYW+E8nLIsTSyFaQqJpPMVT4IuFxinMA7DbC5Eed98NVjiGh
gX4e0VW1jrpTIicGa2JD8R4bkoAPYrE/JWOldZM1y2aEUwNI300c2a4qOrzVrDz+D1DwFhu+BlEZ
aXK9Z0WALOFVFQ7Z+8QP23KZfXoeIWwA3zBWiqoZ3w3inwmf2ELN5lLj0+QUI+jxlRWaVgpU22UI
x/G02XbUafxPN6ABmshsC1CFeJ6pjSLFHGt0E0l8TCiL8beAChp1aSwf2Lhd/FuoSuz/1UzbxRsT
74hdhWuxAP1p9DGVQpc34japzBDbQi9BpCiflLyjM52mToNxysTXgHqlgz9jaBlg8QbGbOKMsmic
MtBAEgbYX+toxVEQOKGxIqPmw6NpSWutzkdGrZfs13CyprOWH4p+GYnylHR5boQgRKRljJr5RGas
i9RqyK1/5LY9XSyzzVOWo75qA8S6CDZEDOcxmEWtmto6PvhIVxVmhMxOa2Dj6EYyZF0M56x7YP7U
VtrO8jAUgcvE9lX6ewsEa2B28YMltPz9KanrfZMfKog2Z5yJVjxBVMMgdFGBKNH170EAU3xPjUkN
mTwZZKvrfcJuIjKDHAWsP+H+UdDnnT5qutbQiQ/f42FY4GmCB7VwzwPVQ2GPt1Q8CRXBAKrqb3Pd
YNEirNqujZ13Ymr5p76DugkkrtycDiEVtz+AqEjZ2JFWmMw41Btnv1MBt0bnm7Mb1QsoIpRmpf3A
QkbbrXKyP5RUeglJzrkoXhi8nF/hh+xS4iuqRvuGpEGUfvB5TEzQ7zuAh3Y4iHipx7tq3zHFJbiw
PPP/BsMLxfFshpXxY21T/Mf9RHle39QKR0XApyz4BcSAIJVu73Lb2/JL+rOdXev+1b2y5eNHpw9S
66Bh7dJWIZ6xkIxLNSR0kasQElJ5btGOgpW5GVYwDULChCj5gmOeykFqzj3bsBJ7W1nrKmuO4mSM
wEX1aZFH112yi/Jgd74ycp6AQ57n3pJZb/6BcOCmZlT8CG3EvAtzKDrflc2vBrKYYAL+HqDuxGGp
5tOobXqRy25WpbHNa+BAIxGsyIx+e1iToA5dS41fGaP3EtMaVBFd5BN68XWYMx+hyufQmvbPcQeI
uhU1AVbr3RjDyUzLdhlMPUio3XO6vceORmKmhoSKY8kcEACm6l8AyZ7vsKNVvncGdbEsqyDgZ8BE
S/+NvHC+32Kpo5LjvL0KhD4idWCxUA4Jv7EjDgfGeUy6grut3UDtLw2PRf+wsVaXuZzgeIv3Yhqh
AGwv26rDHzvlm+lNrN0siuoqf3Vkh3qPjEOrUDTSF1JfeaIqU/N3qFHtOdYeGDl2WFpiGEytdAvf
idtPgwZMNhoQN1f3u+Bw3AjcWjfBnMNIhgwm5le9Q0uzQTs+bU+vlZ5/8AHVDNkK8THAxddO9NgY
3OIpvcM+WGV9U8D2WyhoP+Rq09cmdFoItXQp5QxNzK6i3EkDiAMbzn+lfvfv/t1LlL312QziZFbe
EKFADhuDQXoiHVDyMfNZ6nTbteGVUDNxpX6bB+9lOCFBgbaYfvoL3SFKHQ2TvOM6s8c/dMSM2fGf
uTPek8BJjZt+DfvXE9VxV7aljBcVTc8Hdm795bBAm8N05tk7iC6Urwy02P02xzIKM9s1h3gX0oLF
wrfp+EbdUmKbJliE6M23BcKk5xrwSq3i+ZNEsaAQd0nIpc5TiMSTtQSSLdCrWidGXpL00fnuouLm
hbsgWN5VwuQ+P4HxpfJLTIFesBsuFVHZPygpCmcz9qThKAozHvLd4oBHIjGfCo1imnGZL3+n8HG7
DAkYov0avuHpU/mVMcXHyr3/Rfkd+2tQulc5IdoKqpIkSyfh7M4OBdQ/je/M7MzfUHR15ETm9GZ4
r9l0c6kmKBxRLYGZa2TDk6GJ6nU8NGv6nfR5+OuQz/aSxE+PvBy9oNJJboE43xpX9uXIKd1MaJ62
HYCedA5QqH29OMrdqNes2bx02W1hgApks2xMmYjI9jBa6cqSfXb1/yoT+a7zoWjY0MT5cE4pY3Ia
vOk5o6KAXFS92mqikqRzfMQts2btgC7sn4/GJKJERnzTRJlUdMgVFZIsuL2oXDIKzNyUxtYDujfe
7Anx1uk9AN6KiCNNc/kevftf49wnd26k4PS27IOiM8sPQ6xha4N81Kyn79ki9mOs3Tte+SOSrtQ4
Rp/9VCPkbBTJnlVtsoQCGYIUyhB3omlF4IvNM5S96pldXENg3eR+ZxfQfMPRc0w2SPCAkrbbe93n
i//oDenDlb5olDkVHJGBVtOYcC6bN4kOYV3MBiFYW3aODxkTm+otxXS5EsxfvLqd9+pbQcCEH5kG
hPzMUNOuSNzNq3/wkBcxLj9b7PI/EwyYBS4797p9qsgPcxKN5fmoZJY48zgEaT2ibUOo1dxzToZZ
4v0vVOkHm50B6Dn+Le26yuESuIL+c7GPyxxBwa912sV2zC1PRajbG4AZUgUoB89zJSiZ3yg8srqf
q1Ek+GB5gZJ7yleqCfQpwnxAUxFDUOgdUd2VAqjtzkTfjyKRjFJ+xg1oMDdGeswF31WvN11q9sJW
d2NEKgfSzIDC4Dki87Li1YwYtazTr+LBELnR9Llk5dF0dr9BTne55phnNE3vte8izaPsjWk64BEB
ujbQD8XcRTm732sqhzsmupYRGuWcSkSCgah2j0oApNXOwkyZyFv7nUPyuIIeuq3MwmxtVlnaG+cU
dRdRi4xvI8Op72Gm+bbrK+OK82f9SVRy9Psuwqobkdl7rJgnf73d4UwIOfFvyr0wmi50VaVvbw5Z
Qq52gcQdex3AqavSMM2R4zQvh2P7mpKop3h8kiUj6/9ArQcUmqiCN92yFuKqWmHZ4xpDW0sYccSh
KBSveYEEmqfUG82DhR7cA0Mawbqxn1BOvV9HIaKdVdiqHeBs6EsXxZreJ1vLSRf5EgjbjLRFRR11
JgOA2ZMXFlqh4eqONqS/D560FUbC8doSxZkAVMwkWSXmD531+9dOHjzrhcLtc8VOqjHEiM9bTc+N
1LkTOjmFglCJZiPnvCklB08a/RxFTWeM0vSfqglXn7wv7AGrVyuelA9agCwzltcgZ6jk2w638BVD
yE5E/MzJ9Hvlf6kmF4V+tMXst8KayR/XwxY82hLglgFkIpDzjBlYWWsO+CRqUI/cDR6YNNOuAHXz
sFMSeWLHjpSF1w08AVwdV1Xf5GCzZVmdK4zeW015l6Qlr9ONuKOTul6aXphZOZe6tM1e+6KqTy07
6XU6kyY+nmDiIg50KtAafNde1DFfavnH/CbIfj+HtS7q++QBUzipyR2yCRc4T8g6cQr4BlqPPskn
AnFcX6W4WysKXD9JflvDC5k1Dy6GAO7b6DTz2RupCeD6nhRy0ljfJY1G/Rz4iDk8BPdj+eNpOZZ6
9eorvOuyJJqqMH86ozZy15tHEmIz5CiGenbgIL8hP0QFA3onh/brKFOeiDJuYyVof96ub5EdfMKo
DTmcX4gKGw8X8rS1gCCCg1GHc+1lL5qSA5JHvwV7PReQf7f1NbZI8a5UTvFuiyHIPiGRFa/8DFSM
RzL9CK3rCt/SiXhoe5A0g9Qzc4TlaF1n7xQTKIktPFm9Usr0Bsj2UszsgOZhvww5VpjxU9VhMDJg
96zerSgL+YPUtHCbdQEdkCzsGFQwmjgALouIJ5FKRdaPKknKMXlYLeEc398zJEH7UIyvPGU4ZNxw
t2CjSjd1DD00g8wHL3TCZh8TNIdzO4AEwcDmolgLYorgN/dIvO7TaEhTfr2l/J4KxR30xsEsm3RF
JInLw6CuQef7IpyM1YJaTT6s/EGQxr41EEFTi0oPyk0jNqDdK/M9mFy2H7DZ8n0hx6zNR+h6thm5
q5mNbnSpNnV42PoBBmX7gBRFF6UWfWtMk6xeheZUoPkUL5POSwFqXxX/y2YMY9c1Nk/Qap6UcKhB
6JIrAofvexZ/wFemPstLy7QleTwL34yLiN02LWOoKJJmFgyOvOdVSFzfiYKPkggXE2q6kvkYTMvy
Q+JWmuC0PeeJtYGsshLHXXHnmRdEx11r0EWkn8mRNnVwDbCG3OLSj6vtFTpeEXZQZ9P2pMfVmIhr
1J97CxTSdUm3qUiqZ+bXSAooJ96ZWXi9ZR3nkpR3au//A8k6wLkLv7Rg1aNKw3r9ItOJ4WCmFDkG
73+ofJd6yiB2NzVmV4jxypQGtAe4TgnbpGEa6BIcssiTfAyN/UMwTYezHZKdMe7q5om/ET+02K08
2wuO8hZcT662OLQ1hrJI5+1LicolweoJQSJ5TFFWJNRROhl4gAdBIqlVAEVlxBmCYHOdLEhagyOs
EHIjicmy0D4iFxCRLUStISwPBLjYzwUV6a+eJGJwEnWBd3bamwza5+dzIeK2FDZ34qupdZM3QSwO
qukaUNZWhPz+cwB2GnPPGaaVUD4HNuX0xil12usDEkCJlVJvBvaIJoNzj1iJUsOdy3Thbw0JR6DY
yo2iZc279KUu2u3CcVIPFhELxArQHyoKvMIo5VuNMGfB3No7seD3tAf1XgocPO9Qi7jA3EW/V0uk
xPSKFhAUu51Rn2pHykdAam2gsMSgvSuOV12NFRghY4wnspZ78yPnmmU9VwfjSZ9LrHb7iC3ywqwb
fjsSEfMjjN9hU4uhVU7RXPmnAnWLhPEpckMaKvr4IFrDHE7gZzEssq++Oirn5Y4XWxLCqmybYjiP
Qly9XqfPc+L2xxKylaVUaWBxxuV7Ila+OEU0mZb3weE1EK+8GBqi+iOmyLMNsFJdd9vclHB864cu
1HBdRtHVaWHapT4502gwElVM0r8bFBaQa1wr+Fwk77opDMnSXhC+wIDJe2oB/0TW0VUYTKHeTPMt
T0MJS8/enKSLcLJc2w+BCOO2a6cxjnS9OCwa9CcDnXEu18HGlA5Yi7i/3JdoAmjAtUUdVPEZHSV1
hlhkTCFsQOwPJkd/wsG+xp08puHP2Qs4oyGk+aZyPd1oYBI4Np/cabV+8r9+BjIFaHZ1Xxne+Glz
PxuOlLqWxRe7M5n4SKF+uvcdzsoOyGnVkbGicVKtKKUrIv6IdHgFOdcB6EdPYFl3dbnW0WeZC37q
X9bSrrJcFRUgf8zdgQA/j7Plejh1MYr8HXrmkblN1+IXgVyUkKu8NoETHtBlV6JhA7ED+Eqcqkqj
+JkLDFVL0+hcY4G5LqiLqW9NqKu4NlvRvnf1a5nvxR8OBSpPr8VEMJgdpOrPCvvF8jQqgIUt0Hq3
+IAeIvU/tjrYdRcHl5A/sZfl0oN1mFZGHdNviLvtm2Zz2XQ0qv98NVhG56vuHdevset3JLTTsjnz
Um52bcq1YPCGpJiYZPabzIDOM6wrRdyoC5p/pqt9Uou9QlgsqdT1BhSDBQkVZRMxUksDcvpbqKbO
9LM0E1ctftb182G5YZmCAJImOXeT2XE2VSZ/D4Ex/AMNMNfhPgWtMpo8fCJBiNSRNeeM5h+Hvegb
TVXxKVblc3Ixfxif8xD3RcZZ0nckx6K36w/wHmfjPNjl6YLXMQQVE5jUxAHfvTjCyEVVPxGxKpn4
+HssmiQgm2ZEk/fkbbygYwcm7kvseZsS7By0dUmN13Jj3Zu23cqryW/uCt6gv4OwH0ZruLSNAV+0
tZAJi7zYp5Xl7f+ybsMa7k2Ss2Q5M0qcPPylX1zy1+5Y5wbQL9X4X37VBUqsmmiEJ/25yJdAhO4e
8Id/wPKHSZNgGgUcW2xU5Qp3Cn8NL9jpdAFxwlFOwzVVGTinTyFnDZUWTLlYNPguSrzRHBmXVWWK
YQ+Ft+LQmLDn/UH4uIbZLzi+V/pmbDdW5uSQvcIXUWlXnzlFNsX8HpqaxjF/ipdI3drcMWk6NzI/
fcGOTuucxDogQ7kPipcv26lFnfkSQG+5orGreQe88BOqsPo7OEQzEkaxHIREIvwTNKUK1LbyXqxE
bB6WqueT80/m9fXEpjhrEGNiZeRjgej9FO/AU/bi1QKlTj0/IP7yKGxe5wG5xonCLiQh00M90dxL
EOaeyHmX/v4/yT6m4VVUE0Xryv5boI20WAELLfUAVsX/CT2UupXKrgUQIHN/WdILdx1La60SuGE8
MOHyjJRCwlYtHKuTx3X3pRGeDxLLmctLDN61DNZ6VUSEBihHDeFfRLbz9P3szZTUcmQ4O5b/3v6w
VoCL18CAcp2+JKC92z9BEcQx4G/A+ov1VlCBhYsdU1KVtXeUhMUI4ujmIlQNhFql4Y5mrQzT0VJH
g3SuV0fz5GZ5THg/4W89WCvMecmEMudvn1j5t0W3IJZk++km0FLSLRAM5yWCBPGl/X08Li0XdaW1
Tt9eVW1tZhd1OrHPibb/Pe7tzjJkTLRe4Vj4smamBgc2jTl4pB0z6UwQGkDFGVS1M0w0Dn4Esltz
MLrIU8KZcX4a1Uk4Fn7DlrDfZhiamgiUJHufVTR4+pAfJJOLlwjEDC9y8e0q3JoJFVBiHqebQyj8
6Z6o8CeDUqut7vA4iulYlrVyBLPftpO8oFWbXdVXPgoR113A3EZ7PEVgSP8P/9MH/ZMLtVj76IRO
0U/oWtNu81R5H7MfWpEjzEudEdtLE2OneNnzXh8kGDT8/PJ252O1x/wS4yoyMJq2oWOXEjyH2/vY
Rw1bjnjkE88nu4diHZVMSE9GJ1RhJlDFzOX3Iq79DLudkbtfUGGIH3fv3XZW3t4U3KSPSrLZXSJC
ZCjk780ZTLPwsAP9l4m3kv5uOmSZ6GmWHXnzBRCyw1+PP59cWGLi6bqPQ5Y15kMGOQuYM0l2J0wY
ttGSITQizRpNFjP3zS8cmMnuUtGrvrZ120DSs2cZYR3KErDvEoqKa+MNXnTP8x8vvtDIqQnct44d
a5uAGcZFpe1ClNqQCiaXatPTEMVB9KDtJDF/1r/wJqp9xUz1jl547kRwqxqDiClBboF10goDLE3K
SzD7K/LqbkNyo5t2zExUu9+9M88GXE0ayjLOEVO0vkla/ZLZFiPXqUnX4NUJqIl1fmE64u+gEFkv
evNReEHsv/DXpPHaILOaSpqALj4rzQJfy0twbPFKEFkdbdvYXmFkTBHQDmCwl15iBU8imogTdJ8P
6HeUzf5JOZSJuYpGx+jndU+m+BpZM5GlFF90U+H2y9uaCD42QN3eTTjJ8mQ2e0b6NwBs1F/X9d+c
+UfV8kO+72Lkv0s1Ejw0mNjL55+mVikTYfkbtHKfU60bn7D0/mlpicN6Qp85c/bcs8O6GS6jYdPF
NXrIGCcgAkqTGasH16FFB8cRKVabRiRcBNshP4vrJGbzYXFEVGfPDQTRC0jDCK1uJWo6CqSMo5oP
E4fbAthS5bXakH2OFoPecffIKn8h502n6IPPvwCZ5C1DX2dyuuzjZPVXDMnKAWM5xC6w2xo/Cf34
0aP0Ayg2IYN3pGM1TU8/f4PtjNy19uhhIREzdJvDQa2mfOMFJG8Bav0saFaBVlue2QK/6CprASAi
ijCh15Fhe1auL2bQ63EOm7eLFh5W97bRd/pX4EeRD2ze1zFri3YsXgSmNxTqexHzTzYYPDjapwES
FkinF4YWHhW/jizA2WTorBztwDUD9XxXgAc1et3bcJYU2o/wpFWUmRB5BXOOTwwqRhIK2pS6cmex
2iR5F3r2d98GE24B90d1UiUJNNZvoS407LHFpW4DN2yZHn+4uDOZy2mz35P4etKgxOGI4gRWpukL
Ka/8i7m68RJYzcYSQPkUeSMi8LXYAPlj9GA7/AZ8d4SlsYjqNcTZqQ4EbAWbgXdxlxW2y/69ENqz
TBd+5yoblRl6EcVQhjWsUO1AXAR+9rps2Qb+PmosihZbIQeFEICCBZ2gd396QRuSoQKVd3O9qluj
2po2JmN8ZGltWutHeFzKQMwJx3HjBtLuliP/BdqcF3P/CbUSyi4JzC8ohhI21MO07S5AATDgWJ2a
TkTHJ3BdnEkpbZlse0iNlwhINpUDsgg3XcWFycq+Evx9G56AyMKIfJZO+QrAittkgv0vv9DgF/HO
MoDsCxVvpwNZakVA/BqN2XPD5mX2KFHGcKhGsKsy5zY+h9rjIvjJnGCXaWMW91l8SDA9SKkg28FY
EbofCLFp2RvXY0w9efTezsfbJ76/C6Nr+GeMulg/Z9XwMvYi23X9wnfFdGuZfMv84c/4eXaFWMp5
MSuVzuQVvbKgP13jiOm+6MjuWrkvcBlbyf5K96Vjxmz0Xjw7OUHqAd4z82YF8NSKu5nmGk8fkn77
4FCgNaDPEV45+D0ggxh0la97EGLt4BFGRNODiT8E3ie1iIyvStX+vLWmdRsVAgqDTZP+G3F3OtG8
BxOgNy0KLHg+gNHTW6Y15zxzdlM7jB4TE7ouuqncBG1U0pMJL0Rk6iFslCwfofdUX0DG8cKeUzim
mwKi0yP5BKtRe7NDkv2kZnhCJIIiJbtjCZUdyp+Drv1hgMzsDP7pzi5rD4GcCqwMhxhmYh2XNpb4
Lxb5lNgceKd1hNnn+UsUGe3IPQu8mHdnguKtqF5MvlHOflGBh2WqRkYXdNKWoZ5y6y6xdw70FB11
iXob+AawXnn1a8R4EorzQwO1KejGjw8udPj2i+qKKJs3Lfy6+XeEnoSa/OrvCX4uudlmnj8GKE0c
v4D3O/l8WIYP1p8UlhSbjhUBr+esV3OURP4vcfm+ykAeuF6/8NyEX7E6ZwFV0l/PJvXLbDP+fzqj
kpu2MnqJzXdrlCKe/Mbye3PMIUt5UA/m7nShlPUO+/9X8oXXHZKEFAnTBo5U/cuj0EibcBShlLYA
nq1rzjmaCGW4RDz01GR5+rgjQ49ZS+HGYq5psBRjVIAhF/RrsNPlqLqA5vpgvpljeITNzPWCZs23
9JJIlwJ135HaDW/GZ+7AQVzLEc1jnbLPHiMOY3pQBURB5yqLSoOd8wQAsfqCthcK3jV1QOceXQZx
WAVOvCwbkJF9R+QwSWTEBO0LjBybnmrZ5O82txo3MlMUanFs69MANKiYXp06VOVhtG5b+OMKhoOH
yoVg2AY4m/oq6Fel5ssZ+xzj8bp0kBiaCfA2lazr83o1wvsezkTYxyHQI04QdGkgPKfCOSfaA8R4
fdSdQL6idlgxyHzVZEYOMqEYMk+7Y0SHGlTe+e4EFL/RTAjHYzT8HwG1Q4cximFDYx+AWepuIzlD
zarGfMR2KjQ5j3FrcH9AKo9MITdJrlhmX0DT7Ha1XX9iUMzR7V6uPrOtCJRI7xu7r1N9XkjqQbHR
RPtk8uF49fpsgrmcmdGKRs6WOf10AAj+jE6msaOoyDwd3W71R89mUwiHpyQ1q2yadVj9o/YKS/m3
ohbBaaEUiRoJ259i1MSlOG+6Z0iADYdildrnzjlQ+G2c7KLbr2bm3Hd/arDXn5GocC34cbozB8CD
o0iE1yEk4O+ymwiC1hEfOQtfdj+9Sl9YhpyFC2eIW5VByLD7iiYoxC4ujK0s1+iZxMccuoqnHybp
VAUP7gCcrkKmdpxDhsjbGg1ry/Kvx4bd4ggQgtGwh05xnQ1jiSj99ngebqpez30jC3bZAxpja0sz
ryxcW5/mcDpwn9VAbyeoRwe/gmsTdGrjRCDWB3C1N0G3dGYY31XMKRvhuvnNX5dogNHqp49p680o
8HOjDD8h9lPcMjMvEUwvcnRkA5dTcIOEN6Chsdu4BAUb/ThAnfuq7KG4KbNaHqtc+il1iBWA3nwD
nsMgbNnDKnx/GxHm/Kz20uNlL+1L9CkRaHp//mhRkK4RuRzGxZ+uUv82mhIK06GPOl0GUjxNUgpO
8lwH0bQd54C60fAKiFpzUEgNrOdBFGwPH2aizseNhhyHq8MMCDjwtC7tnZdyBHzC434Unb+jE7Ue
8QZd+782clUsbfPd9CVtinq7/pHQgyup880UTkiRlyOHNPPmvP1mHTTiXB3QPNn4YNxw5UIPpFb9
zkNpVL6yGuriiBveiS50p82U7i6An1s1hU58NYN329SEUjG/PGn1cnoAdPr5JtMLfXb07tPwk17X
DMsDKLHio3oEtgFj1BPRDUKkHL/4FvfEz8fKnhlojgq93Jj5aXMq8Q6Ow4WrntkFXqzzdcIn6uBd
Q8VA/7EEW/IGvL2WukZPpv8O7W1csygVMvP8Us/qfIBYgZ0NciVlOTrR56RNUUCF2rMABkN74sE1
mn1AlDZPCQq2GqhfdMY0v22rk69P0S76vL6oRxyfPAouNkyFK7XJegrpL/mYPNcX9mixiMwaQskc
qZ6hvA+2G3eLAUpCy+60K2wYkkc+3WcFU+2THkxV8rx7E3k0Py0ekiZsB7IjhbmlMnSlKQ4nccQH
JjEeLmSqEcFQtq5tMifj4By2oJKzq+oMrFGK79kQpxN0hp3Mq+pdz381ApASmQQepLhhkSgQYzzm
jrgDf3p7RGUCvX13U78pMAle4dcvEcnLc1cmckJX2Wg5eazi27nI1KkaLYvG1imsJrMp1zQ5IE3Y
Nn+sqYDtMMa10T3KIqz9huivaZ1c0i6j+MmA0w02klCW5azkeP5mN/kNrL+iwEq/y3rf+G7Uc1oR
edy2Cydd/Wmyjtc7JtC+muUNieyZ7aa5vHCjVbcLJvPrtwTsxlHlqVp1OzwPaIP/KcNUsW0stB9/
XxtE6T0NTf2m8Ydnsol0e3tSi4OF7FHElzBbYROcfK3Ee3Obx+mftfqmNv65XzBT8+ANkx5jIy0t
qDRkXCZX9tbbXvTXTnK57pWQO6E5EqIQsRBgORJEC8SpB8O0RPC3wHGRxLn1wxRj2sF+Zla6bYtO
L4Qsxp36+JbHQrHUIRRjMW8gfp7dQCwyvf+jNdwthk6OGjW1xobisqU03NsiysnV0VQ2ySfGi+ta
ecGmMa7nGXbJrM61vtXH5/ljbpHzyX3o2RmReokYjDkX6E3lWhnbKFZoLmbX0zVGEfi4Rc4LjNnU
Q6GpXbVR2SQXKVyXJNQ8zbryyqFyTGLosJZDidv/szEHwX5GIcXkCcq+8QPvC4I48XhN7riCnp3D
fWZCeVCvYEtDNGrt3rimD5kRyef9f73sYDlX5ZYUKNBUVuqyOLIvaqVBrlQK++7eSkwJODvUerG5
P27zMUkNlPqZY9q5irW7xWY9z3YyTC3lfFybOd2b7unuZo2ZXYmATHs8kJSCaEE6F5owO++LENvN
dy83RuKvYMt61dWe8I+Sjxd72ycea76NNBot5Nk9OEbFUwYYLlo8Ij+VVyNzZL49K29EAirmTL3P
RDsc94AeZj6DGtMzIf2Cas8LEetyrRA40M00jll5JX/QSNOmjbIFIzGi7PrV0omSnlMk0nAXZ53M
j5S2j8CZKDuruC0HKOceD7NS3g/61TF59yPf5rYFC/ywNz6lIY9/X1AfhCaggKXLRyWQpgDMh0Tt
9dyKQb+ge6/ba9uEfaRFlBs6nv8zV0q+HKdkI864waTnMsLvaJix6aBkIS0SPALemsehnKgYAYpJ
23mq3JQByxuBWGtwSebvrjWtzDwtA04AwDlI2Yj8Newmsx2oV6K90ctT8Jwaiu8SCapxgs8h7PUe
c7sSui6J6LXn6X6RYHWccbhzrN1LHsjYzQ/a8kE9rY9etHBvj491uBD9cJDae15Wd/RnHJoWRT3g
86wy2JTdPEnU7UAdL6B+tpIBDIghf5LmYKDWAew99TLc+zxnL+xjr0ywsPXSPXGgLtq46JHlUvYV
uEoU6quVLuvW7mOWfQ3JtPX/MRXpIDbKzow28jI0eHyR369DINuibzGzDwG9xTStVfLa6FAzpU2L
jp9CO3GNRyyP39VosWRcbdY5XooKayY3gkMm0MbO2pwX9rIFDVKTJ+h1ASQyy9TmYO8gR3R2I9gJ
eWXfOge2C3tW43HsqlG3xskyTuS99Hf73i+gRGoClNvjTw/PZoJN5QaxijB+Q6pRPTjHH6n/GGAe
luvE3GOROQlnB88+WfyxdlgWuJffpvWd0yXHNhkEizZKl7H0yzm/iXOYVwNB4flPYQBtjI0TtEzS
D/hQHxBaSE+vqi4MXBLaZWw7xkrpxxwdxDq4RoEP/xi3Y5cbtC0TzB8JZaRetrf582eYd2ze4iqo
vCap4lzDfINq29438lomgVXu3HjsXjbroV1adnU0n3ZFK4j3uHV64l39aQfB/3bVur+T7m4gpkcV
gPO2+vG8ZI3k/GHz6cTJTaQb4kQFQ0qxAF7wzl1fhOtXD2nLpod0TevCIfjJALcYen02u5KTn1Bk
rXBJ+fYx31WTmZtocuOzhgoppIDLHl1TZA3kFbSwba8pfBcvpfcgzswLlaCJasXQmSD3skExrLJk
sQWAe/lWbQ9EDqR3KypSDVCm3u4Re9HWEuVke7kA5rRQ+WslhCRoz3qAGDmO+rXdrzWmPyFGOMFm
lXatt40g709RbblbnWi4qZC3+UV7FIL/8Hx0j2jOTKHXoMvPicbmGbfUjDmPx1+1XZPnAB85gZ3L
B3KW5yyp08BoN1oeVgA48WJfUeEXwwN0ykPslZvasru3mAajQTsR22Ez4MFdRngGpPRxDqmg4bUv
FvGXJsL1RH8tqcR6xSpFYBfZHrC8wCOlfSF78l/J8ELStZP6RZQRIwZ2BvseA+db/4d7hgw9XOan
HNR3oGyuXyG1qyHe58SunPmePcENgVEafCELoGowdWP6HFUfyL8H9HjG2S3VGyyeEbJF+OOJCyua
Na09sUwfF911AaHQA8ke16AyEwNkS7ZQ1/DBpDgkvfZJ2r+iCLpRexYe1BAPyCECS9+a4OWh76WQ
3+imZ7f41AKjcL2R39oqFlb40wQpc/so6lUXuahE+J+X0tgHDhmJNIMhaAQn7wVJKZlRcyCZcv28
frtUJ+DycZfSBvVxoU2OsiGtR3/r+S3crzBzDOmbrvvftAjmIq3uqZ/1Dv4ooxDY+P6JCtpYCQa7
ZCDHa59u+2/VmtoV0zOrdj48nd4XgocxoGjlFoC7O8FLWZVmnqpDFpQRKvUAQK4pAUuSQAoQbeY3
aBqgR+JGAvcI0SyS7UT4HxgXx82qYf9rQbns4SzNR1vvUCfm8Ofx65atr8PsJiZUvSKtc+njb8gH
80ULciicE6BRsJUZVZujv/Tv4K51cv7nocDhEYerktR+FK/N/RQim051wMVNpAtCABVWKKRbGfT/
L/jvGw2rF/y5rjCzEG7haMc4IF42CpGlNHzWqVS07EbXIYUwrGINxWylgvfGSfCfOGhqXKDuQkMc
23rJvK1+VPU4Cp6tvyzBqUwQ9rUemvwN0umHsgGsIN8BRwoJwp0tLWhiTHfKV7+GwGa7xJwqlnvb
RzktyHdlk7CNB7Dl+lL+WzGcnMZjioBtDQQcffoKh0MaozqClKH96DkNJbzS6S3pTyj0xCJ/bTmD
8yq+eXf82ODSarL+U8yDaMu/HkQkHga6ePA4fDIh6qA/gce5t4PkFma+wGXaFpdbSYVbv4JpsUm+
lTvJFD+QHjKzvBI2HnImgBf0YYnPnkr+IHScQWkz4ddufZHCVetXj2a2MGdau29Ud7iqkzH4vyYr
1XPYUHB/PI7+1pQSPrA5cO7j8IRTtVcy/CFVZD8F1d+6uZ+myxn1KlFJr6w/DZPLKIU9HUfgudh7
XTm0DPu37Lxt0McOktAD642itynZVC3GtAbwM42BbalwbZS+bRpgs2gViVsEle7vt1Da1jIlT87x
3YYAEmQ+VqYgCyjPaCShwniPU3Afh72+nwOA9atntC2czTk5zLe8gtIBmZC9RXCkjvxy5ciCwVJq
6uz7VkPllqZcrOheu+CnCkEGClaWfsc8zFHhb/obxAMOLkKRkgCLHAnNQpX63oOJT8kxke/SaJHT
BqpN8UeToabkRf4FW2lEpedb35Kvx5ZurZ5sFhzt/Bet26jfqMGdjclCs0UA7jG2W8SZ6qK8e2hw
f2xYgBkI/vBDzQRW4fjQyAXaaFEEn9uU0KXx06AzMtnX5Bv7q2QIgr0eTIM8+5o47WGrjKCW2FdN
C/TmvcunN/bHrVhWuNGD9AQoIybfKXFL6CQIfMiJsBFj17Dl1ZRMa9IkbAe0ywSh8zUh1bXhtGU3
0Jfdnfr3izPDuxr5miGufD2CiZHySKZ6d+otFfTiIY0dI5nhPScGFcm7D+FNuxZkVLCzUr5wLI8G
NnlKYJHQx8Yg07KhApbo+kAa2v/wqTxYO0d+G0vfE+2odbKKyVTRu+I362tdCzJ+RhgRqCi/loU2
QauqgbCS18hXE2DyQyvC7733w2/2sQpN96OIn0tvJlPRqSlUAgV/wm5BB42RHCWRzNDSo0zAamZb
/Ij87eTO+fbyvKflDLLf68xeqy+y84vjiS9u4lCzEjMmQ1HouzZOXoB2TF3xrxzlHc5b84JcsTpd
V2gmx2xoHyTdy6lns0q8RWV7fFoQKC5/aBCGySeqJUWtWhWzRCUsVTj5VxDqh1kT55hQxWl2qcAz
atZQcoBw+oKv0w+y4H2tEpw680CO0+ruygpTEIWqQCW7HmQ22Gu4m+NP6oY82sE52zxsoR7yiego
44eVV4WQgtHUm5LuLH9DSfug27hz4iIbWHO3CR8p2q0MsaNP8DSUYYTiMAzENEhL7kyenrq3o1ya
tJbIwDhCG7dRBLfh+d72pAOSYV/5gF1SV4nUm/6CeYhgUaqq8mGG8W0LNWURArYchrpu+4UFyZSY
Hdg/PUjdUHAfdVLumLz1+AHb84EpCV3elBjqrEn9fy9kDbitU6ERiYnvwkrU015cZjTix3UEfysZ
KN9P0M4G0QJCwTmXSFPlV+K5jZ5ftbMP5MN6qS551Oj+K5Hn7cKjQKdCUFxMTvR+qK6VdcBVjKWL
3DV/a3SlVLrih+mUAIlUgZik/zcoPFxDkilXTA5loznIe0h+OW07zKhrxhxZrUujVVh7UM92BG1D
HN8xeuTPgLpIS3jKN5k6cYDA4pyY6KSL6n3acGiJ47dMMgwBibf01kZkrUIgz16+0wAkmOfmmHet
N45RaKG6+2pQuLvy4M60j1Jb3Jw3hEtgBoL7tTOUfOZi0l/EDYDVaC4UoOQVPYtatFkkXGc26uRb
6TdvLSy99lgRS6hRm73ti1QKwDESgRlI5QmN6NC8a3PNPcvOCAgRQ1kTvoinYvI1zIKesmHanSvZ
P9mBG9b/1BPRH/xcTX/0uoC1VSLymeCNFA3eg31w+1bGzGmbELbZiO1KSlIyDpiLWO9C3BHww6nR
TJXEV/uG8w8K8Tlh974ZQSv4TnD6rSEHhaobfATjSypXjG/ZCvAENiYIFbXcEJHw8hnJUPbNZr0a
9OhNdq+obEDV5f8qokP39e/Op/BTOb/sbQZmAKKV8Jp+TB0DdNaeVcsGvmtCXIZoxRioRwM25aSw
ElSMUihym2Q/038M0fu2YlvdUDiP7MaUq81k6M4STBquP5aBwyfdmCG84zIRZNXhz2K91DvpoQI8
2B/mVhHUZ2KyYFq5bmoczCCcrCj0ZjMCDA9cS4WjzVc8NiyzkDBC0qefF/N518sJsI5aHatveEQP
ajz5KGrqYNhwCpezmdxEZCMORj9+GuBOYl81etLKgz3BOxc9Dyb6yEK9w3Jrj800jIesvEQwQv+f
WXh8Aqy/6dRnJaf89oi06cj56IIA6UkiGH8Y3S6uEZxPWQX0Wizk9PNXFlrR4aB2cH2FF+DWNx7N
6BFoz02Ds7+OIxkpAN6vkcfkiAeVkwNxNA04/aGdJwOqXHM3KhR1H91X/LQzGc+gvG5DLqviLPLf
hAEMBR1ISyGbyUbwz2u5oBQM41BD248FXGF8cd/56AwIJsZgF9q/eHBeUv9owfOz7ut2Kpp+0Chd
AazgUWmr0+Swr8/3BG3+IN4Q+ZkSRU6r4uuGrYFw8V29xitZWs4fWlg0tvmiZeIFaVm7GTAs7ru+
R9/mvydEQMEnmAuSSuRJuBD8QyxCiSdwVdn3CLKk+cFcCNqV8VK7jPASlQOPan25xeOFs4FZlt/Q
WmLt+PMN7smapAtz79sGn/DU6L2vQgXn3D2ZSdOdi4/ljSpkn0nFsuG07n8Ojgl6pcY6ElSjZ9eT
eUedPNpDAfLIQ6NVSyaoB8DdUtT8sQkZGH0c4T43Du9XRYA5fZWTFTpLAbWfPMeK8vMk8gB0RQ1l
tlCiswEYVbvRMZ1K5uueQHBGMDLrhVv+lNqYoTwjjGduw9A0tMhUmmuzCvhe/lwgfvF+LLA5ugua
l6xRPDwgq2vBqNbO2/vMne+uLAsq7t2bqPSKmgtoidh6GFYk5jyQ2PuzuQl599pUah8BzWo2fOVh
fVE9VEk7/bmEPIesJ9peHZMc0m+/zwQ41npCprCbMpMeRIk7UT0H3SCqlg5VmwsXajYyRX/7ey+X
BxOfzgDTBZWk3PARVxfwfy0E8zriHEzagqUnPYTBn0JW9vDQjaUU0OiQle31tK/5H7LRE/oU2UyK
A15yTmGlLJ5byxnw7Lu0CDg3fVbyA0/g0Eg4xI6X64l6XJuCmtJ74Op7HPrvAcX1r+qlyfElBbAN
VZmW6LvDxx8UtQczWkImg+wpibipB99GItMX3NACNiQSVhWFZtyXONysl7QQJ4v+FYyekvjkZFCv
FKv6MdK5e+ENQRGcM0HZWVBP6u3Tt01FrBTByk0FRosqnnJQHpD9PPOFFowGmtmI0Y92M1tCym1q
AyagpFegFIqG6Fo8IA953MAfZNl5cPze3ymGkQxXCHH6RfMN5DEVzrqN3cPMg0XUou6n0uAO3hU0
JLrwHZSQJKr3KfQghzuu0aHqWrCfITanamcgEuWRpFPaAcHDJHhwVCJndpyit1ZZGD7xyKfki0b4
pa6cSmF2brk1TaJ1PiWIwpNn+VeM3fzFgSjhLcit8V9o+tmdRXqarSBj19fvWSQiIX8TsKHPUaA6
eqeO/VUaw44DkRR9Pl57ld2JUlyMkkPJK1W4mEcmKWc88hKNFHnkxPsokldx10DChUecReDbFpc8
tJrtzGOyUEajBNksqbuGGt0MoVmzKb5KiBMOwkQIDh6/Dzf/oJLmspZoNltSZg8jL+j96PBZMl5H
wSOrWF41E5RfIKJBK5KPo20W0knWJv99dZeyErOPq6RIIVJTLZSfyQOyXjeIZc55+FIrpB8WzSpt
smgRn5Rd6yWP8uklb5jgo0bplXjxZ9MXK4H3YK2DP19P4yznAQQDRK4kQbU3voLt4s/ItQsElkVK
5Df9K9iOyUJDjmTvxBs8hHC3r260pwTbMkyQcyWzzA1C/13SSr4tHHrBicE9brS0626S4x6iTERR
xfAiXXgXhBgTEMm04iLVaLZFIaBIbizjGHT0Ya2zyoP/z3NDTSuG1ILJNypanB016pY0Bi0hfflr
8VggZRH1XeRBfCIiiGSxQkjCm2Levvg2zLmmGtGpnG7IFelaOUyMgtxkfO0Brp+2KuGZ9mvYcEt0
fdLpQo6WUger2h1XuXcYqZK3z6ZBnxFyT+V8MG+YWey7IwjfjnYfEp4fHADBWRog/hpvM/MO90D8
nVR/BvZwzzukM95eQH75+/V4U0gJrLClw5OaCs+0uiXQeorzxNGSKGoUunqOcfVcQ4Fdb37JsDxw
FSpnLzV/yzbjF94rlWyZTPCJdxsc1gZfVWgaMHZbICmSi82cMXOLkaB0yvMw3Ou9LoSVMG39CDIC
ccWj7xB+zXpISjMMqdF7JONnOjZqrcFCtOqblEQSIJ7uxqv06A2QSQ+wZGthSlpBeQWnkbHq63Ca
6SJZXGO1MoUoytq491LSjBbYFtb41UsQXRSXt0pm3ChtT1z5vge+aqpgYwB3eWxZF5rX+Vni1qOp
HIEqMHBja/C8W6npRh2Yub6P+pp9qqVx30OucUMCwqaOYkZ4coUyuDb4qTxELkOIM2b7x5WwzGe9
vpvA6RJnpFk26zDaz9gYJur5/uOJae88Sc2qY2nc7wiaxD2r9w7TkO0FSjaZBxF7LFVGvtB72PGK
kqD4uVzCX0dArG68Ev1Di5tur82pleX59ljPBv8V+iv27OMKukuYXadmHTYdFuzCdV2dhefM19f2
WnrZjxxQto4Tjh58Fw/VAUNbki3vvsuxtdoE/S4UQ6fxCHk1Ry7ltEWtX716QCT2JHwMQHIXIlD4
/SBKVMmou+iEB4JO9wNZCcVAax8uYOoduYnBYJS/yFdXYN6Adjjiz71YAoZfS2JbS9Gre3GyEzts
+a80dpCvSDu+3QR8Xt7wJAEO6YtvGFp1w94p0EBPa5pfnMg+S5+Gkvrs3Vhlw1SIGcionYleviwp
ua8tF4KD6iyMOY7FMCE6VxhOZDNqtLOcUtrKzjCDyW8By9SF8LoaDja6F1sgAqT4DQtH3pbYqk7S
40m6cK5QJbhbUgJlxZi2RorQotR+1nigVo8yBbe6s1EgSgFlo/bCrtwYV47yCkZECY79uIfUqrNd
wFr6Iv2TH6udv68mA7KqRLozpIInruf6FNW6R7MfaXbunUUTyBlJ3Bt67nBygPwtwhigUa2zdfqU
O/ogBe8KSmrGEw32/RiClFnoGLAiFoPsvpB8AwUU16r20YmlZzEIMjt0AQILTOrkbArdllo3QL/S
yilvhTErlTvn2+xls7/sRZwBk/m23anhsj6WZj0axBTMBMTpfByuvCX0+M8t9W8o3f7XsuAWuPEQ
ZBtuIiIjKYqYmJlWuvqb9+ctA6eSarwNz2eB/MaXXCNYapVHhL1yunFfx8dnWkJJPoRUjHm+p1+7
EYyIC4FKwCa4C0khvH15U5vW+HEWcAe4ULbKYhAJUZA+qRCwOFUqF+F4nHHEV5mfWxEPPRLRnzeG
fG5df5SJ6e04a4hhZpknb1EZLeUNT2lW7gmPlmgVUVXx2B9XSF7dUa0dHk3aeI5FoG+VoSd8jIYa
14kpuAbTvQbfBNeOCjmebNfMm7WfpXQXKuws4x605KuqFyylXxQXCsxZDN9d1IfEvw0UgpbQJ5kb
C/e96oE6TiVi4FqkxlD53bGdQ2BSmi1i8VqKRC9brRZsvGDcvQrfLmtoMABv4a6w33wMpZwUfeqa
pbb7r3orFYh8VepnTviwMZoqz7Az/f6GWsn5l6RribV6em6GYIBJecnbxan+h29F4B7XhVrkeHPD
h5uXPzSoHGiud1ptcbuXWjH6eAH9nYFoHYXgEqKRjl9YWLj2EJ5gmXintIdKoWELPh2e1POQliEn
4Q36rmHE0LjGY3zSPIp+APgZMJ9xvIBTq9HNdp2/lw6wEj9gN4zZauOGtAoNezGSJZbmhrN1GbLr
Pqq/hy4xtWdqEbU/4pl0K1HcZoyXxGkivmNyT+QMAvNrA/d95OAN9SM/maM7vPHNxiuSjsUPxvpY
jxYoQZGF8Gz8hgKn5XTsJWivXAS6MM3cqO98bzBEceSuhxxSTJ+oxFQUb/hZCwO4hFWS5l1FhiQn
rsFIr9cNi0v35OUnLZ6V3d7RP4jo0Pqkxy/p0NZWeB2chpngI/3Vuy0na74CmHV0CIbWcS3493ZW
lUPgBW2SmNnFAkFVoczt0MfgccLkmPhSghjXjZZD1Ab51YuBiGoZ1pai9U794siE08JJN4FGzVi1
3Amo3Sgs16eWrTfFMsW010Hk1l1m/qB3ebnooNtLgbyTrwLdfUmXuHy+Zc9GI4rOPQzPUEcy0CwX
HGJEBmeY+Eu+XVZWBaVMg4K28Co9WPYbcQzf/wYvScdjQZbimnfqszKLh+g0C1Kte/6S7pfGN4fs
noPgjjnEk5j6kZv3XTmMGK/bgUodp1Mh0DTb799ge9qC2e4c2CtVvGdhm1bNv4ptIkI3vbLq6LA7
5X+CmeqiDaSxx42GfFFWxWovIzp0/pI6VJiXfFpu5w7HQEo9adXhB1L5VPTGneMeizYE/hNNLL0u
XHK8vSOK5Is/98QJED8WJ40OXe35VYLVlYgrbVFccU1hoEFFp1Gl9JTOWpYhJCHrx8CZUhenydLo
FQfOYDuxvw/xFc6DSeqI4AfHOHk5RyGLVoDqxtv+rJLmV4TfxXXgqX7UsgSmDc6dma8e+j351h69
ZQe3iOPnK5YlN5xbvWiAnQC7cyC6LwCoEkBMbWOvT5zQCOijJ+rFOoHMyRg/jUENp4awDlxQKmjB
Ilbe0zrzsplNJeLt+/R2ydeNjkAMWvAld+EWzixcwcgm0eQpoT5IlJi+3x+wzfCX/2a4gkQaeke8
igiwy0+kl/0g7IDkffe0Ecyb9mc5pEpPU1DdDCFE6suu7H/0j35NarNWRdD9/GTciSg0NrxP63J6
Hb507BvZDZmqJZbI/fDFhJ1N92sUR6fs+LovaEsM/H5zy0IaCdU891vQW/081ZbQ+zCXSS4uN3NA
KWu4LdLHVV/8mXj/DL23eH/JE3g9aahWPorcqIV6Lvb8e2LS9CgSouSh/aq3lB2a1neID3vEb20R
9TaKGRlR/AIpTLnlb4SBLt11NXO2zVasmZ9RhYOCxJrPRaTYwd5T/8jE6hI2NIkfS5BHezwXtnNy
JXFQ4c4f2J8i9uFzMg0FCX1eQSv/gzkjsa/lj7o6T3w9CXb6dv88G+sH/gwbCPuCDHk3b8xwNMU5
jtByTgWslfH3aFNnQ51lQfFWlYcIUP3wwhyyy/FTWQXzKiea0MiBy089SqkFJx9czdWfk0eX12Dz
AClqhx2IEkVd8ICWGxF71kMPi4Er/Fy3dXuS6ss59xmCjOUwbNhf3BB22FjsD94wxId+KifftxkR
zVIFdjSi6lR2aWKzk+mBgAd0Jkrn5OEcVRxgD4WadiJLNrJV3CsiWss7F46qVmf89PIbZJjX0I4f
CrjWMqhf45E3gQ/iwQE7TMs8Z/Ol8yVn0+ZZz0+9pCsVI4XuicEiasSCXrGlgz45vRO2vCE3Lhj2
H3g3D0zIpx5qgzBRY4SuYQrFiZvq8PNZqUoSTNk7mT6N86jkdrR7zAE8T6zzfqMn9FaIznAFGOrz
5S+Bf7sXordwqfuEWfKeeICjZRUspXKO7qDock2wKxi4MJcVmZa5AbQJMs32u6TN1W2ztEultiGP
09oY3mq07NkwcP+vZoRCZ8NTjVWhZKaRXkeQ5jjxZ79RBU1brg4A6hr74vx13pJVFxnX50PY2KkP
a21G2Hgbb2edwvClj7aGo9Bqj2V5wrGALA6RGeCafiiqFjBjM56OVFfgCaUI93yGNL6a+lIovT6K
QbVXzSVrLkHxbaHlajNp5zsg59YPxlIxZ8GgjuRkvWMxbZy9lnrw+82VTg9T4EGMkZUTTjuKFpxM
3zZHxo8YOoWShXyczou0A4D8RqspXA8dZVambkfr6NZ10ga3q3K4WLMT57uNv3rVx2sfxkl8JEEY
DOhp/pSur53FP5hEgtAvD/q8CJouSEUlxhbKeM/6YNX66uxa1vKjAj88NBA//9kYSwhOCQ0X82Qb
ijDYWXMjO0G5kp7dcTfOKc/TLpxBJnI/cmMA1W0mvwhmFc6TEvGonLjuDhYBXjXOnCv7Fv68WkLA
NmMgV18kYE6ysPbUwJPGBfFGxqKPxiR8fFFcoGqx6MmnCrjptR9k85RMVUsz0+wuF/9aTgrE3y1r
x5L6WUUhI+tmaJS3pHoGy2V62VmkVa87jGLDIDypsePfRWEjIGiHgs0sjHfD64BhR3jD7OhTNXQA
3Y+z5vTQ7uegzZV2x4ve6b5Z8Rh6uRoUWRtRt56ZJBBeB9+354efaEjCyc9Jur89CT/fpcu2lDMo
Fb9cwHmARplquTNVpVNZ275PQHWW5Q+aZGEAPMbLNrnfRkalVPx31ds6TxnOUVDgjw48qpEoFgjM
/aYWRy3qCqEXR43BuPIxPzV5B1odQxJCNC7bS2iXrAhchn8E0wZaHrjVx0xGLJu0s7q4jLNOZi7/
NtQnerdslUNKwzI2GQex+9w+zxUfcpC+LDSr9h8N3YgcFPVMw2sy+fcDd6zrJd/OWFBMitqXj1rE
3YauTvuA49QqEnjnOglDdRLhR3j4HQ4e+BxlCvBFifQkl4SIPUV9yzmtJLxDHT+iXAbpE6FdiZXc
Ret5iBl/gNk3Nyn/AXfeGvcwkJmsXWUB+rY1YlJ5DR14ZKhESH+Z1oVGYIl2cP1xa9R7ep5M/twN
pmfDM5XvBhQQf9fnY2DovKqb5Mbaf1lU+ekWiKeBrbyl6rP7vLQebqCYqZX4LAHvvITohv4lorHq
70TPZ1a/scxJXMiNNJlW9UY+vru2FS38aXAc22RHHMpjyZ88w12fXKkDWI5Yj2BMQySfpNCHP3AW
mIAgldYrW0LCBoTuZCJborD+hf1g794RoYbcZxmpJ97RDKrH+FuG4qhE6ScR/pbafJwrnTkHZYU8
hYZSaQ0XHV8TFbmnTYr3yqL3OPQbenqmezKllnAWZwjhxR5lQKZpfiSL1dZR6G55mAKloiggTzOu
Gc6U7Yw1F4JMO+YlZgzpRmBq7XQfKc/dlJKlDTu1cWQPsvFResCaI7aiNtTCe/4wOvjjoRUYugpm
cKoGRoDBQxwHI4UK1WaVNqdEQt4QbA4H7RB4ZVDDOEm9RHxS1p0Af/cwHq4F9J/mrRaGiE7DC1VS
tK2AFbROPgSmyxgNlce71ahsqiT1akgkgUHODEk7aN4OQWutVMLmH1gUh5lwrwzgjs02x8oMsecB
GXlJQv5ME535GZ83V37EY+q74gARxxBO+0nq9I1qvyyUadqdlblKE/lXV3gnQQ09oMQfVvz07ah4
Wh7qPtuqAwNfIyuQRJYhDCRnbAZQPnv4mkm/0N0VWa9K4573KIXNSvtDJdqDMa/q1dJhYDBWSgfq
0lsHIleeEma5tDKOeDQuw9rxrk03hGqFR2xLdg4v2dRZmsC9l9XPagsq/xJuAUwlbfzAXtNyJokl
JIujfE3mnXB5zSz9CgtP6AkrU+XKqHlrgt6ixywm+oJC+WRZajfGe80JOs1DSP5T3destHRdE9l/
I2S2TQzwjFBck2CuD625yh8fDbJZ3pCUW8AvQQFSSZ2qqbNEhJPVySRIBYPF6e3tVVYLxjscaV7S
P/Otva4I4neUEqG7b2p43yKQCeOXfdJVoHsOnW+dUJ0aV8qlGezLhcDUihrvp5g4zAmVtF/rR2AX
xnCKWL921ONK69M7jJIbj9ILnWa/oQKUHeXRvx04hSNbQ5aFXWyrhTT3z6+TKPum2PQanPsfICwz
Vv2CBh2pE4hhEMPnBj2/zeKffVmAGHq6WSnVQdrF+hJjTcMtl5268yBzyD2uIKRTs37xxMujkIos
I8+c5L35CThRLYA5UlAcpCW6ftngkK1IwgVrksbzlSl3LDOT1uc4uF2OCNZ8AYuOiHjAOMLfs+wx
ol9VPHO4qkV2FFC1GaP2gGwW6fcJXYT61jiD6xlPXA5Gm7zqi77bT3N3wkONtoV/qX6Th7wOPWZy
mXj7b0PQIONJlcRE0LzmDkpufLCeCOkoD53F2vBKBhsa4GakVTbaQnXJsd3mc4AwlWSxA6bU2E9a
mufAO+nEJTfJ0GPv1AYCgiGJWLlLUv+wU2atnZnNzKl2eYQQ8WtBQH9D0GSdgrnihQj23BSuaRBe
bhm/e3Z6xfiMyzs95PuPx+etOwEJsJ2oW6QqYCrD8xvXHYnpmUQGW29YgIGJbmp9qjUkxuh+R8Ky
E020pm+IBcmEWrshRv0bUcsljRiVmn+kbOCvZ/UMtXMbQEp+4mF5yChRaMxBIkTMyNsRGGNAqffN
oxyPhzTusnfTku4+WaIFGRq8WpsdVN4PMRFbdrMHy4JhJUooL3rtnUWNEe/bCAPFZFFpTGoV6Kmi
wM4nm4xf8TQqA9wzsW2ktKzNG64on70BH83Md5clpOQd/8fjo6Sha/5BmJwuQqwmk/nHm9SRCaNZ
lrpCq6FGWnmkgQd6X8lKbAyTQhfLuM8ztnKbfZGjAkhp+GUZx2u/0KLLQl+xWxhPzy+4bOTOgYfE
P7s/W5zOIb0lbYdStOvPmBkxXqJGYulAaWutW0S9fNQvKya2B1/+J2tLKwUU5X1bCDZJncG4SJIM
Hhm50ay2kIq2sgTreDikEXOD9IDJnZmytsa5RlD/tp0Dk/SSVlLUJEo7Twd/kRl2Tvwc8nLqh0jW
FobitOEUc4W4x+gTCmlHscZ+mXpgEMytwbs6K5h5xmrcQFRn8PZe7u6+haOZUNUj4zV/aa5a9EOD
pEZ3zG4zZawR5/i+W13+UgpO3nc/BSONMXEMpjHbpyVvftPp9zjfCDD7sk/ckAeKDyubna+okmLQ
lwxuVZR9XiWn+hSTzXFeuJrcZSrsRj28j50Lg268WKCUQByACBkJF54HyfBYCvYgo0eVB9jFGsqP
Phd2jYPNjBOzs/MR8QVJpx0Z+IlKoe+Hr42VPYos14cX9Q0PINPfOoZHNIQlkhLkmSdVQPX89tki
dfPGCoEYrLSz42MMmxHLqRBidT4VR+aJYCfQ7JAGJq39AlsdRmbKnj4B4h466LcJHthyBseszE8R
bwtxKCmV1vQDpNil5KUrwzIs4yEavPLzi3Umh65Tqy7xbbe4vdSneyGeD5aisTtUkDncE0qAoR5v
hhKvP4Jmo3+/xDefWZCrNzeQjdmFUFC/kUHR/mcyUwhEloXir2e5PGodxn5Q2FgLORnVVIjrF7iN
sBNbwAsjHYa4b3EO1i9Czp/hF1XtB66ZTZZVFoMpTJT9CZdUghyIGWBawcDpx71+H4xE+jy/RAAy
LRGv9tlXIffGUC1wAfUITKnbBzYk0lUhecHCRJ5DVoc6ss5vuUAMjYvQ1L8WkroftQZfkoB56VG2
u2H9Ency6/DrESU8GKGMIb/fj4234d9AG82LSpkn2hvoU2KhRCeNwAoKv6+hoCWKeRcCiqA5Mkg8
xnfADUEtCm43z3ptsl2XZ9zxy/oDEg0yT5vchA9oX8kSYzHGU40xbFtmQZVJ5ATxNkQc7Of5+M3Z
WgzizNqvjtroqiE0gLMY3KkbEY8G6ObdVpCvQ/RR2bmVwYhSZ2P9nNqXK/DlII1SYgdQWNf1Belk
Eup9fpc1MpXQtV+AF9MhGL59l6NVM54ZtZwnK3U+DwkKajkngE5sAbD/0uV5DfdaP9Ll5WzAevkk
L6nB+aQp4eQidRIsgSdQk5rUHbWFmG8hHNvA0RcCOcAfgUs+iIEaMI6bDwEf0off/jfQyx4hFluv
srOrclX98/jvktC2j7MS/W62cWKizh/9H0w/+UGAeLl6pgjcbk/0vKJxlkPga//JprzSuQM3ycId
56/cFFM68qfJpq42aT8gYmLObUgVBQij0Y2Xk1LiOnqztN76WES+dtFoNrdmUIaC2j0OjaGjG1T3
qpQRzTGa+kjO/agDqBDwvbv6+mngTD/kSJWXhnj2ER+vvSHE6+RVpUxZEF/b2F2Lf2Tu7Y75sSbz
Jg/7LZxCaTs7+wR13BuYdISpncAfii68B9h94VgVqsQaDu1nr4h+xHlqVknXjX1M9YolA156duQw
5qa8SjcXcu44Qnng2cfiyn3weRAC78EKQE0sAqTsFdkt0rBuzr9lwGiZNdKNh0AZhZlw3k7z5igL
2szUZ8P6W7BFiKB+H7kXwj+Solg7rryV/5HYIuClG9/HgDIzezaL1H5Kkf5CkmOpE/zR7sKQpO2N
Bc8quvJlOgKC2t2hXxKFtTsxK68g2nuNb8ZziD8l/6QtiClrOpP89c+BO7AGBm2fDICCRACRfzcx
9o9zg4he9P7sQw9Fmn5dytsXDatmkXhWC/V2+7yqtQzdYXIdRypqjfeSMRN3UD8/BcFnCtPfcDOh
GmTnpHglH+yjo+31Lql9NFRtWnrHsxvx10p9lYYJYykpqoYxXzdT4Js7UMtVfVso9hzkDxWTutsM
+vGI49ZmZnHAuRRFJbGaK1yu7ImDU1OgZRfElhJNL8c00o3/mLIG1baL4NzNMrqF2rDrHRSXq35d
k33bvfNet438WbK/1VSSSR8Cii+pbRt/jkEHlnr35u08AbwyrZdxRldNQqRoroMV28Q86MnDs6Ze
Sl7yQryS0/YH80YSxdMfD08anf1XRPc/Ovjh6RKhbye7Ywv5qOI+n2EQ95WfRVkWJ4BnikZQD/gf
Bdqo7D4mWQePQKorqsmR10cHpswZtOKhaU1BZBWDrp2a6L/zrI7kKtg4Ni9NoZlQmoVU9u4KMJFi
bRE20mgK+c+eJPG+qdcrNmkQwQY/7gHIUxnK8XYeaqrXXrt2xRGF0x8aCHHcLWIBkSme2LdrdMw6
Al0eHfUTKT8YTGGwru/jdx9k6BTq795+fv94K9qM+7ds5FPYigI7e2yNlgJYM/bO2r1GFoBG6L+Z
uE8wsgoTQbhmYww0n/UgpVdiyJstJIUVve5XhIetTdi3r/TE8FQInAEZQmAv7+HmwrcPFNGL7O4Q
SLdUuC6kBCEa0lGOhQhqPHvfeB3Gg/kqOlNE12rqmPXr5xRkUdYN4Eui/s9qiqajuVDWG+UclmgQ
uCTrGfDUgizhy9mH8TyD4RhOdAHj1ij/gcLNEsxEe+mDFy+ZORk/j14SlZjtc5PyApRGju4qfDbP
1JF7Cm3PNQmtJBnIcVKGyd/H/OZntfk5BNKnb0uXFFt4W/1KO1jvoDNeSpAR6lw7VcdNPm8qARjb
qr7wCQoMtpm4FSW2a/uUMQAAku0SRH55nP0ZA9g8AskuHKvJzkz5tYNAjGzBoW6nTo5KIjRcrcv5
QiwxU0nPrZ7MIM799dIaQQ+yb4odx9DxZvj9EJGNtrlyeYxagbrWkKGfJkuW67B84xHpdx91QC7k
Xm0tn78zyCjUun9NhZCi1dWLDP/HmXxv7oeUrCyaMXOJ/ayCF8ldY1Q7cGECl3eu2FSJpquqTy+F
bg7XBahVrqeGlughThFbxrvKgQ/EQCUnFdsvBS10HWKy877rS+mXi1WhvzcTjfjKha6cXuCRyIDv
/o2GXCRsTnrf/a6uGrtygC6gci26gn0U6bE619awkX7M82gdfwwkx/mdxzhcy1aoMokV1aiiM4Ot
FTrtICoLizoF+IYc0g3XQqZTWNwxo1H8zu+UMCYqLt0yQm+xP0Q5l/4Bx4WCRmClH22VUVnfBzBC
7yO6N+BdjsEO/ty8OcMwVPJWNgCEBrUJoX/qnRUb/LIzlxcmR9xQDdwXWutqIe+vizlN5H70sXSh
rzkh7XB4k9MU5POSVyEgytule8ySQfNXvX2lmrBiDR7e5Y9hC2xued9AkTOQYtbhC08VAlwrL1jB
heXK/RBheVeMv7845HEo2Kv2DYcJGXWcZVJUaP6HIRQboTUckufbwgYjWz3lkuOwjUJ2+g6aUTzY
dfMVvBlxg6jtvxQ+jLjXrkgBKwCrn31UyRCEuKkl472th4yjZRFUtvpDQKu03RzTp1TST/p9DO5+
h2bPN4zYJPWcI+5WxTXZpIiAHC4cJrAzLHhPV4UtwbOlVOKvoY+aQCavbmodxKwRN+xGt4nYIfAB
OwyfHZ1mZ+8QFmK2u79AnzrH263fkqzHkBaREC3+NxCLrjd/qnPE1eZdsItQ9uQEpR9ceDIeepjd
4JBfZ3BYV4ZLclJtwOg834mtG4TrzMOEJt0KhJp0/fjGRLRt+oEhqM6M/NeKojlWliyn3ZYlGpR7
Xq4m1MqK2iHby2HjOZoCNu/+Q1DhR7aj4mbMfZq4F9GTeTfcwnnetaY+Li402whp1DW61oX1aL7w
z/0QFyVmSENs0na3XzmLHCcgg5UVLlriZWQ+88R6DCi1u7lDzBAzCwHTmtlJG5dpgbATIAsjlDHN
TmibiAYy7ps+TwqXp9ZQ/WnIRultFwRs/zsJtvBYnNa6REZMzrqXIxF6dh850uqOZ5Tx5Lj0vPTI
QB8/nSL4ghakykYghxS/09GEDlGR02dW6z3vjd95J93WtQACFSqb/NPaw5Fz0+3xsviPGzQU8GgF
b0YQH9G/xDBd/L8BiLZVHbiRaM4OIFw0wFyB9JEFdaSLrMRGdTsKe+1WrwIbg17ePt/EumuBm+D+
zgcwBKPhc9haE3zmw4TVSayH0AKvB5LV6rkrRE2tuWBri8qjJx9BHzJHeq3wCA0ira0ZD+CUXjPy
Sbe2IrthwTrzosWQMqj7B5HXSiSjlwCz32wiZG+nH34eWF/9rGFydDZCTedddLK+tbshxRgedelA
2nNu5kzarD9+fhOIbh71kL2kvpQhs5v2KV7r/9t3YoFov5czsRO6I5iBeo6vOybaXXRatp2mm3aJ
jv4jGASyCSK8UVJqABgYs44QDNfEdwkgTW2ymx+LH90Lb25fXFMmIhtSPu1ddbaPxkxYTTGswGXr
30a5acWW8QOJE7B8nHEpkaQDpfI4KESuZBATDoe3GulOy3mCq8NnXPCSv7uSTFLz3CwGNEX/tQ/T
NZrQDJQFn9FZBpVQzB+0gDJGuE/ZuGTOzfaDVAYjb24r5MdMqRWE1iXKj4LifaU8Dp97ay8hyAcz
nmjL1zZfXVWriIoG8wXDbRQEWljCOIWLfDV1SpQ0+2y6Mubh3CN8ouTKJjQP63qvdU8KnjsT/bu8
ext1D+efwuX+M+IIoSailzD8O36setOlarCjZ3LS7D+YTVEOrHBSAETRzErvPLK65hl/3fe/2W25
N2ysyH/Q/hGiHYGViCPLNQIa0w26owNlbqevb9DpIevYa9PBT00BJ0lB0AqvnKpoFTJwaS/9oBl8
OYom0jb7YdRBjbKL1db1/t8tZJG64oBfER2NstfSEwv5TFVrrUtlrVK7kd2lgeR6aZFaO+b83F9g
yRimwIwo0qHFlxKzHOTq2yheEyODGqvObhKuhP+SsWqCxv1/78mj0hGnyo4FwXoLM1lka0KndwYi
KUmJNDBhfBxb3njP0UzWl6OgvKIQYKPcRhz/tw+UEpmbHjKOhuAE4uiE2iLnshQqBur3ekGPtnX7
k56wlHNf+XKdl3SB/BSjd4E1JIPNrqLsPEdHq5aqTq/G74MTJGwZy9M4Wb0LY/s59BwMVQyJ00iM
0tudt2RaxfT+iZ/evKD6bH8NV5FH1aphYuWjGsM73dWCw834/3fnXBXUNBhk6DlO8kwkoIbBcihc
aOUVNvnfDg37SkeviuDHq+Q+4wHzaEEOTtieyQ39KTBxqMbtbjWKNg1B5ZtkHuawr/af9bNrKsvg
W/zrXS3aSyY1Uo5Ivrwf7rrOQW32Us3cfcU+GiwdYYdN2o8WxJlu6gyfsuc4hdV512tQZaJZDkCS
Rzg6ckR9/mB5tcjB5wiLw1kLIXQdGSuXP7HnXm4vSimI5hKDeLQRBnIo2/Hzj5gbdLDPx4v5jUue
SSNGRs8ZS+uDZQBup6VPaMj8ts2Vopo1UR5OOkhciyA5R4u1qo/P6z7/tENT6XtoLNtnTFt9hvGk
Zjzo5phIBd7Ztd69gUTroe3wgoeDz7c0VlSo9zwnhZF9SlRAN/fO1fmppP9fGEsuMBC41Prn710t
0bG1+yjFWQyW84+5NaqPzNU8XDCpdttqMwmEmkDVx14fEoZW/dBxNV/vIwzCMagL+2IwXOrM5FMn
5CYHHr5Wfa71e1COnUE4iOQ08DxV8nWcniPNiejOXwsGXzHPhYYcIyVYLXOZwjA8Dj2fcLB10mw8
F6aa4MwuW8b+xmZbxHIth8XJaBaOUUJAPTWGIvmacvnkYPJRYyd5VInv42UF31qmfWy7NMaNb5bI
L/fBTxf74o4NmxcHnW+B3Alvd/M9QSOEWXWm94XBxm3bYmc0Z+9PnPnumFMEhTtOEcAWujlTaddD
psCz/qnbUKcf2yKI/5sUrHj6vIHVLc4g9nZwW0Uwriiu0pAWFQqFWMmUWApzia6RcLAtHzRAnQ6k
t4/genXS82fwI4OqC6kr5N7mYDe/9BxrluATFXzAej19M2b3p5FS8yR6YfRQ21udX1vlm3vBStZF
NnClCGob61J+CsEkwFOYinJ4/qDvuy0GkEeXsWcVJzSMpu8W98BN6RSz9VUveeXMIwzD+xbvbjK+
bmtj4lzY2sxHuJP1KIBEqHMgK8ETUqdZSmVO1/a/gDizUwcTVirqNJHlNpeMIQmSdbXw2Tvs6nV1
VRjKdrR5gd7epUiAEcBQzXNlCZ+afl4PS2yRbn1UU4S8cUxBZ7TqXc6zqTUYAGdKhYiGD4m1NPNg
cF+0J/1FMaVCdNr2GV7Ledjh9WD6wJZETPGZ2gJ65n4Pd0GHyWPPzxK+v5emZZ4/cmbMkJHMxcXn
Q2FknmqOEzPgxT9JBLoJ90UVBvT35T5CAqkLerb7Kk/WoQfrItdQzfr12HtL1bzbvN2JIrL/xXrE
cRQgkiqYJnXrGr5/RjVVnX8dG74VZr2Y/f05uwXjSWau+eDmw7en8Um4S+2L5/1mRx1LRxG5oI+2
Z5H0Shj53lnC5wKqE2SyVfsKzetKGshpGl6U/oOfjk39HLcxyBnhoMu51c3oh6fkM7yx3iff7lFZ
2Q1vyZ5SRaOZnWTgkXj9AQj+E7VDK/NiXWGLReHNeOLs+geLsUYlQOdEIp41zTx02JHs80eFneEJ
SZ7Myu3P8KfNUrSoACJTb0l5pC704EKceu550Vt9kKrJHzgcO5GYQOXicU7zN0hiAW2zHTXXPVG9
85kdvaCG0pdpPKZAeyixs/B8nutI/hYEAD7Ou/RSeRiGy1kd2f3MaQuS0FQRqzmygWx31+Vqx6j3
R5UvxNpY65Ik9Lgf4jZWN53IcKVgwTyX4na5AejzevGhGxe+NZmIJccUEqHdL3YlWKPP97A1szQB
5Oeimh2qm+CmYBu3s7QpnnEUQzVQ9ndbi5XjVdxoaF+CtQ9u2W5weyv5lLCwL/+T/VcPkS0O0ZDN
cd5rNBZsFnqEHKlokJs9QPzZqtXU+CYiXai8mpZgDhaCgFBSWuKW8XGxSW0C78b8f2PuEYgN/3Nd
qSSXsvJ3KmTK6qUuDv83W1wg/pXXPZEQyFHk7b+kaAMH2/ENU244IV1sdwyfyk49EcSWexckbS+9
jUFhF4pzMXgSMTJWbDc9+EhP/W0AqGTAKaNgOVaKd+h6kXorsSmBRwKXpnKE7RnxGN3oWKa5DRlL
eGtXKQre3lIlVohcsQvQxCp53ksagawxRgCgqKrzQ+P/yd81b1PEYFsid9Ju/7IIo3ehlJYPb4uD
80wDs85nIjWP+WEadyxFaMKaMAk0Kw2NEzqHboouPGleSG9zwjm/aCIYsg8JvLq3XoU68X31N8hu
jDoZlq/3UEa5QTVD25tF1WacrG8YuOutQ6SA+2cWU8PU7ean1KuRKfKOgaHr+uS9HpEpM2DgfCKW
gaW7YewpXec2DHiS2TnLymhv5GoEJJOl26Zgjh9r4LS74JnKoHaFhE3hROwKcB9K2UOPGqdhmF7W
GdKnkSAkiHoP140dwKP8tdArG/5GpTBpgDY3okTB1J/plFy+gR3EAcrCO0D4H5VTFppwC9ATJ9qi
dENS1Ibv39ntSaDIJHZTTdpy13gqbCJxv5eGy7cV2zC8mkSQYVbTW76O2sT/bpXws/CtICAO4OHy
xz5/RoA2qsWr7cFAgvaGKA8M6Qb2wByjOBSYDtmhjRzgDdMfprMCNHTu3wJLeIHcIQ6zqkUJotSp
n9PveQc2RmZ63yUz176HizaBE43QryucPrv3dF5loh+S97PRTt4DLpsphBjwME/xIvZMZYULZ5mC
wSeyB4XBcmfnQnSsl22aPfj1b/Iqffr8LutUND9TplL7+rcrBIEmbx+6S8H4w+p+pVC33kbHqMrV
UJoe20rsKUPt9qgYRDaj7QdVYY+0as71IX3Gmrz82MY/lTqkRn+aTiDThn6lD+at4t/ZZZIzQL9Z
c40Q/9Ao94cOZ+pzXb5g2Ai1SxMO/FFOhbbcuJW6ETEAG8qczrVactO6eWh/9PbL7Icxh12fLvdE
SK/niC1ZlG2dmjKpk3wEqKMz/2UrVdBGiqT8WZCsXcNVS5OWciQ0SQLm0DS6PX5R3OKhQ9YyjFYJ
f7G40xDPNzyPfFSjgAQ3EDYn035hls7LJjvNyBXBa7wnhEWfjHUolfG9pJN/aZMhptQjmg7Kw+g8
e7KhxQbqBJJ1YQJBYwXCixvJ6Qc50LnJOXK8lPYx3WDKIBpKavZshXHwcz6ENIkFh4CrMAnVYo9C
KNAT2KUw2DA9OIwZ58SHIQJJc4wymN+526bQo6wJnvsILCy0EY/MCw5M1D2tPEMjjce9RKQwyO6N
mjaF0guurqON7tmE2p1OXe3qGxsTSHpSVwTKHJL7B91ssHmqob3m0PgGbitPwYDW7amAjjAajUU9
tDwzcHHxW6zzmgGAFpF+zngw9ztjLuZDeXP5vmPb7UfUSgM9T80lBsTQ1JjczPZlFxD+hfrZt4SA
WvB8DpqFjAcRjU22p0IsMyE/v4iz11r84mBvAEF8yK5JBT0oD+Dsw9U1yLWpI+SKdbkvDznRUeJ4
5AvYuFrUvJWsKq74IpMRq+4uQ0Q1GbilamMmIPeSVEveDJtNeRlExJnAL4lxuPtrbdB6OLh0T7+3
5QEGVQBQ55Te7eWjQg6StQ0kZNQEytxrgwIhpRgl8m2vfLVXqX1IyTFMHVf7LxIBrj5CrPzeH54g
/wxzm/H6NK6iFocz9XBQX1jc4DDC4wnveJn/s8bIXFfJ8RJeJhj827OPruCiTYb/obqIapmdSDWO
4O/A5/78Ut/jJJbo38401UMFi6RiOhqwj3FJoBdvbTIC7AB2JPZur/GRib5C5c7gh/cztXdzHGfF
f9iYUB2b3Zpx+K/P0/Kq6mubkOkiVnUqZl42RdMpKgiglWDbPzzhHzghqvWa28/hjnYhjiFgH0yq
HFqfcFARnzEDO4klWqIcMqEnqZCV3t7Qrf6DqiQeTNbiIfhKjdlgJUIzLYMFn+i01MJ43kL1GUTI
pkQJCDRpPCC+Z05ptM3yDGQN+tjooh2hNCQTyBKazu5PmGLg2wYdNB6MBW5O8esfWAeQyjK3nUcR
G2Q7Pnj/+8xWQr4CAgotM7P9tQVSfsj+wLKhRlRUODWAjDlEwGlW/tqDg1O2nrg8PO4gh0vv81GV
uEJG1Qmupxbtizo4ZdVfhc3ql9sBZpisCmJuk115cWuaFEucVb8Rn0+gabA7F2uNimwe4hh4hF6x
R3HexHbn5DwdGJHZviOFcM26lbmxLtttM2Bw2RxuiQrNeI1LHZw8jKCTcRBwABcy171kHU1DL22N
62o0XBKRg7pPFWkPHIk1H5Ndgs7kiWZkbH71O+cK6rP1d8k2V19zPUT/WTQCAtIEqeUWOZPE7dNm
QtSJ1fpFssID8nF/V7qRI8N8J62xTxlRIQWLvRRN4luU9Gqg6No5lPuTQQYKz2cTVZw4duHiW+HJ
8FpHV5Iu9H+WikLgxU38jzIcCsSVP37ciWCmuC3jBQtJPdf/Mip2oxlv6PhqIcizzSFGqgCLi9++
FR5LqX8nBjkQVr/wnASAZC7wVUa+3tpNczBRqePYUbwVp7tPv8OWL7S8jsyE6fPx65FFPwOy2akV
wWbMdk/VGqb8Ht49Mc5jx7Vm1LzdiA8tWAVrehpktVkBThQEq/UoXteqZ/EePBJBVghZZBaw63jG
HcwHEeROQF5xPmGSq3y6JztnWSSR3cvcqZjdZvCHMDo7gIK6ITRAJbMEginldclutnDiVFwWS0ht
lPIE5dfD4bFG4Isrkj0uLNMhfxlKuYr/yEudln85FeTSYgTNxlSS2uFdseets52wIrLLUjhFsyYP
pzgYHW8sClXo05LoBImQlpHmAF3iF8RuQzvZw8YiGuEkaItRE5TtDJK1XGQx/jV8KtPO6UUYwoY0
afIMUEfaTUkYtQEDcp+lZN5I57+I7FPg8boYKqe1BSq4PslamwmXMTuzNwCZYuXLfqOyq6/+7FMe
Qvj+N66oaRfsEoaGe0ie3upv3muZxp9shqyy2MTfwfFMiIrYddIB5KLLQRWQJbTpU5KP5V098d+a
Qu1xwUMseAyrBSa6fDU17+pvJqfi3HjZeG7gkODYXGqMtnJ6ODvIgFEmM+zrtJPa8cMDvQbaZJYi
ONbucUCsJAqVpfUP6x0l3cLh+/n62O/uH/u0ITiuWWEz4TTPudhlGV8HfvLV567pdleZ1VnbaVhB
8D5jh6/RGEZ3UaRTED/8ipdZUs0ExHBeOqPO294P0bz6BfUNuC7h0Vuf1lmPir7GYH+UDB3+l9KP
beoTBYa/fP9pP8K9PwWU2oXV4nAl1OId7UAcZk64A+aazYmwEYgYasebkgj4GwFFpEKd1T3ZyC8x
2B01oP7adBBURBVAv56NzBZeEa52XYSavdKv1qBTfIIz4oQUk8IVDux/1jkgWQDnjs86m6imVb6t
JUeJ9AsJcucSVzgaycN1mlPBHdoJ9sjkrNWBiO38B+L+CfA3z87G04KTrEznooRDnGkcqJ3dwVNM
3PDMj9qtWd2wb5IBtsMvEmvRPoKqcss2Qx4F18LSMjGnwckr3LZzHhPiF382aZw8sc0jjx1GIVdt
qlxvukOUfs1dbrzKVuV3t1msGF9RNW/DHqbV3WeexcQjYqMARkLq+dL3oyAXCSzSIB2OQ8PXPZSh
x3hmqTpP9bLR/3UGWEKwaTVv89bXdeOYVkUXrC7+SkGrYgGRWwpDzRh/kmngTeKObD2bINrxr06G
q6kfK/OF5Xcmwz8AFkVfIIhlzXgJa4hH8ietkfQAtpHqhHPjaG/YS3jwsML7AIkxug/cY2xs2MHf
a4ChaZftCv08O71NJ1aIGuTEAtrUSSBa4LlsUTcuj5V/X3R6tILuuQ/TMUb7YIPASxX+Ww2hKUl0
rVHO/zkOt1Nz66TZM9y3x3P8zdHR4YiIf6jDxlWg0unZzu7q4J5ensafM5lfuXxkDQ5vMcDVhds5
08FyavWhrAULI8euSogSevwn7MS/LiOW9EtcKJfvhT4UEWHYpJh3CPQ+Xb9mD+502AnJTUONNQMN
gaei93scv9Ozh4rHtGZYU0dkTMTiyD77Vxjqh0f8VwFaBQ5y5BYVw4AG5hPhF8lZdl16HwXkTDOP
RQchzkyJH6K1sh2K39r91kWfns8QKmPRse7SfISc2r9BIa1gGBYctfptwYO39FJUXHxCrvYfGNRu
QqDKR3heChsimuLpYF7WYWEdu6ZBJrkoxhe8N92T8EOZqU1RkxMuj5Fde24gmiVZVr0j5RNuh6YG
7fdQe2ApXzE/F3jRVk4i2HF6+IzkVETLZAY2L9V7soiRTIq8NM+vK214iArrAlv+9Rg1Gdkm6kUX
OwzJdIbjuNrhO9zcNitVdtj4SmiHUBSoLxexU3U0UkqiucNliByXatvtZEmEqdyteuzNRZ5R70yD
V5L/WeHLSa0dLtIsqOLW3muZuLoUK7OXcb+0/uotJ0HFdqvFUAEdKOAs9A+2CB45y+HltKnyZyC+
PDYntnOuTS9RM6PbABVgoPPzWxqvQ6wCCtUTk8EQrrCtOBKS3J4xL8cFnITa36fee0R4ex3ewnL/
T88QqCnDG3FHy4zfZYZDNETE30t39BcfV4n8dGlTv6/nEjtw91XFcoslN356EToQeW/C3QRWKdnO
gTMHsikNzv9yumgpbvbi3HeHHx4iKzqX99gtSKfAd5ZC3ubgARwn6JZ8PkMmIx+nrT90ljzkMwkm
210/SxguGiNwlNXgNW8uiLGDdu0I6K0zS0QLid75UTtLIOdXZsCCYaV1Lbx8EsKGYzkopZJpQOPk
NQqJY/eh5V6fT+Ldw6m9s6OlfnQTN1JdlKF76RFPcD9cv3kb9gzHoeAD1v1E7H3Q1rQFZmaZN6dY
XTzILtgNNLTrVlpE8hJHrXmaF9xm1STY+K0NhOg4UO0YTFiG0CwDBF2SFuA8rz0e2dtTrEa3absJ
VwMZ0ld9lv1Etzrn/3QD3gBNDU9ZLqmKY2irPNxVk8ZfNqJIYB12lwsuSpV6jdwpOMI62FBNO19m
rZRS/hLGKUshQKgFNuaO+4fNsYdIAyaH+ax6rMfjw1sWKw/9kp6xhLNqODIf2zQHuRuuDkjMUhID
JqOOBPjyziiicVl604IyHO0dIkTn4/i0qYpZYXmtrojRpbAKvNDxOIicRA+3nIkdRuGC1/wduJey
w44i7yjOhqy9LeqcZ8vO/0q8naLaMVBOt2RBePgGVEe9BH1G4yVli34y+aacPImeugVNbxDyZ5vF
J7gf6wa3Pkh6S2+pciYXuxtgroocJ/e4KlJVGouAUsHBwXMH1ctza82+NfLakmQA/s5dBdmCfiEv
YRwPOXwcJJs4iC/gFsVM+mu+PlLI8q1ViwueISmmY7Ylq0eF2pL/mQUmJBW2Xb7ohMfLy9zfzsfD
Xeanf4Quw5oHGeJnMRHrmjwepvtSlbZTysyT5+lq3Vv0D/bCeZAmVBWIdxQ3KQXcQglSZXtY5i7w
5vN+kTth7Yvtyk0i92wtiAC/ifkogYOrXGmlCyqZX4ibmcUCWH/u2qjGbaX8so1Q4nvWnqaljZD5
EpxU5wKIoCqJE5BOZA1SMjwlEGMKji9JlEzrtRrJCXJx1HGINMEN2GnUZkA4ci81tkWqFmGlxJlh
0/IKFAg0+PYgL5N410G1SN4yNEr09gPFuu3HHeSRpm1cT3S29jfZ4URJrhPtirVpvRxxt4OUECKu
gSLEUk28d4KKXWITBRf7kg26XHZLu9YgGIBLBy0vyWO1Vpp8P36BN3SI4IosJ/MTSOABAQKNNTUN
eOwUD0GsnGRSgRiu3bAZqSCC3G633GXiLh6qVawwUYm6mgC1uBikr5N3xHoDtDeNrC2jVGBWPHg1
lSbJu5HQbewpyvo7Rx3DkHhtqlM8bpEmwK4c87vNXatRiTUyRiZXsvw69wozLl5pfKSc+9crf7JQ
61Ck98qjvPRNLTq/8+OEZatGVyuuwtnPHNuW0fzHGJrUqYhD8wBu0QeMBH3c2p74bQY96MQAFp+A
QUn4tl1L9GQW080yjdub4wMIm3giQB4hmGhDB7GW/XshIZr7Zb9x/H+wcQxYb1TsLvuEC1vtB2tX
35oADpsA2JOPBGKtFSztW78s2SV4RNfi7/FtHHsawwwoUc8cTVXe9sH/2HvHuSMXRXkqrR3RYiv+
fslizjQ5LleYgfTy2equs9yrM+24vOKpAmy2qRo6mbu/XV/cHdVai8Ve1hx8u34zAQcgeRvrpE4P
jvOD6i+HhMBHOE2ap00eRI39Wu9xAF2Lka4LAoSjwam2X/uhZUGjmHEe8yIUjQdmGg9Mj44uPlGU
Yaq/sloq1+QNrAH5c4ECXmYwFLat7BM4WfKTIjflEE8nPiwFsxBcAOE46K+p6ZIDljLcWVJpvuTF
RmR+hgIp78IVBLKk54UGFki7e/SAK7Cpl+jJP0G14vJENiJ00p+LgxLB/8XYWGTwZPP7QS85k+E9
JPYaVoODSr7heFP+7YeXFQUF0UnR32yQvKSHpkCZ5LVeqjfLj/s8Btd/8UJm98rx62Tni4vYmu1q
DQm+BYkx8L5W9N17UM1UWG+zqiy89iWikt58dRmn/vud+gVG0GrxJjClRf6ZQESeRCMmJcU9t5mH
TbpGhvqif+YTMyqy0W/PPF34PvxE/2BGzTbRyLWtsySGCZg2vAK3UkH6MIm+/EE+R5LRXCnE/P8l
NYNJOO2wxYCKcFc0HSamIxFvWv8r1LV9IU7VXrXBDg3hyKUJO10ffRaXIJOsqYvGhR6L4XNF6PaX
4weArKimcOFu65q8dguR7TmWTUtuIJG0yUoXtAH3t6gZU0U6xlQwGCtJ+M7PjhWeszd69Ae31zJn
sMufZ3Fjd0hbyHxdhcWyfRZtRDoweWz8tT2jZnYKYaqD+nq0ihPgOd2hGt02KMrHWXZ+7nRq/TBZ
Fx0U95MwVTBF2gvycPnNdczXHoTafFZx4ht8vts14/eHgCCVslbNF1vsSGPKd63gPL/nJBlVbP6w
VwGAycI8WhgnKWYmeqcZnFECC0Go2O07Y9Gmc5goV4YDXvG4wNMjcBaqjtOCdr0zYdrTODYDYdg5
Yazh7252mG8ucP6UC8VDlqtw56innGOK0BeJWLy9No8Cvpx6Gah7Hl8hJW1NhvNmySt4megELVoo
REIyscnQctPgq+ZLBjLAKLQe4YkJV6RPTMeyUcyhozldQy1vgKl2r++WVTSPCdwZaFS6GVnNiJSt
50PPez30qU7naFVn0umgGrPkikeTs68acmlfoGU0w6F+A2+b4ROqMBNErTC3p9gDAlUXXinBe9mm
/6sZtPn81lG8aTrhStbZk4nt72zK7UuvJnAYEq3sab9hVKpkfr2p4OP0BdpthUZTueJ6L4siKd6L
akySP6m86FvPUkXYfZywxIC8YV9xEf9eQwPB0R1QHEriXXb5yESW6Z/kBfMei6X5UOL/JLFPIRFA
w1yZwn0hq5Cu3Y0lTwGQzihQbyXMlfyivbeVcD6ABUcG+cX3fBEsK4673dO4cGC2tcraAC8xIUlH
SC/x1FiprmDzKVlS6xuLy7KH/GuNP8Pe4M00QK5qKddGWRRCYcKwaFvK1y1ueosWR2FQhhojOWsj
Tkkw33SH8BnhJ2+fmm9g7vKJWNqVP0SHUwcgIDIIlaYNzyMRpj/ZyIaQlZls7Jzeh2ooZIk8rBAz
966l6gnb0TT7MD8/l4SmbJZvKlhNejAxeGfCfnEeLR1CTq5q65HO3bNRCJ5ckPwk3yzsrKuxdpFl
t+kR5CPoB4VwVGJDkcyzeL11c0DoEue2LE4pOw53Hkwe8CBj1wAyQUIihwpuXXcfZ61QxwiKQhYd
zkVu2RZ5SDzZLL+2Mbali+cUUfbCpxmhlyjnMfLCSz8WaTZ9L8b7kr4+GtBp1fapc+uDOvj1wRsG
h15HVfDnh8ppbxNfhQwBEtaNvd4aK8Hv2gynv2UEmBZ7WROSwT28N1ykS71GXWFR+tBKHwSoGn9p
WuRpwTc4QQlyc0mQ/oI/mLnvBSGv9F27vci1PzbNhzUFfBV6Jk3YLwUAjws+dkbOQ+4F2/4kFviL
blbQIrlyyHwpAeCh4HUBTHFohPyye14GbZMqOvnmR1q1gCW5cNs4vPrcfqg/NlBmcBJqrmSn2DWf
9faSKYF2I1Xt16sN6xutBzQNSHTEvJYo4k3CaSzCBkxoFh59CJEWHfAQBY3vtJobIHYq3H+goosd
dVCfx0gO4mDUUJrjkeQ86y9RDVxFmu14H/NA7VychKiGpyuNFdtadJd3m+xCGkJDxgHlDabhfS4g
1Qmqxcw/FAJkGL25g3RbRK/5LxUAiTJSqIWRdeVdS2+5C4iL945JHM67ZKkZHJ98Qk49j2r295mn
YrTYYG3UK4m65171TfNRZlgK4cG9fixk7VvmK5MjnHDfqYE2DaXRF0+F15mHU/cdrWcd8bFCJM+I
FP9V1VHDFTu2JE5bLLS0WTm0qHzdNk0y7H4lr/nZB2fP9yhUw7O6v7zYH4yokVYLLXZwaS/U3Dgz
NvjoYAGYB9DryCIICuEjfHP2ipYWr2Dr1THqaiiH2FcLRxd643YIsAZdPYv+KnRtdRQqsxOSD45s
ZH1UiZPacpb7EwejrZ6k5MFH4kMt2UalWxPItmbTkUqKnujuYckVPz4F4E7gGuTyxECk+u/JNeol
ScL915tbnTNLDV47q59GdC1JEroblWJ/GDBjM/0ciKDqEUlwkHnQT05h2lv/MrIFz0PIO8NXOpQ4
6fYcJue/7Nh8kDMDPqwKHXZvpV2vZjnLMILjVPI++0pbuds7gr1UZc2jyCuchp9wNsr8xUHNI95u
CdDnnpbNB0qlQMO6w5IrMo5Q4deDfhKNT72jUrZ7SeWOcjlouHjDKODx/8zbZMKvCXknii6+iDKe
vvik7rVMTtZl/du/55PwmS/RwnrZnKBgpoZJ/XAQN8EHslunOoW2zhnvgA14cxZ7KjnRy8fuNCoU
33TCp2UTYu8I5dUSa7apfMbNjSnKDnWWSHhA0OFwa1s6XA4vS9U3QRqFpStfW/5LHmwPBPIizxuD
9gvlCvSzbVixQvtx4vNOTITQgP6l6mLfy+3NIgtCBn8Mumq87NYMWWCBIrInEa8uvQ3nAtcWRnkO
EYPDcV+fvsaX8KeTJeWylBGpBg8g00QF+rdtKl7VHm0ZbvUE5p6rFmPj0sL9R/Vpira1FQkWIwOb
IwsbI2XbtyfV+oRRw97obaGOjlFX706IB9FIrxFsP2nFe+K0c2bBNFJt9enV5SktZyOQOR3jOOgr
SbImdbHzgV6s7mCj0wlZbpeAkzWDeZ7TTHm+hfA4j+Q6Bqe6ObgqNdCNjcw8OfSl+OxX56lDIowi
k8Y87TVaNHG4ZniocAXH2QrgasnJzejmE87vOnw+jLeaH0gEii74Dvz0N8PRbTy+2Lr2mkYxATZi
vR+aCFuYlxec6OyWyw06x4Mm9e2g+iEkNddOkO8Ef0EUc5zQOaJfgRRH4nfRhguzyLgxM0i7ZT/a
wOycm+FEa6045HHnJY7hVpA3VHcsE4oYCPcJoAVJY8auS+qUU53sURJiVLTsJBSLvvxTGSrvEUaJ
Lx8ZYD13vO6Ob8QZN5Ht/AUveEmOZhbUlXwDs/x6erNmZjSf7sPVdBS2vTdDRmgremetASs/C4cp
sjzmHRg6Zvvu/uai1jt3uiHhlKXrzF7SFQyZourV3yNjIVSgc+r31PzCBm+du53tK8E+jAiwldBy
qw0Ifuyf2DkoqMHwhFyQoU0JbOrB+aD5jqVnukAJa/HcjyviwChK8Xfb9k/VDd1MrrAM17kPUP3a
5n8X/yw+2xdzNOSLYpheJVsLH7YR8MI6fTq/mTQ2CPXmPcUvmFN7FrDgNd7KTBqxn1RE0qVCkMQP
6PObqfEuRvleBdVWyXtZwJUhaDzun83cer5ZAiUeb4VNKy4tW1nzyEY0Y1f8V475dQGJbOseXsB3
LJXVIKWteFvLGAMNrVPW4Ir5zX7sJsd4ok+CnnMXTrFtyYrtiQTC+xe2CH35rBsfoiSfulrmZN5w
ZVTD1oC3pjFCwEmYz/Vb9wQznSfiqyFtD773YKugmKHB91MFJ03dlYjiuH+iDFlstRpUsPtJP+gT
2/T5NIRQA3+60s8HPnIBZImOHT/yLFNlNAxjgWnOoWGuy1T9d+1qLlJzZotgGOBrIkyiY6/da5am
ezPZiSbpQx4cHkc129Ir29oyg1Bc7RV3DZIbs/dquubLCbr5e3iswn2QoWlrO6D+UKEt/fQXuiDL
qMiYycm7ozbTYn5QKV2ibVMO2zKhXNsKPgkqdiyNFDGAeygNjCX6xNxGrrywWOBiCzsII8NDdPx1
tPPEZh+lcuoZLCkIf1USJsAdOmczxPNKiBoEBHBh/69mge+33KF4XhqGNNVzy72OGmieOSZBoDUi
dsqSR9U1ZpF5AHakBasTCpIw3g3IE3s/qeMhvteqYRx6tp1Pw0LIVkBsePhtKR3Lhw3iS9r85YAK
TqCGK8KM4GG6O6Rb7mCe/vFqNawD7Llb0iJaSP7q8itu4x5qBzEou7qc1d0cZCBfh0Ph9kEwhE0f
v8zGo+xeTtnrgJcCHal5g2SLEh2Ra0w33TduHct62zwHNrVL+bBHcKmlkSAYDGJL12sNFR7rWiUc
CITZc0JI4S3iBWw3lA2049cV1iQiLpNqj6s/ZZKcUDYhx2d4BKOygZaK3IRaRZ6KAvUvka/TyTc7
OdWFUVC1HPo7UCCupzPF1k/L1oMbU3kvFWuGvvlMPHfBBlvUjguezrtwGPJjHHgjgHERXbqUvFSq
87dT8ZsFrcd8LLVFT6T8pqWBx6nLPdSTp4sQyst+vy4PbsQsYN0CUxbfCmtTB5tMrrnxoh29jMl9
xRUk2R7FR9a/m//HragZg72jENLtE+GehgHeVTCiFHLO2V1luXLegYfgMqMJW6TNsDryuIQr6Dz9
ImRWm6iAMMwjGhcOa8s+FgqB+cIx7V24iFd7hu/Fe/7w1SrZAme+lQFEdR/YU9CCZ8ZRKmgYWbnD
J+FhJWj7x0Ck4MYeGM3sDMU/3yhplsCu48Ei94pY6qj3wdbEHDspEy4tSQpc7TqLNYJfO02e8FWl
nvxt4gGc4RMToCsbYldFoX3wRfKaMfFhLXLG5LFirVx8h29TQXMjpjurE8UsZTcS/13I8dl+Nv8g
MNYOSFKTKbTYNEVjueEJLhkp/6VjIWtY4Y02je27TmU6vWcR/oFxbtaG71uGJV/aVicrEK3GhZDd
Wm3c2MKpZWs1mIrtDISX28Q7zxEAB7+ncihGjN5XcZo5MBuJ7T+BxI+GwHYKcjm5JQyFVse1YtYV
EYW8aoKDNMr0sAZOXOYhsdfA/QNTqaH6VQgqmkUqWwPofLKzlMfSkdWz1kWzifBPwHzQg7L8uQ6h
iFIqRH7Yyzhrg89nShyKICBXXCWPA686qBkk5d1c7lpLBON4i7vTfYyxRiCnnH5HW/ZMYagWhe47
85mVFUlu4Ol6eV3oq2N8MdOeMBSjblYWMcMhFE1RP+zNoukvt/+oG58dXY8gfl1DGbw7dSx6Zp7l
IMJvTzMQt4XBZ8W/5IHrhrN1KPApyirC+m4+i/Fky0lPirBFjGC13JrRaUcm4romMVLHNe2RAJ/o
I3spmbcnNH9ir2E3mCGkTl8KkvxjLCSSWE0ettnmguF6mSj7OTVZdGeE9/x5psYnH/Z4sTUSB8VI
yWT6i1V1tug0iOOiVcCj+HSilKKTwgqb897U5hbKL2YJG7/PEjLGtD0x02RPtPYS4t2YjKnhQtdW
UdDaPLreLCvD89L736gOfVMKWgyF2lsEgpWZTnzjhfZVE3rAAISYyO4hT+CrlyemhRnYWptroaxc
JsQyxsu9zPbFBKKQBeWZZ+cdSwL/wAc7w2JG2AGTHyIzujMPttQcgEOD613sO4kCd9dCRStXQZlh
wgm3jOxPNTFPNEFCOZvHDAb0tan80cMHXKjEqph9JvSsQ9HEdSoxC7MHv79y0NKfeVlNGENISDv5
zer7mi9InbmcUArVda3Qj5Kmg2fbU0W8azYhAEmdXr9KO6BE2QeNO5X4bvmwaL5MHwW1U0pOIoQE
MdRA8siafrmjjlV0D7sshl+7DLQFL32i+WSyk8NverC+tp90HHfFfjW0IwTfjsd2tpHp5sfu2jaH
QDtC0Am8PPCgopN5LqlsnGg5Kh6jg6h/mbQF2dxfCMBDXZ1FBoAZU87qzdR1pCRaaZZEstosqM7b
4i5zsmA0OovdJauHoUxU64fLZx3ufCoohyRc1p1soqkn8tyNrzbKpqQ/ZDAyaD7cmSj+BBofIuM5
P2Xni7vx9FOJ3dSwDyuz/bxdTbQgSw7YqW17xsi527wE6Ndvsy1clAYLgQe4UuVbTjXpx4nJ4aXS
Q+cT4KAcY+CCAWvo0TCchM6c7uYUCr3mA+a/vjn63LMqDuaKJf01jJNDkl3DZg+KzC4A2gY2VvC4
2bQ6OYcjTQFlHgPQxnSsrS0bv7wzqnmLAj0HLXgNaejfVtewdo9RMEhBUYmvh1uWcPE2nAdEGurQ
xEurykOGnacOT0aAbFDFsHUxGaixJqiEiyH18SuLfzrBWsytiR4CrPQGckhq1gk9BECiPvn8RkZr
h5M53bsOjAA+HQruBrUOseUBMg3ROVMAPkzAqYIbO3s+o99IMiHeWUuc8LczJe2vROmXhBssJNgS
oLhuMiQZDcIOffjmD/qzNI+2XiqW+Y0D0XZdsZIohh4anMMCWHyEqz8qFtI8E9ZMIPd116GnVDV4
LNLNpGqWEqKsr/whDaRGhJ+VK6mtNWJqThNsprElXcUq7Cfxjnqu8eO7nohPjb+t3s4mkHx3xjCo
qu3/x8BSkhGj5nZSQ1drLD2EOYJXVq7m80jGLGr75shMcaGrfAX2fyIBsgekoersnsl0uALfUmEQ
RTLgR2621HKx4LlGmPycYTNQkHPCPV/iDgzU5hjRH2kqjjX/42Ck+1sFZnmk4IRRM9Gi4fqM065C
FfpY2etyIg8V5ErORWgQ/RjEjzwRebHa0W/I/yLXAO0AhPcXz52b0Os2gALRA2xpY7dFD500fkV8
Abr7875r30uHeDhljbPdcHpsaFlttKJdQolJe6YRlHOQhXbdVE8DTE4ulGkc9myzComBNTdJig1W
qgF15CRkA7C69TgggIu0BrQ9g9AvrISRTs4WtFNaqT6iqKRqqJiWK6XzAFbyiOqGP8ytIfvgIIDn
IOV8/bJEqeQReFBl40ilo/FYKQE5SZjR0FyGYtGBiHtH2LhwJkhrCiR/A0zAywgfhFLnXFQz0QI2
CJjtayKb3LIzmsnIK+PKOQU9/ybqeZZk/EQQQV904MRfvhz+jKldSkoHoBGOrZmpsr8vCq7/KNQH
5IfNzVz4/EVDXVrroJyszYL4xVsZ/ydlBJcoUPi7BqksKcdZwqrGXPDqqOxl5UWPRIuNuNpQEYlX
4VffDmBVECOIGceGfbuLAPSaorReBh3bPhDBDvRHGb321VAuZkwHiD20qcOf8dCyQS8BvhijTWXA
7sCraqhhZHQKiYuKqpTlWDX4icpE3vfMEDjwebu96mhtq8newLY0vlmglX/Ba/d7ch3XIAFXel6h
IsEZRCz7YZbGn9eaXKG4HK4YrDv9sB0kx4TUX9vKL85s9CxWt3hUhwrG3HQX53hensTnU4h6+wuS
Zn/YSVKqU+aIqy3JAkgGHy6LciyAkERyqRXthc01ZqpaklU8g6N2hj2FqE0OGgRZ9KOqnInR7RNa
+YEXHwlJRBlLcR+TgLhXH987eHrd5Rm4RQmlUsho7a0Qj4las5eQBSBmiFen2BTT5uMABF7PwqJc
VQlpek/HNMo4tmoafsg6V7LcR9D94OueADxTFqk98hDfjsZPhkNCAdV5iRrZ1LEwN855OoBhc1NR
A5VG7dBPSGwcxE7uYUckSPLd1y1Zz3HLffAUoLjI0dN+QEUyZIta3/29o6y5vvKwQ7YNSTA99hgj
Qa7j6pGq9sP5u3UsfwEWQxoDl34DfyQmilGkgGoYUzA8l33GJGhhvAInqw8WOp4BSyvVOBER9BSK
T8uSsTCR2p15M/g+wNzPX7MIntrd0ffrMIrI4tojsgUgH+qoVtVVSS9IueWSgoR7jd8oM1uUQGfS
Q6C+vO+PbIJ5tlVWOo4gdTAi2GP9BBdnGZDQ0mT4C66mgleVXcMSYmmLiYVDGtvJJWuQ4CpezjGj
blwfu+Xn3dm41jJCMc8EMEEZYEnltbHPjTH72loqmwexMAT2oUXeoQ5068K28UMeONZQBnRZbh8H
3YR3h4cJsHpuaI4689a5hhkqtAmiVqGV3vxr1wUw8t57DtGJ8PgTxwA5B+FM6Uylad5Xc5p4Z2EN
RShWk+oEdDt8iM4/4EkTDdJdYAyHYT1TAQBYwBbGXD8c/bu/d02fVSYcp81fZrLixYVbEGVfb16p
K4mQrznI97fYF8DWvaNmR0L7kLR5Q6loN486/kOwSK2J+PJJNrS9Wt/Z8kWKWO4AqvDdahUZ4fol
ajNbIIVlHg/VQvMNEqfhppiqx79dYdfFiGDFWwjqL0dEMXzwtLpQW5rrooWUtMc8S/lvEBSif1Cp
G9Up/KCFhZhcC/zqkKf6J4gF98xm/6hfPjv4H/INE32uBiGmLVzfQWpfHmmGfdjYEw66ZGK0CM5w
hOhUNah6jjylV6HxkUTAvh8wyKOjzfxp7BjRmlQg0U9xB8tVKYN7K+eswNe08wEwsYLHTk75jm3I
eCKdWVZeQXeHdzlCJtE3FUVYnPbkOFYjAjmc8F8u6S3c35scsG6uzRjPdAoJmt631L16iq3seXvr
OFccRrWAIkXWGZLC97BOx9/A1d3byElBE9N8FwtqVv2UK04WgrGe+9pvd6SFyw3tm2l68jvFdia7
YoQpWCG+M5CPsxLJ8j87Uv7Oo5UxPcjAv7rDYq8dbTQqMcSeEaQ3IyT96N28bYgMbi52/7n5BFON
NmI31NipgCJWccxcYXQJGvDloDSV1fR3Xqp5ztpPsLYWiFr4A0Gzm/V2erZk5Sf3YLo3D2/N3Iy3
Sg9lZ+d+ZsEQ/U/mqcom/+xcf1Qwhv5t8+wySHn3WXKSTOkjzMvKKcP2t8lx0gAifnZ1T1lRppFE
+LKTF4jekOnc87/Oz4RtUG1kapAcfkLb9Bc8EjWlRXtaclnQNXcGWVCy11ou9tISd/VP3serB9q0
fHX0bUfNO2KgygbFmM3To6PZ2O/3QTIMXoUIYLZffbJGCszV+oEfRZ6R4ARipHhC1PCWOxXPHjJK
SvNDzfBT8ZsaMAMm9n6U8n6txW8Fo3Rz7uB7NNoaVDtt3mwsXbbUx9v1GP5w4xLaHCKWE5fASEMg
CTpm7yC9t22tt/g8S6RC7flPmUz6SbpfLxLg/+P9EvqFyb8AQTtb+3s4PaKnMT3LzMu0Q7bG+rI/
/5BgmnenLncQ2K0tzzGoeIQ/FS7FLUHdQlLLQvMghu/oMkzdymldByoYRrubbHiXM90ghcIg8uqt
KQuz/+6igNg6lhOKg9N335J3xjcxKG05yZ4PdWnsbGZhFrxDIlC6J5VdOxJGK8OB5i1Olj4VpeFx
L9pqm+1983/fhpzAW2323zHTShysq1OzYyR0qeK0QDoP4ftoxgURxn31fO3UcrhtEDBX/crSa1rl
+Dk/4eq6ulkalkNVX0T7HF7xXp4sp65MTF/aqr3q5+d4JyZC1/HjDU9v0BK9FbP0qvzN8UJlI1rT
ql8AAIDopCOhq+X2qTNBi3c2t9k/u1p4pYaOCsJr6Dl6VP2pSwx2/5xFEyIrswzAz5tqUR9t4VGM
qe6ANgld2A/wHwZVR4dWvbsTRs2CYY5Yf1++ofqXUqeF9Sa77szOBDMp/6CmcD0Z2LxUokbWo/F2
FOr9kA3sXvbKVnHkMy56mwuEdfXJX1fmxnCGra5TIGZqzVNTei4tddI9ty3r1JCKriX4zOUfsulu
syhcu/QmknE6ME1eu7xPDf8zDgqhW6W52Sv72fGj8xHVFZOiCyknC7+6FM9W3dldyI0ZDPaDkvGk
5WApu4K1ULZ7GYmnKuI4ux2QyI5/J3r9eJlcSBvXMYJB6jIY1851ylZjuGyZyfSQrOjGbOar7NiV
n7TAfUfHrr3kYLLuTsmfoCAxlpdVyVizJghg5ULbksfkfkjAl/FodtYZ9opxth6NC6e0Bte0VCOU
3Useo5pFupwDxZwF/pO8dIlRk8IvfmyCXN/1aDNgJop+ojIeI7dW5CD2DJe58IcUpoxq9hZ+juMK
zb1WHDyHAwYTVZFHP9wEEGK/5+gYVoMkPqTilll3FQQS4Sa/RXb+gz45lbQN5fE6i+Ts6jFYv96M
FohP8t6h/mRE2fVROmaZHftq6MvKsPvgukHHtWNvSFkYtpA4nK518EbI14YLJKSeIqpR0iD/eUiY
xrMfJgUHvUzEqY/k2ExgZbHLdiJI93m455+R6rZE44wij4gUAGgA3u9Hsr7HKh4WZxzqXAYDbslO
QAG1+UYdtJfD2NMyvMSN9pWDshNgLAuZeKYsoqYdjdC2PlGfJFuRG2CUjE3dcSP8IpvgQzDF4ycd
AfLErkr6gU/0P7yM/Cx11lKelvrS+ho+myvZQ7rs8w1Rm1AU7OLRqk7ERFsIfPzmDpwK9Dg9vP2+
dimzkk4NHYAMhD7nP67ZhxyZfO6aoW1MgQl/qPsv7KZ/gia5c7uErOU5wWVeaSBYsiwtTAxmTDt2
cGPIZnMxSaJMIRHqfhO7+Dli7oPdGGKV+PWsy1DwlBSPg0IXRwg3bZA8A2mG2T2+tzsPuDxbotxt
2QfGbVskHScFqVtofxfJ5jpzOnD+czYleGrwVcOr9suKOoF3tdpbGNXoF6GM6Yup2yj06FQPT1Bw
KL/nlSKZytBMlZK7MgXeaOux6BceDFkoh9e0X3rDD7mGXPg1v1dFtciYrQx4Pol63hzhE/v57e6Y
ebO6YV4X/jOG7LGtsFXqF4uaqKw7l9caJVImuijFttN6HGMXJ3gjPXry4XXTSOERJoBieqzumzb6
1tP9GhiDuc4P6oD2uG5ds9w0g/Rz9oHZr/C7f4UIlUqCI+HSwPr/tMwzQDTT1bO8VvA+tqE/Fy5N
fjfZxCd1tFFbrqL9M7Z1d2fsaioQgWMPJTKxe+HqJS5fYEDN0xdMjzl/SjBqUP+w5PEmJGlGDGsx
W0U3TZMn3LkwPmfJdo+WUD11kDg/c58B25AbF9C+p44s3x4LuxDwS3olJ/OIbY11gbUIKLbL2AqS
fj9SPlQUFUYQVIsIGODBRHlnrrAdNWj5iy0PEXmTfEMGfwygUHkWJPIudQtUic4eFqBTlNIBZjzl
9D9OFHqS0k8ytBB2FHAJEOuWiOV3NU+Ndb6ltk8gJ/R0eBduHSq1wI9WT4ifK3hvSPU49f2maKHe
yM1q3nz6JRwhhXKob0uDsW3V1uXBvF2sOGzEHehXy2fW41Fvzym3W7a5Cd5xmtjzg6et8zR6PEAj
5fr7KGpj2wm7oKak6OnaVGecfuj+zD8VvltAX6eQ0NuMeR52Yo/IJ+wLJu10xeDYVfhIRD9Z4Rvq
Nu+Pq/0Vrwr2K/2x7b+/iNHmCERUW/aarAN/XjxCRK0/BYSFa+78To1/THdt2uP0jZzUv0kl/iQf
muzXzuLxRShhYDdXsw2dW1BVEYzJcQ0LI67rJoRyNXsjB9w2ra3dGwuZGFsSC70UPJPE7UlGHg7w
ip1TTswRr7/XUJZwP8X/JInVCYoUbrYWXSdi5gipxsl8sxHtu21wrXN7EB5xFFAUI9nCLJzWK+gZ
HIPCCpLmsZRN2xSuDxH6J6cMebPAB/BDQ1Re9ynMYC9cxjzOlrnQh7/MwY+25LoQizd3OYYCW2v/
ZLkNxbFAGJpi2GdQ7WwLFB9WN0CvmnRWGoSx8NxT0tGFyw1cqZCEwQbz3FCxjQ7KHI0XouQWQTIi
cJlPUt8ev8BSP0l2fKn2Y7czIYZcdGHHu6y6KCH5yf9OBFu0juJC+eJD2AIpnPeKgb+TI2bLwuIZ
tbJHfjp7soEcuTC10NbV8S09cROhd3yPJ198neOsZvC8+Ry5MTkVEYRo5eQQekeH0XWThye/VmS7
vaY7zwOm4NjDvdPT7XZnn+rWT8doQ/B9ifQ7StV9YY0VxSvUsi+Z8fntZEpV0KqgHPkNJ/P6oqy+
gesNRcq68mh7yvSLn9ek5VKRumBhDfA4Lxgg4xO+0rrQMKaOe5bhWAi3lpE7v0GBuQYnCnTUcoin
fe8X20SQn6Uy5h04HU/Beaje8g9KsyoOt8Mgov6hDIeuTuACkEyk18IPBUacLcSOaivc64SIk/zq
xkvsCbTSQqlBarLJyWJ6WK5lYobAtAHaLcs88jY6Ew1KXgN7m6Jo09RWio16cCNI0fo5hN46q14y
tm3AAS0Mk/g38PIlU8+XMcO5aKibR6lKXbo8s3XmdzKzUex2OJWj7AJXJoSJGtMrMkzAjYcFo5oS
urhTG+8y14kxYvP88dR+eI9muD4a7zXLxEREUkyuklFNzVXza4z7Ll4SE/Lr7NJzQWgyILkYSUS7
6OzS0g74BIYi4DjPvBjpJxsrxDP6/tdF6sI5zsLYtNsTaXLpQSX4anemcfpGyz5MS7DU7K/WNCuH
xhJSSoV4KQAbtWHbSawv+X8WIgm31z/CkXZ3QBXFWiPuJnkfOj4/Coy+EPiyEqKI6iG52ccnk3VZ
aqSzqPa7xcZV9VAkHZnlb/0AKe5bGweoiuCJqBrV6gCRbmX0lBfWSw+htII3voZfXIoGSHB8bAyp
EUr/aPcP1mfJsucQY0WNt745AY0Aq89DW1s8v/MbAPVuCKf6XDDJAMTqcS/rs8yMSDiLkTQWdOao
90vMmYZZs9IuFEJOuJp/RZcPvEBmMcQapzOrbUhMrDCFC1hxXh1jveGA+/GLD5BOITL3lYt3zz8b
ejnEl4ZnrM8B9/DxHfjOlgHC9f9dobFSca0G3d/yoX6GMxvlF/Oki3yrmZlFnlW2+FXeIv5dKfBz
A+YMUB2p6wYMn9YaS1/PC0Y2bUV7zC2sRinjsrBSLT+1QJSQ2AiKTh6LTwXqqzgUdUhYVdlgjXEd
TTZ9eieNE83qmUnBIqr1TY8Cv3Zh4tzeNvhr/D/eNSfzBbscxk94ouZxXiwRDld1MofPzslDJcw0
/qEYv8Y2JXWGBHIllG571n+BXZUsu33msTx+ZGuYRTK3LgxZDRvIqQzxxZdcURKR9j58lNmneaae
gvvPiZnrJYBigzOHEO1I0tX5WqbinZOAi0qgyaDUiX8tJcUxwKMW7z4xYgOkL9G3kdhn9CxGu3RX
UfID1TrkphX9c2cDXrkbveX8n2LJ6Dt5m21st0Pkcw716NwOa47A2TANtz4I/Npj4s06ZKj4lNJL
bwJ7FrhuEEwl3O180SAg2t2Ao8jLP3ODiVl76jYSMqBRSAEGkGVT0FA0AJWG15VTHbjbiJtejpRq
Ok9/uaQrz+BRWlJZMW71k1Z7doouQiRltCEy5VcZFoXy3NAacCN9pkGvbYq/eWPq6kckBSlxzL5Y
cONe8AehEvG4QirK7+/3+LoMzBfYktbBPL3F3ltPlFdz++AL1mRF7sTBTw/1WcoccPksjHD1zhMU
X/C7QIkgpkpcuWRD9mpSL8XV6eQpP8IuNUVUtYraP5ZB2qc1DM3cJuQfppSIEBcqIVn6ocW/rPGL
LgeIHH8b9m4Shv0cVaT1KJoxGrHqNMwW26REoxuR7Stav4B1zAVM4DqsfJbO9YMt7fe03Zc8y1ax
cA0a9miowk8QCbgu1NqIi5wkznK73gcqX/wUzshBMLBptQCH2AIzuUXanMN2qiRHV/yIGweu5MRk
F3KeJSpnuKIXEZM6FzdkSo5HrIzMSr+Kk2VeymdM76WCXwoqXN4Nf6fHgWsQ2evjQgym1ycsYLBG
NjX+g/Bg7SALZ4M5eUACb2HKPK00Bny7LE/XLp/Y2i2gutd/xs43SUuBuhFV/RD+2bwyKlcOVkSr
XgM5oLexZ+kFnN5EK7BjczPHSU2t56TIuYBmoPAO9z67rIbMyc6qds/nsF0xyJEJl7ypDdW3p2aI
N+3KvKix44z3mWXff2E1G/FibaSDjvLm+tJZzHrI5WwZiCY5YAqq2DUQ5Jl3hwxVqnCQfgtkjC7M
YaUl13Llu/n2xzQcwlm4iAWBIgNhtIBSYDZ0zPyYcHzZ+1V5UbLD0npZ6iPAvQiCpesxOGzP8kCh
1mTiQdHKKgUo4xDkZsfQDQ24/0A/jB/WdJ4UUuCXKcF0HK51+F9kVfrV2l/fFsSifp7GBrmJqyd1
zi+865hB46+jv2+PR+DoYvInR9t2w5iEMf4S584dqfcaPl9p1ZAZN5RuIkU9WOFFN+BLGdGug5YN
Db5MmWXysFhVec7OPvGGawPH8B7YjjRiu0w3BtAPStvc9XHCezsNtCN1T6N36oX7xo34xiPFhEyt
PgK1TdOue1Ue65EuOsKEJO//88a9uqH7gyxp6/iVhws9dMoDaZILKLrqlTvOYtVzhgqVakRFIcyy
rzjlxHZwWd/stcpNSXweSruO65rJX47kZ7q5DiCNPhskzcmLi1yBjYPdZYiLGsegIjfy382TspmK
2EMnUfeMQDoN4sk9UqCyJ6PFyPMdMYCO4EgpXyuQKaZZubHEI158qY/s0KtC4bQNE0l61bRyIIeL
w8bppc1v1dop7zgJ6bkJdOWnSWYF6JWOWKaBdqZYXPsTFObOq9Ja9wDJnqfUperpteeHZ/IDK8MK
p009GzeVGyVs6mIPGO9bcRk3rULMxNBwY9+JOKmVLgEkKFosMlFCf0y6VeawzZ34IY0M7BRR6JAF
jds6ywVfC6rfVJeUT9V1UbNsQcDTMsFxW05u6ya0MmLvPQXBw43IzG09rJbzlTYY1ZQ0mH6Sg8tH
1WCnpGQcx0nXDn2T/hslzwUKWck3OTZ5IRy5suvXATh4SdpJmYGjz9QGV2bMHJX2DZm5OSnKnemm
qTrW5Y2Z5z6nWzpOqzMIwkpMzMXlMYxiawtizvKup1SXGmSeAa8T0nZWcoyjUrWF01aXQk/WrKYI
DlZfvlLMnYkpldJ8O5pld8kroBB821MRbY8jrfHs8yK2mSgFi5WUicf+5QQtSCVIZqjQVhML1HCA
kWH4RUu5BGV8WOfzfVvax5+xIs+EUjQfwFXtwicfFSIphtmhgpAUiSIPo71UzlAtrVc+BUk8mDQI
pCYOpYQSeFEInU4i5yCJFhpAW0TDSnYhyCUoUK8iCgaaSRyf2254Y8SqpaSp6L0stGe0aZOtiJpx
mBvxPoZCOomr6mpcy+fcJ9wIUM69B10qgGMwwv9iDr5sauUmQHwATOq8eYX+XibqvZpEYEFtjN59
MbVF5obktklbiF6rXcHmiFa2VS1rYOogXT7g4jFsYqO9w1GWnIsnuKmLjuUX/Cfi8OBpqlCug2uv
qWnL+EwnAJHCMrU+D1fFoYg8ffXrptWAkNhEFE0OPbBfxJ2K867J3d8lIYfiKapNy5fwSgmQQp0n
tfevj8hlvTOyAlKlZ20YczXimvrAzfDA8srs4hOwWzny/Nbhc8POA5Kad85OKHX1jXhlSssVZR0n
fIXKS0KQJ8rm6E41u4PG3AXkkDThc75/af0aGX8MOcXvEy98Cs2UCJxCUj3JS1R6VbPPF9UzJ51x
0sdtqMxO14plGRSNIM60nIXLlsvFjA2Dfbl5vswtPk7xUujz+BU3koRK3M50O2eYAaR0nPunWzTR
TyicYUey/35me79467dsGZD5IDGwDH66/t/461Rgjd6XG/X+GryQJtPyWq0WQEZQImaSICt/ZoSH
FoewDgd9Qmnck8HRRs+jheu8TNthx+r/LDYRnzje8DFr/wIgRAeOoFN5zxziY+2oGorYCRNYNGwz
iPFfoaazTDj8RSquIZJdz2tQmSbJsvbeRiiOTKheR4k/LK7KncBKrBGg/lDox4Q4rNFXrOey8ve8
/72uxcKkXBBY5VnrYNslMYFtlkXBhxq9yoEk4KbJ1clLgPaWk103DxRiX4JphcIhNsmaTcHmILYf
2RWQPpluYqt3OsUjseOrAyXTh/CYHmgdss3yc8t6hC74ujR6AGvRG0GJL71+sLOeDvcs3oee0OAY
p8Ibl0e/rGUc9X17NowjaVx3xniIILoLzQMNTPrd6iQ/CUpVPZ08jyV/JSoa6ILMjTuneFmV8i4d
y7JtQWfv5Etw9DRtc3QKKud+j8LTaM+wb+2Vnn9MGUTsalkeGpYGMcwxySKUIYWRuzPNDqOqhNo2
UMwxl1vBC/O3BqI0+9fnv3AJzC2DXGs5bHTiLR7KdhVzAphKHmKW0iCfZmGx9G3MGtha/gYuIpgU
edtkvqTTST1On8Oc52thgKQu5Bsjgfo3D2ARt57+U0hUrbCSu5V+avJdk822W+9eFYyQdM6nk1JP
zGzu3KNQNpU+/nqtzilags2kAV8dILyJbLjE+wpt2uZgSBD6bCh+B71XGR2DnW1DfAF4QgpSXGqw
/zE8arqamZV3o7QT/CTBtVTJbvnOFhyb9cr4jeAxZPpjGKQoovYNG/SuWZrgzCzJokwCYyHeGfTn
CDnc/XceRLapMrwG+ot/P6MHKBIj1QHfELgCpEZk0f8uPKLJOVHEcLMEWguwm/A+3PeYU1f+Oe0a
oq8qBBKgrqrl1atZR+d9m4jeu0TWkBzJ0hPF33pOS806n7YQQS1MFxjSorCFgx/qZfZpzj1IAP6C
diYoVLewTLPa5QF1pEDLPmQ98othGkr/GhnuXeRUlPmHgO4auxmj/ceK8FjgyZVamRPnbSqeLQdj
m+AXrGAJH293asCg9ivio8DJ2jiWI/Dfr+6uUM8GROBvsGVEhhoIaY4rMSE5JfTTqvg8IKH/VaGc
a+foIMCkAvJvFyOK2yNntBZHsYkb8Z52ifvahkNKXAlTFtqhktGakvJz1BP/vOae94Jl6n48aUxR
pnBuhq8ij5X+7VH/JZCIz4Gltbe3HRgFsV8nXcbCmnr14mFziKwKuZi4ebO7TOD59HjprkqNhC7/
rjGd+QCpx6uoOWCsqD6YJyKcFYDwB6H+N+UlmtNucmbQVdDDFhzHmQEFVwTaYPkiCdOBFTWay5zv
wO+lO83M+UK4j7GL7z70tJLrJX4TU2r7CHKWH8Xf2+/5LDX3w0CEQKnB7ou2mlqLrfUlmaCBA94K
5nBkWLyzJYLVpP7RKuRpsXeGJGb68ZsTG5v/LokMMV5MDiqfyv82LX9mMX+MuXrDWTx2h8Kv7ZJx
+ldSNc3aQCHt/44Pb4twKtOG6ggHauubs+JeB1D7GedTN1QRsEy7hKkAUmwSoUWB2XsTUegtmjfU
zgCCQzZDPbmyEKo+R3+FQyxVHcKTOhsovOV/q5yVBFzNRC9CN/DiGbaQxxKeUUe2QdwYezrvKtEG
vXVvhKub3ITi0H1ca3KgpaQsOK/P5/Mi79LYABVdc77H7rEIp/MW2POb74pKQRcysP8yf3UN7ay6
SGRy9xIhOF3zKXizyaWRIfp+2P1h5mXBFNUVh09bTqcPXQv7OmpZX33nXAHBQ50gO7mD2CENqVLg
DERMqKoIxd7kFybbADdRj7HOTT/Ab7KRsCcQfzXErUFpBQsG0+8dkh5mLDZIuP5AFYArX/yeKYgL
BfxODKsXyp0ZtvFOGq+d21mt4PtmDUIv/GkyZ9pbUvPTWG/eQQdPQdL+EvAnCa5csu70LprlsD26
K8m5kZJx4GXZfTIXXAjso5Fe4HAShM4D1Rrj5AmT3RFjpfliC5QrFBQaF/ikCfZYBzJrut4ygY4Q
jgJKh+VNzsTVIQPvlClROlioSU1/NqmYpVeAqpW5L8INQoQJOS5/+69ZE8gvRCAdOde3h3dIpOv3
soLHpiDaS3HWPMLecmmSb4hMVbFpj539+axUsXUgSB9PHmr/5/nkZ+8JOVKtbncFJIGQwH7Ndki2
/vTBqYqobn9+K9LXFnBkjYpI2gjeLz96LO2gUmvmrhbwB6V5+G4z56ZkkT5dMVHDXlA37+AB51rX
qZGHhzWYVxa9duHR70/1J0nu5wWjUrNoclljYyytK01RUaa4KmGVrHgLNUw6oaIIxyzdgTmSbHM3
goKooQSBkNygRBX+qTvrl12mx4liKOpM76dkkQRRPLpKFoix7wN09nxNK+9G4fHCWzjOPtBwzK7i
cBN9cFqkw0c7I0tAUZwM1eCOF9myJVTgzpa/rRlnoAEdCErx8Jcetucoclp9GqxoW+GqBt6Np1o4
/yPwg4KtBQh2GwVIrmkA2OGSckqULn6MDL2kfYTUpkvkRhlDA7JkSBCLAU1eZO3DEKazBUsMcVsL
YTVSJMWQFDXOO7FCekiwlTcUdilhuJPpTyDNX4ty24TUmGXkdMRgE+26QB2EmLf5Dw1y5geVbqLP
9eDEru+wQuQV1uuJn4J0YrUnK+ih7guKkyEgfhZjwy/ewsszb9sPo1epS8m/CyGCJknnIWQ9C/z1
dGDT0CGE28CSHpHEODcMvZLDA+2FUe7ZOh/jxrFfaqxtXt5iuVM52jZ84ic7NEzdpb3bTPv1Vgjs
sBnmyOR9g2nAHHLRZUuyv4qP64GRbQBxG/IAKvcbGMqOQxahx0UihfZU7+okNtSy+Ocp57hZnMLk
45WRjlgvqCVtoQLMFmv7b9eh7vA68BlBSo6RmpUG92xTEkc6gb4caG0vVqCw+CWVawQncczABu25
HrlwicszFnhgc1GW7ahsHErUiU6qbrO6Kf/GVg4iBfKXzo9yZn1DX9y352uHebfS2XpwvHHqAe92
wf8sjM7FNQ+/bkmAgAXRAf90WwLnh7ZsDC6vUOtMpf2z6OvZwWrTVzgUPgb+n4dDMXvvHwt1azlN
L6itl2xpkYDiIeLpQNBA8Uz4zzn7lXjIZ4xm8UYF8KgWkAnhKH3DnU2WxNyEKkchvr9z8yHOJs+Z
8wmn2Q4Fg1G6GjABgXAEfhZWsiYiECdoTrHnA5s4RFB/fVNjRvfl/Wnj4Kt/4y9Vq08FWcp4cQoB
VsvXaRmbghStkuwKOuNvEpiGP2HfsJ+qmyHms8ROmdo73DRLkz2iff11tX0yDrQtnFkj4dUIxUES
Vt90T8ZRMnhndYdIlBAT0StftOf1N2AoWzAJXRrFweBAup09qe4AXPbecHuqdBia1vv6ODC0zDPW
TJScXPoEBnKEz9Ibz0hzE/NmkLl6HewAAVTAfttpAK3agI2W3oZYlomwYsJdfXgX/8MW6xRrAku8
rXoJ4a7q4yqm90SPkJaa1qY47UnuczD2Dw37VrFkm9zut+BZuISZ1ldSgh+sMpHiAbzHmdJ2us/O
FNuPJvCOabF8NIk/7GDdiuDvhCbMURziVaKp09kde9zzTK68F+lLRZFtGgWwBhO7Z1rVFYKb1ZAj
UrGyJ1CJAm45FSOjhKsroy+ldrRZBz8J3LMnpleW/szlWTUXgWs/gShhexTkLEIxt0eOLEmTyvZR
4NYeQx5q7MH+GdTC5XrawLvvJkLE4x9bioCateGqNkCgw+cj05Hedo4UnltUGXLwYEqPtP8NbM6G
5Zr5IR2YvlgzJFVibz3WGBWdLuyDTGPQ2C1ybHgIDFONKc/EMWlUFnxFzIx3PQ+f1mmXeDGHwv7q
rjttR4nv10eWCCHFJu3ZaRMYalRfvRsOUrFqbz8ZKXkEpRPakRwBLI2Rj4Pwdld2/95rmUr+rpKp
d9xkfffmNHUdqQgyKlbsd2UN8YoKnhqQn419tXSCskxbpKX695ucAiZFMaJC4Oz1xozSkd49g9Ur
LD8AqJLZumnQGrS8HgqF6pKtNvZSP80uywKHsL6uoEFcR+tanGUD0z6PeWZAEWP2FOLP+WIHtT1I
huJvj4BRT33GXLgpy5fMa3zFWYo6rp7//tks0UC3AcuC430GS6n4Ja9pabNhq0V7WNj0ZvH89qlc
/cFnML41PVMwSSKEr052lUJWvidNumScLI9AI2ej86QKQB8gyMawkr2pwpOSTS5h79opbjhKFoau
kVb6Yyrc1ZVkVhdF2wNIn7ej2DhRw0v16jNPqqAyFLOkOb+d2D2cSepIwnbJQGGZykmJtABdWlqU
xOFyqqRhgUHcCFxq4xvxiFY9H67mfDyo7/ud1XELMld0mzYNEZ7jdyNi8tMMNbCs8fXpF5en3O2A
mENEet/NBWdh6v6PJXR0TVqESoHtcXkJAQE7WKaRiRCf0D18BAh+j5hAa4QBOvt/TxfUWkc26Zn9
KpLqYc6ic2ehlnSF2Q/19o7gxO6deK7m8KeWDVm+qMb5jDKfAklcp7gEG/GjIQP5SEizTjnY3sri
CfEgCnF2skvM8TC+JJ3dierNBHVEVK6nk38jWqbmtfEAqiF1qy5/Oz1zgCGjzhhybwqxan2vVsNJ
URJbiFJzoD+RiU75ipULT+os1k7XB5pxs1A1Yjml1m8j6cTwS4G19iBKZBMIfMPslUEELAVzjaxq
vhVGuW263FzpEHlPD0rxjZR115qNtZIHMeYfOB4mC6MY6itFtRdy1RrF0kHYj570KaKeZgxl5vT/
7AvXXf61jqDzJRqFXYU6cSoVvnpyuvoqXglQo3eUi44CGZwT5xLdWq/VD28oDIA4dageb9tsw1+T
CMvZEAPNZuBrSAszrLuBx8opztd6J79KpHROJ+vXPTWGSd6dY1RQBgNUh9an2T/TSUYMncMQ7poL
N5tU1+519b+S+G0HVNiguKen75Qcr3bTSLYFH2bHvBCjWL24+lf3rS2ob8IHrUvJRKcbuf9v7Zow
qloWlF6SAradLfUXp1mKYhuM+RgpUwguC/LKz7tCreywZaNFNLwRXbhACmZa7qXkudbS4mOSf7Px
6H89DJsY1t8vAqkGiND8urI7qDuMXv/6BsH/OhJwtLweR/U+XGx/7HJfXmGxImOp3aqfAPR1tFaq
tgAU9dd7Y9pHo1mnoy9yyPF47Kk1qo2uwVflUyG9BjmOJExwX7L4Kp9s+yrvhVHB4O/HhzZFUUBy
mtCWvDbEjPaqGn7qsfLf8bm29oCdES6ppGuw1FfXnxYxwbV5w8ef8NRmLSi4md6FqTNRGdRjVYOb
bk4NkDGK4V0iXbIHtCcABU2bZ0mbLKyEDlfjkNq5A3K9rvTsI/RUyu/AhbXdrzhOyVF++45QBqVn
D7zn2ZOEQwqvCgrzaorbAg91J6xKIo/LVkMv09k637luCM2Em1vXZeK3E0ieNpYn4gDBp598qtle
2NlhzTl8YrahPRWzQs7KFVLCk8qnh6Wgxat40rVmnKx3RmrwgD3fWwratRnDcu+bXubCVRCxXijO
iZzh37KoA7IsAuc4jhUMj5KuVe2Vg3RTup8a4J3aoHaANiuMM6WTCR7rPE25yo3Z6sHjyJq8+IAf
XKji33Snli8lwOcrYscmjp0CHU8W18Wc8GfWkZTqDXA4uORZ/ra0iRWdbU2zKJ0LMihCfecaoyHG
Oq/lbhHxlP8oUvwEcYF+ZowgfQjfRCbnlFWd+E3L/Wm9JIVjQC5wnSK5oeOj4BwoVEPTNvrDEG0E
ERCtxSjT+FUgjWU+jP3CSxKermLCAl8UhXjvUxq2xOo0RAgqN0Tu7NwQvpt61JN5yOclYquH9e9V
btPuMgE5PDi/ohabGX4IMNTPwgjONNdPXnuhO04Z2yjmdKllpHQNx7FliRdoSEdhFfuq1TrNde4h
8TR5tR3jzgbuWeXPtbuqdf5W7wpP/3S/iNE5f3ds9SHGDxlnBeIBubmKkMJB6JyQeOwr9J+nn6a3
6xizX5FnCswKsYxEXXIXPIRjLWyOrdE8npeEbgXv4BvSH9MMgYd2p4laK+ASLKf3jYyKk2OfGUqi
xcA+yiUQDv9lS0X5LXOH+a6gyuNcX5UXzgW6IVYrr+wqjEG2Si3jVi7UaS0//ShC6U0S/Uhd/y0A
KVFZUWcVQGqyKHgfKRW1cmKs8j/bkRgDKncnlRWza6L2BvdvV08t6jM+OmttCNMUfR3EZEHMdAyg
XqgqslcvRX4RrKDjiJcGSv1weNtueobiyDL+F8Vxor+I7K80DBmDfHBzYuquWXg6sXIkCQuyEGn6
lfu4ZMkjukErv7Ds8jRc9ObRycjaGhU5Nu8oF4i9OQhsGbQSyOtOKHzWjYeV6IWTs2Zk4ME42mKV
bWQ3+oJmIM+nhdIRvCb+y39JQAIk3gaFnD2IL8pxKaBF9Yv5VDbKFoEoW+vJvDVf+UQZEPPbCzW0
BCW6vjs/6NukOJ2RFLkpNWnm6W3zIFLTkPr2ds3rMyVg8REvHJelxea5V3KmELXIXZL6NBOFRLEI
x6QLGsAJvC2mdGJmZkYGByBj718nWAsAqPZJ6pTTulTByHnt7ubqC0/G1qqsj+Wpqe8uzWuOdaVb
ziOBpvCc93n594sjhxpb+wLolOXj+BOsfPlUdWumWNxa7c0iGhhA2kjU1fAokvxyPeO9tPX9rCnG
CxljFrigGMkfuLjmVDPtJK2sdktKgWM7PISEMOKjRJ+S2NfY6WAFdGJuzF1dx+HwCPXkWqFDAWgA
FCihjmIuVKx142e73ld2FfDTnlQqzqLUUn9GUeac7uBv6ZywSzyx7oTctECpNC/H+zJEI0HSYouy
tZU7VS8PlzYOCFC0GboHQbHW7JGqUWW67Ekv+WW3VTckTrvjV+bSWkl69AtGeRMU8k94ipbuOjt3
NrgeUxIMKfq1DqeP81stNVzhgja5uT8xfu50WhT6NQegMhYvAS1DeSLfl+6Mz/glhQzR3EcDXD0d
/4HP8agcCfLWcwEPeK/gHl4+Kr60nBwb0p84tAFFTQlzMDJ1o8Q262AhhaUHE02n0VpIIXM0gRpj
6Zb2uXBeNAY+08HYAZaQyD3ogyBWXSuRV65OJP1ycJ2Ujvrk6PQLC3JEl16GZJXPNn83kDnKmqkx
a2Pt1WGNb4vgcq2Cb5F06VwcALKNceMvmj779Ru6fQarxNCloZOJxp46npexPrHcRmeCL2gtkQXO
pw12g0tNRhxEyIsBFKQRBIi4+tWBBA/P5Br4O7z5TI8mwNYsdxVtjgnyxBdboTrif9f8AT+h2xkg
Fx02wPf/FOWq7JJKtZh32PK/I2ePuEjZ84HtyY9X2IBwUV9hUZQEa3GUgOgjhPZKPdSk2EF0xMC5
jcF2eyH+0amCR+VAeZTs5mIPYfw6dMfhH38QbTXIplJlRzwxZSakPAPwyrepbzxUzA4+3wxowlic
JTUY/k3PNx9U9hnEuaputpMxi1u9IFIlzced2BeIiIXUVh23IY2DryoAWTeHbbiMT1c/SF42TDBu
KH+cIuMnGu8VJohaFOzeT3Ffyxs64ULBq3msLuMXZoAeSSf3R46nWwdPGKOIjWzprhPDIQWy/+45
qEvgkX1Y0697qS9GxGIFVDSE7b7mev/46M5lgmERFTOqbv9F6Vgnt3xQHS87cyce0IFxRKPY/poC
d3D/1cLjEnw7mBhSC6I9ZDZjB4m0o2aiSsDMCfTfkw9TzGsWaUHz37Vegk4Z2Z/U82uQBKc+AfbG
eSjyg6tGVlABQnReV4Hzs2sAKmT6HeIErP35JdT/CDGBfPbrwvb1mLQaMzN06mXnsTGhg2DmH6EA
3afSTsg4Mr1v5azYd2eMsqjj+kzhFef8yvYqYbs85zunjpFLBoM2zySmfT63JM1u4oXgImc8ICHy
aI1u9P9ayCPd/aFa4hM9p4//ZmC7MpuUY667c5n1bIq8hsFa6uJ/1Gq5Wh9068U5Yu2zVop2lQ9g
arD+13FsUEuDoNASn5FmsXh1nhxM+Sz10Lac4myqly0NTN2H6BF/aXpfgL1eanQMvzQrLwODdTiw
mxZD58pNt3XkAppDP+tdchfAkCwaIbATwgf5peCUs5ga8tcnp10RajPe+YnnILvo6z6xfBan8gbM
pkVx1krU43yYShLIGvN5FswtWCzrUHOO8AIg6gS14vmRXSRh/FxOI0mVnceNHQ2W8PowckIAzkIb
iJBEBd9KBCb9/69TqtUAEulah7Qa9QAiR489rX8iULpE/YEaJhLzTELdcPsy7HmKSA9qGKNm5kF+
WRFoTsfyWkHRx2n52eFv3suVF6JEIF+y97/ZylUjdrswHXvu1NOZMDhoqNpFGpaZ+9gLBnQ/oJLP
RVzTIAfsop5dQpJ84OUWojxzyC7szw3CXSUCGBkuIWSYPlJY6POQ9VxzWH41+nYrGmccqCtrpDji
/AagXYRuMypQhHGwyYj3l7+pcHLrKRIhOE4gmgpfARbr7kRefLJ0GgtFBHGIyrzcxI7ZpVsyTGkH
7kw66Z7ybrgodMxYVhQVW5vkiTULUCnSGIsCl6gD8k/4DUYhXXk6NoJwsZfkNdbj+bYqtxbtF4sP
gAmffdO4Bleo2JLK0ikwIdap6XZjjwfCXTK5pyPpGEda9VcXDgK7D9jSDUGODpa1FTOnp8HyNfH1
9JAoFh72SB0g6nuSw4fCo1d4YQK/y4A2I8W8roS2GvL3vnxzxJq0Syx3TpfcDDIV3wPYkdNvDATG
sXKylFh1pXaufgacExFppJJhiLdUzXAk9Q0OrWvF428yicCC/Szg+/5YKgJfcPk6BRUjCutUQETq
0m4JXcPDiXq9EMGGAvrG5pvUjyY8ssyTqyewbQrwFahgt4ttWn9BKDMcTIcu1HBlcZeFB69o6+IQ
m38oIHt5nCD8idYkgXH45YKpsB5HjEFrJISFgSoVKExRKs+qehxOtlA4quWvttLKWCQ2Hdu/M1Ai
IBivmgFKKz0LrTHnTzKQ85gEVQQ96fN391XvkagTAdt3QFIgvq42NYvngC99QScRWuhtMSWwIxB1
dRKXihW6CVPhuHOjf7aEcx8UFCzUGOp2pecGLl8zPuUZko/ekkabQzpTbpx9nBbYXUgp/CrTWtH4
4iwEWaqi9OvRqFFt7J4MS0n2MPFTIrY5bX4/8mP0ZKVaVqotRUXCYDFQqGvaF6/5LCHyiW2tl672
ja+4491h32uhfqr65PIOaHOmvK5gNOBcfUSIfioHkEuRNz5WsAJo1n3cm1QP9b1VldMCSdXCviYS
1gxy4EXtjnG/lYOPrqImlDOFr8U5O9Rv9yBqZp2xyrZcRvXlCyp7g7x65KpcwFZ6n6hMzPUSNSFE
bLTnt+FyLjiLVsvY2eM5DIfxT54AellJn93GMzKz8BDvOGg/IRKo2TSi89EXo4R6qgn7pW0RK4or
370/MhVJQBPpYO31neQd/yBu7CVMM+cTe2Sjoq66loNHwaunB/CQ4grhpws1sv7eB2OHtDvb1uHm
9U6EoU7o9awcQDWkcahKZz7GxaHA+7r6ajtvH/ngc1bofXe2/PtSgPgA9zTzFnOUVPS4noouxoHP
GCX4duhVADZcNiOx0WI2VIPMXPcTQsuPb5hbBDtfP0nbKHcebeN+HWF/hEue55ktcGE+pzPij0Wj
rmwznVPG9ZQl+MC4prG7UV+H/ZnlfFkJYBvERAiv2i4kd+Qtp5amLfZ8tUkgApZn7cluWyC+23bu
otMgYiqUtoXHwz70lPTHvjIb5xiaKqbmyBeq9KIrqjdREnGPsigqz5hmck3tFXIb/vWcAEeOpCsv
op+sKxge6HEYX/aq650KyoNvnQe+98CI61BPnJ7+/XJ+jE8medz3s5hXAcRlEXqFIBNWASJb6PqV
B2ya/kJH9GlzE1u95LgJI3eQ+0g0WZ4clnvBqtb8GWFdFsRzvlYxk05Kwkq8Z1lgnaCHzpSje1iZ
MwfaJhBEbzloJ70jtBiqYi1q5/rP2/ffQWgF8x+ybuIW+U7C5dfMeH+cgS0LQF4PKv6HrVaZr6iN
zaybHi1/YBBc6RgQZZrCXY/iPXJhOtWLksCgnieONcJzTh/mJhZPX+qwYwMdX9JVNTvmXhmJopVX
X1JhH4qB8DE7dnxen8mIitlVqDjrGY2dxLUr1y1KawnpFnYaq1AxjwTXbAl1fLoM2LMTMkPjIx20
a7GeOI25Ilu3TRHF2ivP/3ZIxmDD/TC3jrKs0ZaZHLAwvjAo8JSmCnmIwmuBMxqIiFOlyE6qf8be
ZDC8J3XrIVhB8zwD6EsUTGxlCRQyZ7h52XHShvWZY1bW+MjjX93h8q/Oq6V/z2hq5NsRKNWynmbV
tbslCIt9I1b52r2bR8YqpfQOMlOw3DCkjvCO2YblOPn8qipN4YTmQNzyTHVkX7h22ErK4w0vY5yh
6ChleN6r0Y3kPu6b/M8xC3MWy+ztMc8E53N1BYk2e5opwF4R42Quh1XGK5WHnY8e4f3tKcu2D2nN
68KJACdTYR+vZai/uGJmx1s3Tc9UVDtjw/TqTTQ+AKKSltDxfMjdOYuUcJqAdJ40Sg2gJP9kFKgl
S7K5rclynPhWz1IQzQYkjGiw/SI1qFlmbfjQwrvaK3YovzpWLEAZ+cwsRoHQSGMJKrMt+4gfeoLq
JQxcR/mitDp5rStzAsedNqgSs9bO2eJn4Qvgxlq/P+iNCdrDshIr9sVD5yqG+X+FipgCj01bWK+J
xpDYFrwlqXVKkDpUQsx809hX6oMS/oXaBrFTX4fN2ASmylNXFXRgEWwjvnTnKit77X+t2I5L2T/m
OtWSwycUu6BRCetGwGSxG1ew6U9UMs3BxyXXqs1W0hQemXZYTXJULuSWgEEgwM6VXt/vHMpT4+1v
NR24hHBFvaTKdU/NFFyDdzYLlyUE4OaBZsYR+5w1VUCqyxL2SHxfJckgTtk3NiO3QIbVhjgD33T6
xTuPreDtUXs9UHIGh5LW+aLvhH4L4saRewf8e1nQsmjCrZl5kNGzwWnp12RMbuw6g724n+Pz/iWh
Lwz5C8seHS+qUHy9HCGFDteqLBd2HUia04yP6ZTlBKDXIriKwY0YRtOh+3WtbQdHTLdKsvN67lD/
6z/Xhc6aQt1GyJ1D2nZTjl8SpGvjcEB5xFfslT1MLbkIBWqiR2tgl43Hcr6FDBwyPaM6SSZszwJi
2ycwoum1mka1An0LSDEZmwezZhkSG45fwIfC2WeHV6ryo6//OhwWeGZOQA6fS44qtdibBOPLqrCP
79vHOvqhoPVGAufJwa+kpfhc6f0axhfRNSzeqnoiifwPVPR1z/m3NEB4PUjvH0dSKET2q2GHBVNa
uOoeONn6xjRmlg8J1IJ7OhPX2lx0jSfpoVQRTWsycDIE4Ml4dIJLs57Jostq3dJwjBs4UeUv7E+4
iEtxw1Y26XBedAsIodx+GM5gHbENLPn/xZaLn3FR4cLlzfxofXfa2g9jIHalPqzz7f0Z6SEvtf8F
VtIOwJ0DpMY4KzlXKAuYkgIW67Zy9Nzc95ViI+h6DsCgl1c4RMp2y4+UKt2MD/B94mncsgOCtaSA
PjBupLi0RhGX0LRjGIXib+slsHuE+Ya41QGzWVKlMS7d2qrDAdgAd1IPSNDWIShyylU/cICDfHhL
QDivYdjHeK2RmZDQX7duGUCF/9e3Cpfm831ODtJN+jgXBz6iWJ09rSxl+rhqBQcYy7g4gpTWS4Za
XYZA6wSDz2AhuL5iommtKlyViw1Rcc1zBeh96GjVHEvWuBuhub83OpUihnOHMJYAQGIhPr9Pam2C
F4ZxltS0n/TgRGAPXguooj4Em4+jZaLp5+VDBYcppZ7Q620Fk7VINhhEwN7ysQsizvmFBbkPcSjV
himW78RvBCAPC77xcuw9P/rZvDI2O0/0BTFtAMkUMBUN+T7AW3mc+C27aS6GYVkVwBSuE6MUh2mN
hJgOlG+EHsm+KSbOQqDUnr05X4nVGrzOjk+maXRO6nhhk4jymCfM2VTaqJ1c1oLCyiDRGP7Iu/pS
82gI8BEJ0BuRKvXwEm/o9PF5SolwDCUv0M1IN7oGUJBcSb3X6r8rtOubGy0dlTMap/nq0QnpdnOL
g2HPIDMt9eTg1YCOjaDNTG7YstJxQp8G2z7rxYfhe4Q5PiESf0roafpxuNO0vxf+mpWp+gvNNod1
iEg1PJRduKQqwf5lJPcMId7wTCOj0gL9ijBnofDxZyQHqfAHeZWaKvVQwhI1PkT49B7Jvvv5k98s
E2y/o1Wm3DC+XHirFGmxywrbnPU5NLvAK2Ah2/Le1AMGPz3H8PPBXhTd4x7nvlxKOMAOdhNiW2Gx
tiAbb0UxwFrex+dRPhqAmWdfQo/adu62BEYEX+GspJfcQX1Yi7Pl6xcc1QgLR7rDptFA24bqg5wE
F5i2ngIUU47/hPPuccIae0ogl7uS0bB9U/+Ae9NS1BgAtqX6+GHC7V+mhw3bXMRS7tNB4dl7z6ll
GScsPK3B3rTlOxukCKh2XTqYXfIFtMCKlNRv1wOEzhdBpV+SypVlfL3Lx6QCzL2gS3fkeeBcuvyt
23gOUTc5+8hSJNwcZF+0uxRzlC2dGk/t07TnFpvu1qIzv++1FWhpoQPbUbBB0XF8cxie2HwPOjOM
/cSR4aFH/67/Ghngp13lCzhNxKQYncQQVSYN60Sb7k2nXkX2JrIZe8T0wzL93tIzFwNdhnwr8jMD
fAn/4/DkTL6fcWwdnPbp8IFhlmjoRPrdqBxHUly/4VqKXEkLiKVMELsFt49Nm6qBs0SGJYvN7fO4
2E2s+OOL4QWIyAfCUNMSUwBkr1H6hCXl1ZjkkgTO6FS/TTBTxrRzo+mOZckgf0pv/4f2lNg+xdGP
MaZKqCnNVLAkIN6n3vJVSt2KzcGXcNEv6XM3TNwggB6+H88Lw+4YPXohvm8bpQ9Yiy/Vb1C9n+gj
dBrz0YrLqu5zt12Y4JZFp3lZ5t+nkPTp3mwOYuJjWi1UFELiK9Xh89QQcc7sS/ppyoQLFpoYRNBb
nPK3W5ZamZNusnnfhQIRzz3Pppup2C/hM2I9qrRn93DpM3j0dLfuhWyG4PyxZER4FzmxEiU2AhjP
/lahZZ+U+iwZN/DmIhhNw5UFcqDvvRufkDIZaMipRX27vshCNcDu5zBz+V92Q+Ql96kEMyozRPkr
7ky0XJMGCAEtSEwHEk9g29dBy9+sBm253as+5r27EXiJTCa8BuRTmBPwLwt7tZTgY8z8CaKZi438
JBBGqjFhV+ihFea2cwLRhYI1JANrPq6R9VaawMtWZy5wqswz0RkgLE5B+78ZDNQGVpAqMNlx6xE1
/AR86jV5GyYZzZBNrkg58o2hkZmAXsUoHDnG46q14rsuuXJH3PYjGXUCeAItJz1hpubFA46clEvO
Koi9XJrIQm8y06mOu4QfQvJgf332swu31sRT37EIheo0tlDpv3V0qbi/6/u666+sgIZRyGxGz+1+
sJ5MwLHDwaKIsviz5/uDfezI4/GKSjDMIFv6crmY+VtUD0U6SODSavhi5bTeJNhODZgOVRQCk9eH
NgnmF/vlgNUSX4T4PdZ0XiSZmgX0oY1Ev5WU+O2LLeGWCJemZ2urLdOGKavOxLLQM4zQEwlkvXsV
aOO6pFsfBy2y44tdQeyk6pKBCkUFewQgp9nKqayxmEt/Gyw2RCStBh5ItncBoH2M62FMgaesFvHf
3Xxp+GhetwN2duFlWeVtvL7ZzH/D0VBxvUssiXwuU+Pn+gO4M6Copp7kd9ooMHM+RCtodYdAinjR
T45sXOLD1EKVg9XRj2WArLbO8+b8NI8A17Dnp8YIHTp5MEOhW7IWevSEuVpIQnEUn5DiggTQQozC
dnejRNqfLWo0aUi0G2E3PKx5rfKEEc38VFyFP0iiOZY3jSvYvy7v9A5O8ILAsz2yqvsP4O8i+06o
37nNhmUQhUIZd/vkUzcDWUqaD9WccGLwkCvP3WlLtgWGGoIkYHTJRZLleZRORLJRHOrZAxa+6Q2Z
N3ZmOZWPmupWsgPXAkMhZkUGKAp5c1aWjulVN/HHK7KT9F9s/VEP3FUOvGrnY3QV4TVvOrjjDmdJ
afUr6G15af6lbxslyURlcVtWFJDrcNeMRslY4lnNU9vr4cikdN63RQUki/U7bbHamVxUqvraGybk
7TiV6cSq/gOB/UbCjfy1NEbsyHa5j64ULMhMw0JT2zSBn0v1M8fLCQ3p3CLcOmIE8FuK2WV7uW98
NPi/uL4jFxVLBWv3+HdjtlP27WtSk6dWM2/YZ1zIu4s4jVGegDtixn+lK2+gQAfvcSkHttY0Vdgj
2Kk1rh25Dk0wDOKoYJ21xK4a74eANM61lFpz6XFLHmAasFnzyVVr576aEwwR97xaLR+bKbtu8m8W
G6lmcSsGlLu5YMeXkgpFhoyHaqv/XKbcgCB+hpZxtVkVunTbyYBvc47dSdtDwBdqb5wINmAY5qok
UTEf5W0KAfxN3COFTwHHpTe6rHycA0rU6dCANNfQZvdNADEGnU+xT04AVtC+rHFLNt2qSdiRp8pv
P0FYmHXHznEZbraqEZ8o9CINFZYZGaTmcN1nMNrllte+6t4soTL4RcDB1PD6YOUulUHtXYsNPyka
bbM5c+7Ijr/PWij9PaDzHj1KT8OD6i4QtRaaGcgRqTuupde1jkcQIgPYJMYtAt7a9zOBYNXrvNky
iOKcFSPf+yX7EcoYBR2bHUOOAy4rmjm0Y3Tast71j/eo1KBlOrA0vybS7vvr+HAzfSIr6s7MKdZ2
GyKhlLBZIzRlu71pJk9ZPipPSXCHuzk0VnKVdoeD0OLfxoLXehKx0KxV3Ytfpwso8knA3qIzGCg3
Ydcoqn4Z5WLsUlzdMbW+NyCFVJJhqbXBhcorz3osvjWULTjIeyFEJ+5texChAK3ppj/LGKE2cG1t
rA0h8f4MSIvbiyktazX2gIbHB+ToYrQBX1H8nUzgTHcdh2DiFNdZJgHy2EbI+CssJj8aahLFnJVx
JdBnKQGTCPOFCnPGyBMWmEV7AJv7n7NCaS+kmYYk2aFs31bpINZ+Olzhz7L7TCnyNXxjJDYSBZ21
Z50TYi5sIDZcEXGNk0bOgE4NMsCacyiIBjiKx/tWuhQrFmoqix2g0HiUYa02t1FSokBRKIk0RRvv
As4/AX+JeyD5EofKtCtcDOKxCy7dz6328Ux112Rq/xfXNS5PPsgiF+Irr/tCnNJ5QIevNxMBx9pv
sIismIHTn2Q7Wzry7a+aK8vUkx9WHgtBBe9nh2YXYm3rp6qeKoK/6Dk1MHxbtOUz/jEpkDNXnw+e
vRO8yTS2iYckfeV/uEK3ANuRlQtBetdbIxxewaa0fAYG0G121IfIcCXdU8oxSwFAbywWt7Yci/wf
/h/TDGfdPPgk2UkshdiQ/h/JniYNFNGuiQIJ0OLSshbjYMduXhZwj678Nj3T3S9U1JPdtsWVXFAw
qlu6wKFbYpV2dA1o2d1sC2c9ySuxlGU4AmsV0yH1DyNsTm5MQ90ym/OdcZAdClOGt8RlP9DHv8fx
gM9287rvwi5OpWGEu3fPXneoYnJjTCx+lRvWPGXN21bxsk8Jd6YzgpZFD7AW3efuaJF+VZ5UnlF8
gAsi9bxuBT/XdUHQ72JX+Hbagx2jG0DJE9wIcHkR/s29T9q2rgomTaBZ/lW5gJRE+BpBnGoZtOvF
43Z9nOSqcxd9R1f88RqUud6vW6GCQn3irvmPy8GNp93hcctyre1c9WhtUsJWU0FVHuVfulGPhj9X
8xVOt8tm0b/asH/yK7UOnhG7fk/h31yBVI3iZ9UbX3GZ7kVnVcMRcq0V5ifjmK/+rZtyvo3tFaXx
NyIry8rd2iSzPGR70fhzrye6aNtc2NPR63N9Ef53lJ11sCJDx5PJztGILZfuVdpvFNbfTJM80Qe3
39b/aWSOV7/HkOPpwHOaJeXaqTyARvwIuyagmfcfYPCllUssPSLOluJpI+64JG2u8WLD/1pFqqTo
2WN0gUBPXR0QT6JMzVONDzOM0Ev06lNR3UTXMZlnoTEus1yLcjxACvnNUYoe9Q+q2ZMx42Tz5Kd9
YDjUTEZwCpU1cIAQWH7ICHWwAcUfFSebSZwgGVDzhv4W5s/nNFQ7NalfBdWhIRlYsWMDTBmDHi6c
iKprYzBlasCIG4fDZPSZK6Ov1de2Tay0WgHv1VOhk/Udc1Qrf6nqPoFmwW4rtIenAlBC+/JqIi0L
Fy/HxQWRPnLLCUtNgWfMv8m5QexOUqT+mo7fG7FsgKuWecOb0Yx758ClA4/Fw9dp6LAMU/jLLKmG
Oo7klm3Hyv8X1MmraEUTQgI3URX2tehvp2ZVOkLsmXhtkq10fQ4upaN0sJt8BJPOXDj6pEdaHIKL
rdvjWrFkXZ6ZjGU8auGjgxb+nWbr5UGhofO6+hgiXD/oNLEJ97rh1XFJYR42nsYG9S4T+rfhfvjU
iAQiI1V8dX1BMSh/dakv/1GxLht31vkd7s2jIOPdiiR8RjYG1lSQhv4/xE24XXx72HZiP0DfgjeG
ujn4O8aFj/PRmhOQKbbrgulcaZ/jb0Nf2Rp+viJkEUye5Ws87oEJcKJKb3vZdocvCMq54sp75bVT
CJnD15nZ0E7T01rq4UarKFdMqnm3UbBj0IsxnYV8Q8HUuPU4bL9xXbJGFXz777t1x9o3I8wbc7m4
lnG2XyHBAvhyJrVplnxHD+VUFBmksQjkfq1i6zvgE1c1syCQc7ZBasgDvTL0RKiTzBojmMZAOr05
dKfNQEOuDr4m8WbsJcv3VCWe25by1Me5IGz4f7cKBA624T7ApF3eRodVuCF3+4x/+H75ksjt3suH
CARM3tz7yM+HxrkfwBFcyBDTjs4uMPDEcH0da4U0VCXDSfP1bRck1P3371oqpfKM7hd95YCALr50
3qQASrDDQXRG+wpELEUsXEBC+qhuHZ4Gxrsa7xyvwObFRDFltpB1o6tj2jSCcHqFAlCiBzHSHeVq
DEka3rS9E49qeK74afZAolqFmwpHfXPVGD37zoRAyWyxo2yXyezTvHpHXHdz8xZ38Pnk0u0pPaUM
cOB60cnEgYP5SYE3U/fWEtN0lDkfLG8eIOD2X9oq5ZTHi/s7aTy2+usvZBWA/byMNAkcnf+cp5Vv
xVqqXpU92lSuqj5UYoaoxtTGENS4RpTusfdQ0W3OarB/qMtBRMfuXTBR9yGeX/DL7ev2wpceDjCb
nMMSX1he6DVumPGuM8s++CUjan0tfaTTN7ey01LfXdwKjewuES+3nUVFOhPV0BNXq4hpMh5+GAMg
ZbboDpdz/Mf+NxocfZiQqUazmv+Q90YfYTAKQcTDu8r8zF6bESrE7uZDXUMJ97GjAUHDBrfvyGd/
3dGP+sZTDVbmZ0BeJsZMIsp3RDEzgn3hCphnvSLbVTdLBCfTwFaWFIoR9uBZiOwHhRnGMvPEy3k0
fU+rDmlMkGfy1IsOJIeuua6DJFnb0po4zEsYE/4aoUSDYaKtpzOFVUsHiy4DScGV60FgJ+hY8mao
VpiyT1J+vw+yM+pC4MXc2SkK9Y0tW6yi2O2TE6z9W57yhOmu3i1KreNc7ONz03mnspFMuGRkQGHr
rAIJ70MwFWSn6sasPvZqiDZkn1/T0ARsmTSp9I8Z9hcXHvlD7I8X17RHJ+fjqkgV2aBv2QIhViMe
3MHNr+cdIjcVIzfWkK2WtWiLoGRvZ71oncrRmig5LqJGy+TzL90RbmFWnuCx4wWYg36F8Jdsptxm
outQbA93ytHX2iZh7o2gqHZF6evitEMuc8e5Yf673t5Q4EcUe4EzkkkCJcNcKtM3HctZq8qAgz8E
Tf48aMN5s+GDdS83wk0NtZUMfQ7t3SkvVcRkHznuVnM6Lucps5S3RUPghyhAMyZ15+5a847xkReK
P9AIhsq2kAmdA0GNCnLLrsRWu5GAE3Rj231xpIaz6ioZs+cGsszrfMg8KjUgDjtHNVhJnb9gAyal
83W0pba1hG6YY1ExM29addXDNIGCJTaE65ggR3lHFh+Veulu98zXnagXJ7uTN1G5WiWy71XAsw9D
Mz8CC/62FBVxTPoVeHjYqtCC/Bp1JxmDI/l5X/eGMV/8tih+5DuEgj4DXSgS9S2XSOz/62s+93ES
xm2wyxUOWpeWWbpkgUQZA0st3krjVU/gRXh8QK2efFAIYKHVXEQdkrXg8ywi/DNVjgB/+/Qd3ev6
+3VkTkFzvj4LoXK8GMKfX9mFAVB6sidVLcKYSrjysH+QF0nUZXGP03MzFs7vds4PupKp0WkO2JOx
+UC4LJKfiVEFmM8PKZVR+/qk/c0PhVomyfu8koVtmNT2Mkbzu+3Djcbxby1h6vJm+/b398MKrRb/
reKnfqOTOP/e2QKUtJOO0+kqW7hae7i0FINFAO7eVhZ53XzCO0CFUjgB6/GwlJbhKEgeKeW0MrCb
5hiv7CdzAb6M75OjPJazoocQZsksDxRs9LZbLmf2IDlK7ztjWLL/hOuZ5zu2EF5MQn3LIK5RMiQH
uYS72HMMJaJvF7G7KywzqNhoqZbWrlNTHcmhqxerGC0xuWeQn2jvGiAyfhG2WGRpsWBkFBtriO5U
QjJLce24yCvFLNPpqEE4L5R/EuuxmVFEuIUh3A/o3tLdwJ+hu8kXvzZMNYe0sWUnxm3j9APe+YlX
tingCdiLu9c1XDaOU3hUJYUt/GT8/ibj5LDIs/bWBI7bNQzeMdL22Gx/WcD+cToLgYDGoS5OP43J
XuRqsM+qci5XZe/VrmQhAL5yz1whRgdGedz3Akt8lGftWB411XaoU2evKRYvV6RFWUhcq942aLt+
MVNqrtkEQ50VGCPkUvN3VqN55Uq3pWDeevPfAij/sPxli5OIaM/My8vZpCLjH9Jk8mddks1bX2Vd
s6qmxQiIy8vbIyPqE+P/XuU4bTsfHDZHfdHA7tp2QnIR9D3/JvlCZhuLuKxb39ODttslqIQd6QC2
Z+yT1n/aPzTI3Vuje8l/wZW8n0bZZ+1WUWKShSKANue64HKjD3FW1XZ9N0Bet4Egx91dm4eb3iCW
v08bbuJVssHOmJMe7oD3w96x3uDmy5210lM9uR5O671nor/akkxclsr9ddwisLqFAIF3fnzo0Cib
R8kQxlH1I8CNiuNyoUB6wQftotx5oZzxeI6/Fb7S5HUkLU7yjPbX15oVrQ3dinKlFtcKuQvwJ0L/
pLbo9lKDo2FUMzzNhLsJU+EZXwh4/3FVGkJ37nDUhv+e1Dof40oqQgHvLykMEv8PJMJeiEN814or
MJ+ahnHv7XrPpm2/P3qN3RzoRoqeCt5HYz8K5eli4YIcebMZqvgzRz+vEckbFXEmLK4Uw6yLo0mo
y5UY5D6DotjcgKCnYK1OG8VtOS2mf/G742Qo88++Ivd9M6CVZreAFh2VwCq36SdV42tDccpldeUa
pD+dzX9nnnzyOnxRSbKXumYW/NV3O7l1D6U6gwXGuvyKLpvuGMUN4QPWzNHF18mWG0prn+OcZS3R
+jldVHH+rKftujsxFS57outWuggJm+aVNyGStVfj9Tl+uZNwAyu0S242nybLOTdK7saVIAp+OaTN
L7LeKc7iB5u33cg1tceLhq56rfZtYbSs6mvsjUEzhKfQRaiM17wUgo6+4ocSfWbGKg6nNF4Rq8kU
2z9SwjIx+bK/yAl2Vs8aQObyz0JiCenzaP8EeUmPHGX9o5p1/SbDm7OozNB6JgZGQPx83QY5wA+2
Gw/P11qDQuLBHOlBHyAsCnagMuyqmSnPWuXU9EbzNUPhss46s6MRotae27YcqQ5JsNHt0B5nPEis
1iA9pUftWzxY7IqCReRVD+6PogjRBgwx5ksb/UT1yOAJFE6by73eLDDXOMv2NWKE5cQDHgCIpal4
OI81uBlQx/1eeRajyaJ5a0py9j9+X2YFAwPKY+MpzUxcs5t7rLkvnQFaBrLNgvc36rI19xNYl3+e
CO/uX/gPFob+10woS5oYWT2OEzZRomaJZZxpDpdAvCxhF+dS4HPmCr0s2IP+1jF3F5E7pwZPptcE
72cVRd6a0sO7d6dWbdFC1uNZh1t3pk+fHRSaUAfcO0ZMcyvx4WbzT3xN6cPVwi62MtdXwPzFOyM3
/O0SLbXFB4/skD34UeoKuj5fnnaLRRvkim8DQji17mOwsQk4Kfb0LYYtHZce6o1HHiPEWNzLPH1v
L8ew7DdjN3cumPU0+bLUj6DOURmJ66uU9GDnC2pIJ/Ns+98pru6cELlVLlZvLPl6Jd3Te+RmnLn3
GujJJ/gsnyXCyufZ0FdU7RW8ggBu8gS4zEryg12sRDRX5pAw6pETaoRSoAg7RA8CKfORHXQ1RF2x
a8n/sRfjoW0bOtWyxL89lkDpQDZPh4R6iElYnyj7ikbLXPSSaxEb2c2P0Fn5zAbzgh29pCocquCS
nEoaGxEmatHD8wWF7mmXh+UELkFoMVlAowooHwTCvmSvN+XAkQJoAp3fKTi5YWDVEvYO4xyxc5lL
GEt7qJqnau8h/6TK2OWz6Zi4NqYpqqAggYTDiD05I+uwjyfv7yGgklY/EmDgft9j4A8AGbEZ9nyN
H7Uh0TV1kh1HabohKMHyeQ0vrO4HHaj8Ihn3FZSQ+LC7BsGp6FIUZRGdBXpIj7nchvpLQaV7EgV/
sQ/Gw26WZNNiTvRo4dsLVH3sy+jEtR0l5/KxO3uLfi3mnp79TWGeMmfSRVwiQu0w2fjmLk3hTrJS
ZHb80l5U9hAOnmI0RqSU6HhBbAXKewR82FYsQBMWGhw5VQ8+NaFsKzqoeFnBvaB6Ip4iLV4plIyS
BT34WhcwWZg2OKQOPOfF1htgGL6M+UZaWWGzXWfiQ6sf4Kp+PI1KNKaLS2GDz+VCGlUFMIS/mfyF
ZVLh7JoMYAUorqMKUtcPsNT2gMEoFhKnW+wA2jCWE+fBJPUMEVIoOzint0R8ezWg3IBHmP14A8+v
kcB//aOCLbYgZhmi2vCUPivvAWHIVYx2CHICJdJS4UlKc2oZO/zSJGt+ymYTrimDdwUg5iD5WCsv
j8OOO6piQkI77kXyRt1jdNFFtjwXgjgL2E03dAPm3ZJNkMTW9Xmtt0raMj/cjPWX+mdGjluHFTHy
0KrJfP0Y1ldQnw0SHPoHUFrJgVb4Pg2LCikXSKkOFFV4SXHxnY7VSKOPGTwipOM9cM/onh7FM1r6
fa1RIuIdDxAS6ieesgaFG3+ekQx9lTlvB8iQa33HGDKsf/HqXhktCkUQ/ynWQ56CJ5wx96xgsM7o
iluvodfdOaOASqM/z+46ZXuURA4lVVLoEWqgaoJ3XStYscXABQb8g5JSFTbGFBNQNKeOCP583OZF
Ndyh4ib0DQGVpw0J7rF+aFcovXghZjTmJQJOZ0EsgE60mrrndRDry1JY4C4CVwhxWC1plWA3jGKE
Oy9Hmo6OAX0bg4XrLoB2gAf3/ncFQM7iyrOuIC7roRv1HbjDpmOxGO4ffgra5nc29jLD+BKVw/6d
xI3fH83zJ6pXYaFrmPoDbpECgOQ15tpbX6UuHkIy4qDgU5yB4nxHfYWEHbKv6CtxFsVFMtdBBX/S
URO4QQWV4inHLtD7KPc5P4ivB2dQ8JadUEJkz+DC7Ol59gykW3mQhl5weF6aLnQs1cVh7vYHvYYY
FrJYzZxngyBcdZysHoP9VpbRmWsJwE/Ay+lEr9djEDdHEn+wcukuWHfmh+HjjXu3aaH+q1QX17xk
YqU2XGXHa15xNwfpa2Z1MU0ycgdm4FjSMonTlCZnnPHAvF1c0gGQnQbzV5w2bGOg2oodR0HVjL97
nLZEbBXBL3x+EVWlyT3ibAYV+h1bd7i+GGWuc2qLpKWXWHiIG361lN/ermDVRuFilCZRQyuhczrn
tKQFbl1t98+iu0PbSyt0v50Pj2dMWBtRwzL+MptZ4zMsjCZpoojZWkkQ6n4hGN4NqSL8tZFJjp2S
tv6TgY/iLQfloj7mLngsowg3wz+bF3933e59g4TXpQRV+EI/1VwP3KXBRukX20jLMPMxBWfiDczS
k6uPsWnRuW/sHeK4X2Lbx3I6maVCDtNtHzzy+v+T0udYy4S+aZaoHwMp1KFE8l7r+eFDRH3eoZh2
qqB5aoARrUQqVhbvu62C2dVmL6Ik3rafMYvupyRgCFZdeO88zVBVItfghr3KtzRPXaPDFaRKAK+f
hruGt3MaeQCKbGL3WOMLKPZVr90OAjqbx17u/Yz6vGbZyDUPHeF4gAT1l4VPIsGxj6IPXDGF2a5D
Xc0f3ds/okzZHrDcuyKgpPexkcwFJmKl4tLssj9WHnja7jQABZNK9ljj3Xh8zwJZCYVtLIYV6avA
q3+h8fc6EbcudL7CjK5CKkAhbAVBfOjSpAOMh3VMMVq0ONLVEw5aTdHaplKNarZ/H3GLnDBxcygi
xivmDgA316Y1qPev9BlO2RM8GHrpsprwd4u1TfWPfxI4tBXzHs/uwhnBNTbakyd/ckZ61eHw+LXp
DG8fzHfL5X8nIdzERqQ4Gie/sjretP+dFXGhwPz8+fmsincqzKImYxK7yfW9pOzQeIxdzJirXW4F
ezp23pYNzRwj7i7+Ei4nwJN+NnxFfVE8bUIiCGVAs/Lub4Wc5BfLwKftHkhyufHbpEX+lvp1E8DW
vFead8HRQcB8EVidC78heScE1vW2YFTZ9C9gdX+I8k2zJNcGSjbhw7THIORUG5TZ04CUHJhLtvWn
XSggRexC6gxuv1GusCHo01JIMFyR3Ree3t3TR0vc8+gu2K4wSIu31PRuwHvqVy6PHzQOPh1P60Q/
A4mproQ92ey0+cRz2MxO3S2exmXTEJU67/bicNeX0rBuasopkdlX0XKHHlqJPiEMeeYtZHgyrpPj
kxc1QCS96rOG10CkOEbMR3bN4HXWsR6lJBYdijgZVUOlXd0LT5Q9qRxKGb1DBeqT452E01Tpfogv
RwNMjDdjv8bl7cj05Iz9QC671+ZIumXd7qZvZGOijixagzJ0yLkzhV9LXWeWkM+u1jmzzEbTfmgI
tfQ/nUZnhBxK+rCWC3vH69yevn6alBU7TNLQOnPS9K1y06M959IMhUwJQornqfRtL3UVsLr+Al2+
5SitslN2qzRg74Hbv3uGv0Of0r0Y3aKZ07xWOcm2gJ2IA2WIQ7HJPHQdbvzsACRK9aMIfOc+LWre
684dZvxb2CD28T4YMuK3TxRaK3erkP9EvrlGFItYdmSiJZ91yAph80RZgtSjL0F7gpmhnk8LtdCv
t4teCRJKY4Jp9YTRwXN+w49JGoUQKbHBlzEdVXC1eLwSVSLJ9xla9OYfcdWbvy48IM5yKXNQiftC
4HvRA+wNwUub3TH9HcoVmCBO5/7rvOZlAlO+wtjAokHzMXwi+KnvnFh+jQxeqV4XjOeeuU8o4CWc
DQM32zfVPk88RHdjPPfo2mV5HG6OV2QZVdmB8p2mH15cx31bv21Z0+Xytkz7De5RFQGXAvtphO77
GUqndFoqhnblZeP4AMs5BBxc3zNG76NBiBZZtpa1Ay0Yww3xc8yKuheG3x/WRqqdNisTTQntr74H
G7BmyUpbABh0XHlpfFTTVIjxKyuLojY+21RD5e+vqdOafgHN4HudjSg+P//Q4Yn1lgnRqF1f/PA/
LbN6eTygaRf9+31kKENfhxQuYgHwdmabeGvyE9fGD1LxYgKQVakOEy1gwb5PMxaJ9K4zV6AC4u+l
HabrcPoCjgz3d2Q0lC36bOriQIQ+520pxuCuqhIAKrVuAIp/hXmbcsf5yNIAC4cD9p1NQ7/1XG6+
kJ1U5D/dNA5qfkIF6/VxDlKtB/N6bYvFLNpoyKx0AFPBR+OVxwyPm26B+vXEK2NOr4J8PepfSfJ5
2VfUh2mrID3BY6VQfFNVkCCeYIzOfqhm2rR6M37kbPNSsx5KSWgB5T8vX9SZZTgvAU0NPZVORK9W
qWflD+WEyB1HrPPlCE8/YMAk/ef8X9K6tc2HzIe/fcGd0Nq/2wH0Qp1kRXclJBKrwVDdMeJMTkn6
07u5jUl/6esXjC/wEXT9YdiOgEXHwCbMRA9BRXVKAk5YGsOmKqf4KkLJ2VNMjNolmf3/S97/4FJN
0YmHYtTxK2jiBKN/5hWvGGYKoN0vpTxC8QzNwkMAcj6kak8WgSYlX1OIjUBSPxaDBy2s/1Tahb4B
Mrhheo++7s53ziBr7GghIPe7G5+TLsj1nQZ2OhDqtJin6GxMlhE+0Z6a4k99nrVwXTd0J6/LKNxF
9K/mbjSIemrqimUh/S0ZT7nbSN83jLwuReSeVr1Xm9eAxQkiYDEEKqUlfR4Hu8yKDJ8KfLd0v225
RjwWSzxT6IsIhw2O+nhbmguHkD2zgz2Kn9PgLlqDd0PFNYJmnrPhFo3TPBfTRlidtB06NbhWA2nf
pRKfa94x6uiHMc6O3OLS0emMemLRvUA8H6YxjdGhmiO8BIV9lMoT5+YFhzyW19nb3ayd2gLjNAge
VTkA6o/17m2mSY3EwAn+NB8B85SlugMBwTRD+cdyRyPS0KJy1HzbH+9DcVwk9uJBaKuc1kbK7Iem
vFxYgjhxJNHKs/npy+MLgX+2q4cF/K2oRZgOgc12EFF/aaffvY+csa/zjdIlf06QuT87muvs/1Wj
A5YPf7+6k2WNn/5lFXxDZlQUpsnYYWy346c2qAbuVnt8kHpwC82/emLQqv7/b1JC6JTZg3vqpIKZ
Y/lvTZy8cxOIG9D+E3Vbd4iX46Qi+xIFTyXnRZhpjs1HSfSYpMQloMkdQRIvKRB17uZlfW+MfAjz
zxTt3Rq8zu/UrJp8rvrA2m8n7/ecpJYA/Elbfgb1puA4f7sRDzv7WjPH0vofaDZnQJL04dVh7kAg
4tCVI85fmn6940WZkYkGZzm5xd6tC4pA7cU3T0U5vphcVBlz99WDIMZTjeal8CZJrOb5BoOXARQB
7tZxE3/BgxizTH1dOQyxcGtqU2C9ntuj9eZj+PMqYldLuUVAJ85ZfoswXUHxAjMEGOK7t3cwjtil
duXMSdMw76ArjdQ/zSZim23HUntiq4pnCzG14CCouKpR803wZcig7wKrQyn4FQiSwuxFjXozav2O
GdJZjd3GqGHeNkv7dVL3W0HEYMXBCJGwM5Q/4+uWP/UF2OxlnajTiwMzoypTpIsmp1Av6fBlq7Db
dUIrSVp3J2qS4MtEDrgMPTDhoxfED8c8Nrqf9cSjvQRnqur8e32mEUmk9hRdHP5FHDVY8yisPXwa
yrVLASGRdnffRDaSrMFIVwab8g92U6963TQ3CYcSpo589GJk09YLAhtkHwTLMWNMb2+MAockI6r3
FLJAIg/ANrXD9dXHIApV/ZI8gigEL0qSzJ8GrtqaL3iRuOQDjIMAf9VrxgCHt3dvrLxr3YlYcgth
eH2OBV2JRz/dwy/b6gd6vCwf2QulB0fYyOxWAqGbnDOFDTDK4xsf2+k4tO/bZbK+qOhZGP97v0L2
h5rDMkkhzRA81l6OQESWA9LPs3XOfZsx2SyG6f8LRE6Mvpg5nNs9DVB6eR/3doQZwtKUur0vIZb3
4/qKOK956NYskoV/Hst+nupzGpW+BOXVd6nJnvPvIVoWZPc+AU9/Ac9W0z53L1eHaKmR9zOZhRl0
NYwwFjlobMHaov17niLZiFmuQVGBQW0jJyicDQAUVk/tbjchqlWI18KmZV/J1ZSEk0W8aqenqZ+/
+VOnCRidOaqCUd0fsSusQomloKVPjzCBElRzYRjivlbhvv0HVFWjlvpPM0fqJ++8xKZAWfX9ShBL
G5OYgrTKxOQZHu9V0cGv6eiEsMtZEmEF30P2skqUtZmLSw3F6S2au50GcD5EbQYmgh8cAEiTpSXL
m9lWwzGtEyKSyCPsHIIbbsn4vgdSso/2ACyA2wMUKSWse9/r2zK7pqm6jMzcEEaPUSraRpk8QEjJ
V0lQyebrRJ6YPQAOWc16YZOFMCWvV4D3Z6g9OThnMUlt7eUC66tdrQEAKSdcUe46T3RF4LnJqEsv
enQYI3/4QepUEQNAc6RYEBwzk9UkvaJBvxk9JtsSzyLThR7wgZYA2TQOnYqUuywjoNVV7S1ZD4H3
5Tq2hecbphD7bxqpE3TdVPK2iIq+1oPLV8+78tcizW6i7SvDNjvZ1Y2de2JbMAheLCDCq3VOXc97
UJfE0C+gDm3LB3UpVymRiY9V161wXnf5MJndpVSm4TgXhAC193apN7VFeASx4PBHL9+D8bk37TCo
Wpggm+hojFFarD0kujD4zogpbsp/4o6qtmfgdn+zRf1eMxQlsehAR1eGyWz0AHNQ6zrYYq7e8qOx
jCu9R3Q7Wkd/kptSFWngta0DbPjUSKz3ssEph8viBLlXjYpwSl5lJo3Dz4f6Uzsxlnk7LI/qb+Pq
f/4My449QpNIugJY0a5dPjaJ9HXmUe3j9zA1Gglog30TlY5Wnn7h2NLWa+U2TvPmkc2O4mNRVsOQ
SzhKP4J/dUnEIDT7lmyLtrz3K3zjctqQeLIun8YBGvH7pk36Qs0HHRHEATizVzRkvj/9Nfr8BwQx
1En9/3ogvDlBvdD8f8AANPj00Ib/AIw4lqJtGvjQFaoHlPsYqD5J3bmhNebkpU+a2eKcJgesdnQ4
HDxmyjZUvZLqG00Vvj1zVP72/A5KgkYikVwKIjFNQvG3ZjkHN7MtuubZPQxQq5MhCrXkcy70YTIA
W+dQGd19iuCo+Crzq6KlkKTdyrBCi9oCXL1n6aeJD9fHbogTRGf6ciKci85mcUcM02mcJ4Svrlig
Ybb48e0sWARz6Fvy10ZJegdpAPVr7QZTdonHimC2HnulWY+orGfcnOgHMCIjpyPTTwVhhLnTJMda
Voz85rhnpKg0rtjRgLCA0d+z+2QBVsi2WFBX5RjIWpRDZXkSXluacCvIInBFuJi1Lcgia8CQ13bH
0AnWuDYRnUFwFG/48TbysFVxgO1wP61/pDSMDDiZCRAbXEzza3vwxXiAMcZRNKGyFeE8sFhSh/Sw
K/WtA7VVcUaplgm8sf8AK1tIlFJN0wgjQJGDfig7iQk8I5/Z+IKx24qMEJ5UBqAr9RTRP+8eCazw
LGyf5YIgZI1SbyX+ZSJD02h3IQz/j0ejFQuixEeJp+8aiq1PLRv6q21NQjp1f73V5TgYhh5/93v/
fSbl4xnHgTgn5k/fh6RDp+sOuSjE+vX2OtsW7C1N99mYeqHymKauHftTemh6yW+SHPAyeVAQ4ZKp
wHE3gtt2x0omBHww84KkQyKfU8FAPYDLUkhIXp9d8f554l1UoIkzjKOBB9fdpQm2RjjguWluhBSG
20lB6iVYwS6uutRfVRleqMkZNHL8mrxC9Cw9NUnoXeUGLdSvrcHPDktGjF86NNT8GkNShWgtP5K9
fNgb2BAnJ1Fmu/mjcoDzCj87mR3VP4XjELmDo+iWK3/OMdLQcuZ9Mjy8/nsZNzT4sz+Yhq4RoR4P
cdPOD0C8zry7jtarFEHkjrmU0YKus+hT1Y8QUWvYW7JEVzrRZEeLUc5qP9NtjJW1bDlsZmssQU3t
lqGAYIl/PxmJTuixAk7DcNwlEjCdT0HkvzwbxgON2lHFLqphzhXB8YN/sHgtTN0x0dfmqhWgmXoP
lrO83z8zz2L0cSuTVPvWV44t+4017Ja4bRJvzlxLu2p9XU4UfyfN5YfULFapedgud4x5+8bWyxms
NabffTfROSDW2+5MncYe8DLii95vNpIvM+7jmKS1RE1F0uBbcGCMoTXbG+ILsLcp++TcZRJdj7BS
/ZwteuIs5kINikgm9kjgoSxRUsDRI0wvxaN14GcESe7f4gTybtvvUWcGfS7K3J38Wi6c7tYGxGce
qj6IzXBwnWhzauIlHUctqxMuX1Sdb4H1ZhMQYWNvLMN8DlH735T3dY4/jWaJBW9/2hZ2X86g8F4a
i6ElVXiU0hjbEpNwa53TM9ZZ/oHOAn6jafh8ItQdWtLxHzJmj0kGehNS0ngA4W8vslUtW2JQVDt+
dkhPGUYyeFDHpyyVIutE1B2LOPfQNCw8aUN+We3F3K/6jOiPWqGhYQR+ZYYg9Q49zC9+7hBTdD7A
l7V+MAYa2qWfbRFL8dZfLrEVGWJhs7TH1zdVIzpVvhL2zwSN650Ksw2D07jmmazHTJ37kCP6TDXb
WAu2ru/Uj2lBQsLvxnuSZPyfNQMRqc/Ty7jWAX54kBRXW/I5qyJMtQRPRatjZSCs7TpbaZucHDiV
h5lqQ0gVIzxGijm0IUZsm2afeWoib6uXloh2+730na7oEz6s5blikaVOtd/zo6wZOg6Jk5W6lODi
xZNNzWdT0mJrrLomXMeK6hPwfk/BponuYJUSgOyQ1vzfBne3OsSjylJx1+T1rrPXYN0FPn3WDMpS
mPFOYEd3JtWTHEiJyYY9rkDZ8T+XFZUq77FXOK2nsqnOEr41td2sG0RNn2AKs2oKKbTFNGM25EVl
YzhKxqCmvFEU0iHqehRI9wKGLCEIrOJupL7PtW+HqGNNy/K1qTRkMC9MGdcnPgjAYjNaarBCLV33
VwIwKDsfBHgN8CshbIr8L03pBi+eFxCDmePiq7Vcd+sigLpyvOirrhYrRQFy4A9wEr79JjhIvjIL
/Zd77VAFaPh0dB7drXvOAWSvrMp/QU0O+1FTEeqevZ7o4EZbSZd8x2Q2BktilfyTHIbVpUruohfY
O31WZ/uYhwt3yJisxjsXd2kRLxyCakAUP0dtVr+QFLXLRX8JfDQrWAyDXvqpvfTW3DQMQhQ4Xl3I
JI6RcJEgBeuc43QGcawRl8rMIE0WL5bWK668X2eeni0QkObMVv8z8vuQCk7BTCyRPxVLmmCw3mxU
GBLgcAwqCedpEBV69qzWQmKVb0B5/vbIzZIuLeZCiYu/79M49hBAnI8aVKOfEmf84DGX2E2aNoZu
0ZzCNBXivo94CFjh+YAwHKxqkAg6ggCUAdTLKQ4HxzetJntB2HVP+f+wZk0LgHw6j2Y1FLZYGQcz
ZDT2tl57XYR8Hqy+svkzMCstmp+LNmEuJVAOaMfoxHBcqbowUA/A+q4kDghnPAV7UWmdctFlMtCy
ZoIxzUI0kdIIF9il80sJeWpkevfllWYPgXFXzpNGYuUex79N7rQWCETsVZlj4dGW7DIfliT6OTJZ
n1L0ACfSmwX7CxClkXZ7U/Rf9nE5xQZGFKu+sQZSGuUIbMnX6Zt2UacQyRm2AiTFFCap1uU+pDw8
XT4iD1uoGD/SWqg5X1uy0ATA4uRbw4Did9BfFyWXg64aXrbyXDEF/+n7F36gOgCNVNHMkCXvEMxh
GQzxeml2PMGGMZv/W6QoiGhsv9xVRG/IncD+AFxRSOiDIHO4FLFHubPiTFhIqULf/2HmzH/1hudq
Yy0yz+iQ7oVnP6VA+VDFBQTRSlM49haY3kBB9GyV5mFQ46JxfDQFhxTbQLSfu4IYLygIDmuXrrPE
6FpJlSSrb2WwjFg4tLe5T6TnqpwoJJc9Pvvurbh3Nf8+sQno//WH/9W3YUpzBy8bzd7gxJ5w7bE7
u14q8p31qeNwZVV8xdMMmq32FRaIHFh5zt48tnzI3SFmqhM/V9wagH+YWSwauzTKmhjIBeAcNBN0
5h6rXIwWIiZlkUR3qOHS6hBZWvVuRlkyV6Vyc44z6VLHvdG9JNtT8xukt39HSD30o26rJeexD8Mw
Y88DJZ9JkbPdaUkAQ4ZcLNAo5MNEVNqrCgFUYidXK1mRv3J3M1SlIv5fpPsjfh4RV2OQkG2LIlC+
KDXpQMpZ/wXc6LO7pb82v9JxRNdwWBRVVWScIdB16YWkJT4Hz0a2Vx/xq/F190p63Q5J+H3Pmpzl
YgM1mveTibkvvHW6gUZ7YNjtCWXfAsG0Ponv0IueoDBNVNqpcog38nDwxz9LTT9pXqA/PzR/Fyq0
ww93Cu3zYwhsqEXDh4JkQfKUaGhjaKlrtUfRwFLeAneO1gW6t/eV3JmcPxrCSIsAeZm+0GUUWLUB
jnyYreFpBnMFwECzsbOzNOxie1pV+UbIDHScX47rhWMyIC4QVT1Tu5jyF/udCu5TvaZV9T4L7ZC1
oJ+ghyKO7e04OzmXu9HGcp6Qy0wI2ZIG4ksdkceakubvmv6AfDRlXxgJx2CIfJA59RShvJyFbjkB
E4gwbnau6coV2981N/Kcb9kUPki4t+d33hTEH3gp3kkvMV3Fk1tY7Y6/CqDe+HCRJaJGeUmsfap9
Fy3uT3z/P/HXF3o0HpjSfh2EmLWfgNgCW3iZT/LeUXilD5wqkiuW88mjsoa1UX7qT5Fmpb9Yxcrw
ATOIV9bcKr/oPcQS8/pCGRb8262JejC6bT21c0Cy07ymVkYcXUk0hi/jBVckhSyQGtzditQHfqG7
pgFTiMhPmAQoo7cWYq8OATl/QT/bmfNgmE8TV4b6UeuJa80mAex66gu6OJ2jJKqB6yTRkUp/IoUt
c8zDPgAJEkULZjxJ2tMixJPMiFZWNQ1J8kB5OripAQHXuNusaTxakhgHB0Gdu+Ho+BW3BoIZXq/a
NG+BLcoedpG4IFSbI65gTr4aNPb+9AUvm5227Gw09sPoaczYzmHomj3OSBSFGUjWXvMKJC3k7lxh
d9I6oN2WzXGtaVXpkFW6rKUtCKaLsEuUZEy22pNhzNIwqdaZq/9jmRiVZcVwv8AvYk7rIbclXVcm
z5a2DZFIOyH96B/QcjXKQPkeMLV9HQMNF7j69GmIkhYhRgZF/3orTjDuyf9olYySjvRoNWbzeBo+
SWOFeTDgXJLKfpFtxTgNI9LFnYz6EBSG2OryfjQq8qnG/T4wIvzBdqUZpQ0n6ISRm8yQ0PyBva14
3iABk/Hsr2tePMBgyY1N8K4netxQFdvC2Kfc4ucy4NxYkrrNjP61qliPQSnmVV13dq/RuT5TzbuS
bQ2+iUkwqi+deY8VMwR6CxuEAaAttp5LTzpwPvehOfMPdV2VqFOIlsbQJKxPfVrc+qmKHZjOekqd
aGIjlcWhLuIDIJQX0E0GhHRuH+FvoWcsqgH1hUNydZ1UhXMT4p66OcZahTHPJzNlz1n22wz/JHJ3
9sz+UFBqD3A+NmWjyfPmpfOEt0EXJriCfi/WE5l2oF6VxFsl7IBiFL5KIsqdh86IZClEHTNdvgEy
+fG+W/BkPpvmUF5G3hCOSTFU6w4BSEgKoME5a8yBbfkT+lqC25Wmtgkqpq0IvxuJnhIm7QhTw9P1
9T/RmPPxVrF431OBKHL6VgfwjJUSRmeIRPmgcLHmwJxKHNqlmbPVlMIC+FwfuHn7NNreRVsm7LbG
AUwwQP6biMZ7A0LOrH5p2gWKNZON95HwkUhc4WRNykBDcGHLKo4c20rYE0KWxYkhgueXi/6Thflp
YmsItD6tCegticcFTZg4VcjFyaYsk8vhuPw1wvnhm5hiiWA1tmKoa8C6kv1wsK57n/CkaBfH4OF+
Bnk4MzG6qfm0w74WuuTprLEExvhC0sPHIgW4C742aHnPv0kwEEIZS3plIa1LKvyq28pf02UbvUeE
6R6CalnRyCvSwtdFPtzqTQRtxme1jywwEhSohLiZ2QlGs2BWZmopLDK69JxcuQ+Iv1dTjh6EI2Wv
rcGq0yX7snWTHAgKoJAZpNja0uM7Du+DcJIPX9bPYSgIRbIQnrS4smNp4gubGPzdY+6/x/03jyOs
EtWoTSP2JP0GmtR31L6NRr6dFtUVjiVVspPP5IgIK8RXK44Vz/Xl0ByOqCKXbvW+A2Qmv1CWm5ns
riBQI7FsDy2lVmGc0Wtdu9kouSPXIdysBt+wCuYQhLCHju7tTL7HSsLqHvRlcgN36+Kne7S92uao
UuD9lBGFtBpo5xTHu25tERqVJqySydoUKk9ryHpG43rhS/fk0Jvc5Yq7IFK8rrjBUHLJnPzCe5Hz
ZKZr/Ck+nUJW2xeo1pvXy/z/3MVpHCpc5fIEcnqN1Ab6dxEGN8p/Ygxf14kfHqqBW6f1kj46WPA4
I6WUHgzX028Hefa1tNqLrSzlOoP8SRkcmEyu8XNyLE2fAAlgDYodOn8aTF2N4bn5oi4HI3qvV3AT
HA7UYzlIEF4XNFYkSsPTjiWh65asqSMew2Y3P8KRMRaI4ThgRO7fkhTcrEtovhQmii5UNIrpBMOQ
sBySVJuNQUx2HtzirwynoHN8zTt3VJchVhkuJ2cHiDovps9VdSjzSgRi05OxyslZFIVUlJ8aRVqJ
oeDZsfz+cNPAGiyi43nIJsk3cWMhnLc470k8NzaDt2m7v1ngBiLkzRH4aAP8VuOtwDjIr30pch5S
XFx12z8FpC0lJ3mmAU/NzjkhnJt5lYE2OlVKqgIujNELbzeEoD1BWnRShckeD2x+0jtMQu6OEnii
boTgKlQA/RqaK+qhjhrBTeQ6bEuiEuOrr+ewU1jriAWEz/zW4L/baHr75RA4aUys3BfGP1y5JoVg
UFNgJ9tujYEWEzqtNJoUbqvLVf7edHcZsxka1+k8J1S67Yh5wWB+ZQ8JvpOVQKwjTrOJ8F5TAEfE
MpkJHkz/gyceojlm+MdosJrzY3XAs3RONXM8nvcH49VcLaCzGTyEgXJzYQC08qA6ehhFn0nu8EHX
dOeDx1Pn3R+1Vcp2fDsDAwocIXwy27yLwyGiTYL77M3KJrrRhB1DSKGj23bQ2QCdcE++e7dsQolT
dYzLv7zBlzP7GpNOjH0yWxhhvY5b2o34qFr7U8QOM5ckMzmZATL32TyGgOADyZqeD+8ZJG2+m4qF
7TDROw/cTVyBe3CTX1CVpTn4ZG8nbXntuA+hCVOEhFcrJCndiYBGvjYOFuz3BCoUgK51dds9wQ6p
z+Im84eLMOsTLEMZO8l98KOmOusUS2N8a6loFxEEyYmqP/s0yu1r/Zb3BCKF6z3G8hObwMWO1OAM
wX20DOl2cf6OJfh8G00rd7KSvxDS34q11nZ54q3DvjXNjqY0QLdKEEGJP1SlFsxTzThLyoMG75ES
6INNbbUbdgSevOcFBgOzlPSDTR1mvDJefreJ/rpNwPhmrCbT4m7slI1fSjOQ8qzBrMvAUKiHOQK2
0OJl+wJHBwCLA9saNFMjU+tb8eQ+KtTXdfX4oVl7Kc3WGsNhJHDP4fnAqKLISzvzQRZP5vUQfoDn
7+WICKtuAv3wuZhhRTF9WC1lKrEmFiqH6pLl5ErKdPIhRbd1fzycn5bfNe4jcH2OkeId1v1GhHzN
SVw0XSGtrkoOBhF8DKHcUX19HeeojGtSjMNBwP2SSXr8/6U1/6I9sa2kp1zgHlEDM72lEtQF0Qku
md8KhmigKuVR+vIgXDUqxuDW4fBbT4x6CNDoym4w6ROCv6S+0dFLKehCKEus9gDnXLUdAYcHbRTW
PmeQI5mfYZXFGwBV6TXrtzLrl7S9hChojV/aMiYXVdIcG6QRVHczUwgPD9b9ZAZQlLeMEpkiV7/I
oFYjOs/oVgckasxpA9SzYP3OQGeumkXwRj3q0AULajyoIeMc0vZqVVgJtrkjHHQJm7r3XWbgq0RR
dUHjSNKtf/HDcZJVGpiv63hlg89H2JUbUx+XZmhBTZgz9A4UKZ9YS1zfvO7Q8hnk7Hzcnhpg/y/d
lfCAjvCaY6v240dItwFGR4apIz5iAb92P/zKmR5nczKi8dbdSbb/j2HTo9Rub9gS3qOVgt0EMCLw
Yy70V8ySE5RL607nXtgGXEJ+QbuuvHyl2n+JZo2/mVxj78wC1qz8IxM6Fp3k0xk5PV7aLfUK/R5I
Eds0Nr6J5+++TKtuBanIb6oWkeRpMevytopwC0le6XOD/iVFR1HO1ougj/qu94RBySycR3VadC/3
8jABxoHrh8JYCYdvE2HOoHgqhegIpIlCKkLam+OqxKeB4uLvLePWLrvnX6vAWBmt5TTDjXgNO/Ir
eRGzC6rPPaaQGBP0PZrgH7YdL8Z3RW9hHTeRnh4iABB0DA50aHZcifLhyrFAuNRZKE715qwjgJt0
peefKFyoM8kCkcRma7tzYM4vox70bLy0i1Dv0WOefm+CgLOOHdYN3yMjdil8nAXdW5C1cBgUAabX
gwFD02QX985KWWHPXEypYy6vKFJgBTft/vTpBZbS/JTC7Qju78TGa0oSvw9KLCA6fp1+zYSMifct
nsFHMqa/kDX51z3BqcLYHnHv3R7n5T2nxYUnvOsOpXI84D24mp/dK6R8aDL6rmK8pYHxyBDiawwh
ADa4T1FkBagkL73S87zpGOd7oWufUcALwvrhtQZB4wI2UgVfdEqq055Rm6WYoqwTSYxWd8iBWEPp
gr6XQik2BBlk1Cua9G+wQ4gCnl56O/RBantOYKV8DG5cJkJDtf+AjQI1oBnaEpPHwQCcLs4cSDfe
sckimezMRe6d2vT0H9GfkK66Q2RjjbVuN9rTn0JTayluf2YnqJSAM9Wt4LMfP8WSQeezwpnsXHpn
EFv3XxIyGhbPsgmqmDguVM/0nu7dVs02ntco/nxzTbGc42wlH1kTRuLEYACIbs5Qvh1bGGJFZyfk
kCEOpLn7CMwXmet1ivPkPO1ncO6J5ikwfzaJe0e+qhASqsKpTcdW1WWu/X63D35k1/mPT4bZ5+eX
uxPIeli0yJkQZNLedcZrOpHcTBT8sh4c4qYX4hivHKISNwGeAcI70JoKIul8jWR1mZrFMQ5djdIs
8DI+JDcvbcwGKW2MZRgjV/DEZ1SBuvFtYFKbTABM2lqC5Vb073K9zb1pg0OLo/3zgFjx4wdNhYwY
SlbVrzTLebiIEKxa6Dpusrb9TIkco3940IUigjrXevzdCVc8nUNQfbFGMPY49vgMKqM8TKBOVLkW
anohwkbiCMSajQXBWpC5y3xSn+ipmZTmllawwJS2Yni8vHVFZKg1NGBxKJeLnv1mtpQ3HgN6+57M
Sd5syearsraEK7yy044hamQ5Y4AYbGeJNdlbYMumllcS/Yfo/byuRkj6d5eSp/DWkAqajviCE2Z9
hoigeqTDdHUTOMdrMqhCNoB976lPRQF0M/sRQs9XglSYtGBrcMmi/jkMSyHklhsxjxOUyl7cJqVg
zB/o1ILHW+kEkEnGB7bT68kxBRs6Kkw+vzwQt+FOmE8g+Y6GP3WXTzpCKaIB/0dXHbrFH0GyhyI+
hEHjlNZsSjALwzW5TF+o2VijuAGeMs2xTzcopJd0r0X4epe8vbEnilded7DAZMUR2fNroZgGrM4P
aE7D60x4cc37PMECaDLM14U+IJcRCXH226gv+4snYvWbyt+Q2sRAPpzrvald4lDVe62DMY5OcpaC
0ydMZb+7KORLC3TkXUtGSzgJsZknahPSysrRsFkovtAsgKDC1qO6HjIcXRbGak0bo5+KHMhOm/zQ
yHBMhW8LeHpZ/Bu9TeVbMCkFES8Mypu1Uj450YOX4su4Mn8CLEx9ZICycRyZNcNMpbOwOeh3iZe/
dh37SgTN/IQS+vPGv3ZJDn2y7hCzCq05VD6s+d5K6ZV3sZznkeWmZuDlRTup8jIqpLm5rsSsEIIZ
3ztDO/pSr9KoQpHsu01PPxmeIkIBTz5Dr6RoNrorzNs7PB3ZlSj+4F0pjUrk92X2fePUrR+vdQ3F
8YIjSdbgxCBXhHh1R9+oiifO7HEusxK0E4CBzTY5lCAjTS72MW4FzYTWZcoPwZ+jqOE/DZb7ArJp
0e4sMLfPIWU0RrosQF/k7bUjnTvz8dQ4lsHo3KDxFVN0yy5lFjALQRDzYL4ErX8dovUC2dqAuvJu
+gdjvi/U5Tb2Cd/6XihRqfGuJon0LhNjQ8QWHHXvfEsLt4+1mHtV/oO9wojNdEzBpjmhdJnssPwB
qRayFqwx2giGYk7pYnuOs0pxklU2boHsPM9DjkedT+P9KEe8Mf7uf2b9Ckd+2ip9VY7tepYOC14j
W2fehovcM3T6pVHM4TrBxUlQ6PwX+9Qy1n2/7AznfXjTIrxAYunJEAC3vXL2JTtrCMG+yBgc0glz
XxeHKrrGhIZmPSCe6f9gNAZIXrXAKsbKoGsMFtrKxJuA+2SpychDBYce97rVPbnY/HKqFcJQRre7
6hV/MIMag8pYzsAFvdfEUHkn5InPGlNpOig0CIKVMM/aKKOrJBADKTNaAy6dCbgVHl5Gpv3DdlCV
iW4FvGKnsacX9ha0e9M7lqyOVENMVRBzdQwAzmBvifAlVl0hMySJNkEDCRE8nqC7FGGWL0BHCFPs
5ZVcTnv/AR2NmE7BuXtew9AYnPD0NfM+JTbljMVdGPZFVKL4jBpqfpvJL7FuqKRu4KBvEXXtOSTg
l67Qj6wIbYWzRrYgWHwnaTwxzhuO8NIgA6In8HVGrloya4YXvPe9xHSfiTyke2oHgVAlRSHTO9gf
K39AiXGh6uy5R4HhGUDcP3DXIOWDso/VMafXspg0nNKvE9fQs5XTFvTHDjvf2qQZlGI5RjpFW1EY
DPk43supqsn/N6tSwsg5LwOFHAqvQVqrg93uJKgwWT0ogMgiu2lcjuTU7ntbIrvRb50nNVWdkqaR
1RcfFyUhDGLNWWyLYJDKqtr3OU8HnOvciBYPHwM5tsLhy1ay6SEguo+80pcTk8fgDyLUgggGfuSj
tsWsLmzE/RJCR8OWcI0bbbYWpFVopgW3vGM8oO9JnemQuhqhCfQj+axEM0Qjz1rtLh5QsggCccnP
qF1VNhmnzsso+b1GlIW2TPhBaCF01PHqDSe7MNTsbvcZRZHQhQostZ+gtVmHkoWRjJ61nd6VxijI
/eBLO+usLC+kcmKjRXA3eJPX/5tn/lKBGx87HKGtu7uiOIksvsykG8brS5DBJ5c/EGXXC/po/Qz4
wCp2/lZPF8RhJRsEa5AubL8fSn+zu7D6B758KnDY4iXq1zO4fF6j/dWKSaj5NFSUJglNmshYBQwX
fdpKkIGqjpXD4k3MLTlIWjFbG5ij2K++BXzO8sC+pJaB/suwnjXhZb8+lK8ofvA79K/SqiH7Qpq1
yLBKGL/Gu3LaUGMOzu0MBpojU6XFIhGTtmRVeSrQAhNOt9Kq/xQvFArSkSDfV+dGGPwlVKWQqeeV
vHxF7Y31SrD4gQ19pOMDsGk1OYFLcu4lI+PXlYmCnOth/VJFVIkwcMLmy30BO/1szb6UgvHYPupL
EI4PRCJFcAwokgXGo/oXOxkdqWbSp7dHabyXK8baEBYRWB74He0v3sOVaiSDgIuaLkYtpyL0wTlb
0eENbNqbMiiI/zbMVHd2yHJf5VW4LtDTI5glxYFmwRZC7NCTcGtAVaLejw5GK8Ir/ypvA71/B5SQ
bn58SSvHqqQMlK03SAU+KVvX1ddqXhKq75fLYNgMwc7bf5C9rYPL6HnVsX2EWQDSk6k5t28uNI2g
5Y3OJRHYk2/PJPv3F0eUr1/CcdmH/mZ9WNs6U4idyQD5KlOyPDaIatseBKjQv5So7AXqmsxVnhIh
lMCjL39sIG3Qne+yaGzNguiMgvvlh2TT63ekE/VnQw3n6ROUYSwfvgaIxRv1fYbzkzmjZnUConep
Au6NwyOdKXHxd7UyfOqbfYtGA3XBELFDtDZuf5D0gXDhUhBv4YL79k/icoKYmD+ikGRVKOtyS52t
86VNT5ooT0IlsMGQx3oBasvugxXvWXyUqXREqMXgPwQYdi/mr4aNx2qYC4G4ez3cPAoTxLtdG+Ne
sBTWII6HJSazBru/0Hh9/GF+IUeSc9WGuueTeznAz+yfoiZnAPkiKmtre13YnHzNieTBU+QVVLhz
0j+mRdGqYfl9EEVWqYjuRiXF+RvBbL/5cZb/om64q1QLvLsI4T88fsax7GFRw+Pfpyclrm/LkYWz
7b1pDIzS2JX8vjx0H9txqVfa8bF5KMVWRIIs0K74hQj3JnnD3uVWr3t9zB+HSMiu+4Qtrp41A1ne
+M0h6KGzYJyvw0EFLCHMRHkUxOzJXlas1ZfWgKlon5b1H+CUoYIkZETuwnEwQ5t5rMEhxxeJiRK3
r2lbh9ZGbqGzrnOYqhkuMEgG9cdRmZ21zXfihmAYs7HKhLOP9nyraf4hTOC3kW7A6S+esBbFqMRP
ia9pXt9Pz0pm1KJmn+3ZkJAJ4HYZnfro0h4b6tWPWICcz+z1qQhC/GDnABdc4EjiEL1d48pj3ysZ
ZBAA3kwTmH2525b81+wHqG2wAuP3wjkgz54hqfcjm1kR3Pm4If7cALYxeaKmn1LJV8dvm2kiyYcW
h6sAWwidEyuV+/mb8vlAZyCpWpSNhS+Vds9n9/5pqoOfPzvdOyhFk1OlxO7+zw9v1EQ4LzPb9mSN
PkCqKj5lpmb6aiUuRswNG/GIWiYphUhChoRl4zswQtEz5G1UwzPqitbwu7lKeccKZcJ3KoTSPPqQ
VdXZuNYBJJU1w89uQL9qxs3CJehqqV95UbPHtePp8dnqaiTQpooEFMFAc8NYiygQj+1vQUa9tb3Q
Re0KNForbYGy1lEk4Uz/YVLkq44lQKu049f1zP7ZMecyFWFhbX4lKd3eCpmHoxLuhQkwCMpz9Hge
eZXBhzShAJUAY2ISfdjJlHQ1C6R8+Iq4Ow3C5Hjmpz4KH8EMwYrNnv6fBnNfvV481eGJsHUUHYSG
cilCznvsvHHfeCDx6MQ4CbtKIJInA0q3MhYFrHu4VUEPo9/YXq7rHqE9O3lDsemwl7yRf4MY5+n0
pSEaCxP44OymKxJ/hxxj980djogzbMpLLmEdsBBI4G2w4MUO7kCYhS7t3E4H4pO9Tmc9WaFCQa6N
9hZOnM1yFEXjaWLjESCrfyW4th70TSyxfKWSi9L5QJz4/v1tDbDueoPqoWH6M0xW0zfbgW3ZEWbP
GMLILRsgjWQdnr104EIXi6NMHIWAoJxEWC0kobSrK6N8AuIT0C5fTfIE8fPiznTXXYvmXpPKTrfS
piqKqkzADLS1HCcPheYjPRAVkYMKPbKBNrY4hqUCn5BrWRjVzn+VveC307h+Ep2PTDvuSy3pHfq3
tSeHkB4vZDMMrtVls1BDAzsy+RPGLn5NMn6Rmkwc45wa3bEs37VUd5xB4EhoYr0cGAvwUMTpA9jC
KugO715jBxEBh/DpCxgkkyifqFJNkN2um1bJivgKKVEFnBzon8GdFlJ3uhyiC6MtMAk314ouwawW
GWG9XeL+8ABQlt6tuZFDNLYqJsfkTpe4j0N9NPrGTWAdaUn1EqEmV4bFlRB4GlvQpBifT3gcT+XC
MNPY931/nwFq+CYS4acdiH2AJFmWoXQGz35mBt8H2c01s+FFJVI00oWqJge9xcn01LreDuoSMbUN
+2/5qymgrPfTP4FSQy7bLiTHt2DHWvFrgwReSad0egDHmWSkVOnRMQiQyrtlopQ4WIr4lB/7R9Az
4B8gn63DLbUAcpLMHEprFMmHhGPsKcTduH3FYoNp5fMhuoUoUwExmi5xJ0jkidOsGusEezkWx4Bu
cfFcjdouc2yAN6F3fSC1DhLvIcpXG+Sq12RxO9KWRY+MwG5104YwOLd43ZYGKXaexc4Z1oCRpFfM
KBLjveMkmid0lHqdhyXzqD1f0rjQOj3E5NuXflBtG0bLihT7GjYbOodsyuVy8qv073o1T0BanYfB
s8Tz5F9RXiyptGP+43Ggb+NEJXJhVYTuvlRikT4MWCPQHMAdY4+9as6eVvATWvaSB9fy0MzaFIsi
zDgkR+euHd4YJpQ6K1Pj8geFu719MdI5gjGvyd0UWQ5GRQiiiYh8Q9Z/eRv3fb6oJvc1+oyFw1Qu
+a0s1W9tDtnPx568bhSvTB616VboseF0tVEZGM0A/H09HmURhVOocf0KpZXfE1YqJtMjlOD1bIhF
PYu3+8Ne6tk4Iz0mlp0r2cPUubFsj4C034fjQXbrzw5MmdZD8af7IRPusePHkRVwddmfnFxqlm0L
pkrT5sz6pEvC6sEbmKhVzVJmFNzg1ixkgYq0iVLYY2AxCh/MVDg7GHz/vBBcKWKB2BK4nQ9c7AXY
O3DIaa9OUoMoOQGtp+h+QfY/+DBB9ptnzNnd0v15A72w3IxwgFisggIa4/wLBY0avDJn7dezd4RG
5DTWdG3Y/avV3XRVkgzn/5OMz3hcPXXL+GJe7IQkFJuxyNeDInh6PwT08ndx8KFwweyNheA+SuEX
CLqBm3gby71WMaHXztRocntTYolLF+R/GEdjmHBAOLB+gWs5JWVOyBfSW2w2CUvTJRKhUUEPqimG
qpawcNsEJZnf6h5scX6cRxIqS97ZyoRzFVRdvuxRfORBdQC0qEUr3XZ4lnn3BSbF9ght+eg/4Ncp
IpEuNETZmEkqu1a81XsT9Wkd8ZVt36zwN9Q9QHqsmaoiFhfcpLAjUu2A3/LRKjwaP2K9g7emEK6k
8deaq012xZeSnM+ccLnBeZwjagVGWJRMmUavcLCC+fQR0TAjl3WDKg3Xz2VK1cQq9z3jByZhDpbP
8cch6qiTcqqZQh0yWHrnlO2wj8LRi5VBUt+2xQRVZCA7vqUXG3DOM0AdtXbiFv8DqRbPfUMXXQZv
SwXYu6yNDjRja9qJYQhVXVZhUQ5lOPviIKau/0fFSf0fIuw2V8oLsFIQY/p4kEsGXVg8jqQsObCr
9+Nj8/LI34VAJ0XmaeNbZZgCardp3F9gLHY7GxD3dvBWYL/uFm8e5MacwI98yEKlH+Ij/+lEgWAw
U3d1gXaI2gukeycrF2660Rjb7bNyQvtnvVD+FPXsjSejBI5U1J4G1S2RriPKi51okvdMU4p5lAOy
vuizjrhzKSaOZUVVCi6wCiLEF9wo3p+m88+j1IWHosgGYtqAhB4AOpw812O6N7v2P3fsrrj8Nl1c
xvyJs/n3zOAn6jAPEaVDDN1tS3L3zqlR2LHZZmJa1nxInj1XhcxZXVvnmWryO3pM+suIRkeliPPR
F5Jb61z4yScL2E6HPlqsyKKrrJ3u4i76Fe5vgSuTNx0j/2mNmDGOYvIre9aQzwh4yOkB0QPSnywz
8S5gBzyLEHhoBkDcPc6u9r+Q8ukzmch5Xae/1iioaUxnFlzCqfkNRAKfFM2w76yFcEkw5G9cNM4T
pqu+WqM1ahZbr1tTs8S1wvkEVvQ+vBbdjtNRXrx3aWyrl63STp3qwbqGvrs+JeB9cCoAobtXhMU/
Hxq6R4lGzRgemA1vOuh6AwZFbXeKhnHqhXaK17Fp6Zqg3puHL7FELteY6CmcieueVS3wFVxG7ysY
fyHO2yAL/hXiQl1xqyoxo2ZOepu4RqSxJAVQM5Blx8Bh539MPErbKKpYdr/9A9o2/t6qaEXvFNQ/
kVO1qlImmKHtCuVdxjW7JRKkcurNoZrgPtwYCM5E5p6vTcGmOBwwng/QtkrjeXsioofwPz0NCgnZ
RCwEXlYZkjrO+aTIa6TyScDxQpRtsaQdagygFs6XpWjxAYJp27eIsWWCtr4bu7mEv3SL66HkLSgO
b0F+qSveyXi4hhIPspGGCif5kWS6JbhxwmUKRy+CsqQHb8pcgdwyTTPcpen59nmH94vc2NKg3nJw
j++S1nS1cJx28yXl16bV0GI4cT2AGbNoOcjwYicVmRTXbssgLvWQDVOlXioTV19sxyYcA1+B2lwY
048sYhf/CQSx0O41o2uFPK47eeOPo5UmkeiUfZIGERr6Sf7wKeG7j059w1K5uqsLUvrzHdBqn+H9
cT6Z1Uk7qAupF3e5mLQmA/BCKRfbA61Y8KNJNUH5eDhed2y9y11Z7aBnEQQ2Sg3dGjBDs9zHEo/i
YeVxLhY7ahVYCztJ93ctu3yfZaf+fphIBHbLLX5WGy9U2EORQCg7G/3XtrVUAbr8VobyYFlG1c22
UQyYW5EjTjgFbwG94gKwew4lCIAf74A+06JnofREISaxm0tcBK1yR1Iy6IxP8yCXKZ/+JHHiAyGI
ScPCVWF/VNhU/vXkB5/EG2q+IAn2+JEyuOeWngAwkMoL0VEB2EmRPLHyvxCw4KN+zHsXEZZ6GOtK
eGxiHPvHfSQqlfcAvRMBUDCuwJOQLboFPpzBYMJiovMYdIVdt07HC0S4BYOT41OGdminz2UAhx3f
b96/MwUzV7NOpUV25eMHk5RnQky6FeBC1MuVK2f63utnM62BSqaNSkg6khtLAS/G5JN0pfwdlI69
ma5SusYWynRlJ1Mfyf0Nsj9ilcO6eXijnS/7Qty6Tdvt7N4+eMjiqtTtIxZN3qz2b76T1sEfsdfM
DY8CkBjETGDPDDMf/iVyL5n91mZJnN+5QI/CgcO93SYqqc7KMVTbyvooRxD1p2h+uuV2IK3FNxs0
X7/pIcNFzSCSnBuU7SYDg3olh2O8fbqpv2anM8H650tmBz9dZIq7tctdgy6UwjEw609zhtJGoRkI
4rW8ypsYg4Py8kQO7msDbmIE5pg6kDVQoIv34SeFOGCt7z1pQLr7FwHUgOVqjMVt6XcENku9P/yx
dsp0H2eePRtvPTuKnZnvLQxwbOn1IagdoXMes66Gcauf7qigkNaPV4dlcjLSuNBGK8l7V+doTaim
HEo98/k6HRxq4TwvyRAKxo+Ivd0J/dEqV5tjzaWcFdwfwVJP1b849mEKL0eSacOUQpCytd2a3y86
+zmsPsgH9aCplYuZe5pkVvj6isuYjllAwDJLsEqkfKUaLv37T2+fvY/W1kh3Z6S6wpDMP8sMYZA7
vZhuCIYjDnRjIAagoKi4xKobRiwGDwxTHo/tZAvNJ+Uv/eVhcxCNamgZm/z2NKhO4VH5KSgxnYI2
8IOpz4JLrr1KWeH2jkqyBlYvCgkt3tCX1SwSD0//iTBwE+t/n3UoNX+Dq7GqaFlJcXy3uyVMpXNr
V7o6SZByKdzlzNh15Ro7aTos9VzkqdUGKhyihqBEZUswAiZEDHugLSK0ru1LoXhhPWzdxnpy6875
1tccvOMOhGv3BXTtKma6BBYpYGfeG2ZI3eSYFwH3ZkxxA583j9dkdzD5OYUFK0eWF5egdJc6+J4o
64yTGwtTjpD80vkOeHbjwx/V6deR7J++9Xz54qDBmpJN7vGSsvg06ntimzD8c9uC11NE0qV1B/Ej
W24YeduLEThDyjjeF6lDMEO3sbpGm7G2IaqRtncbH4rRLdc/hw0FKgIPIpUfVbjN6mak1l8N4C9c
m8SDLbG2ITa42fwmONcmdLDIbboEcjPh0pV3iH1f7KXOWc2RdYTiuXVmDPrBHON3Ew2XxpTZVnhk
YqKBOKMn9gckpIL8ibxXpwq7eAQS+GweRJC0pOwM1X7AnOTM7z2EeD2qtyOOGHkf1r0JknE61e8t
DW5jry0Z/8a4TW3DL91DB/YT4S181FCcNTBXisiqLIt4uPLhAU3EyxxNQF+zo/MFG8ZDZKVN9Sb3
+WeORkdsuJjxK8t5YtBAyf+m3nFIfrW+cIxBmFWi7bcazIgkBKLy4qLMeagtw1GJrUoYJduvEWpj
g/pBOcr7oRLTdr3EABUXczVSfZGRNmwnJ+N6WbN+tJB+VmpkWKSC31T7h7i6hQiuBD0oTTsNIqNy
WsglAGNF9FemBkSvyrT2zKUOyhhxWVR5aiba5R0ACTp2IOIoqKjaOi1s7z86BZjJeSBHzPeAkYHi
+1N//2zFVqaYfO9JAniaksf7ODBh4n7QWqKuPSwUHgwkYq73Fv8dwKhWpG+0/cKx8/oeOA8UdlfX
crjKI4zSJJ7chcy///7K+/4y7ZRHrN3HWuF9uE/VAQsCVCj6jYCmNZX/vLw581yUvXj3BF9Z2gL+
nGxm4EzHX1TBhBT0W8IXdgpfLW9Ob00EvmoNIwgwNcwG6ojfKLWAM2HXYvIjgc6yIRixt9hzgNWF
V05RA2g0rXP2w1Me2c5D+ndxMjp9pTIsqj6PJc+K4MUpo50+Vlm9b88oVoq47H48KX+lf4DSGWrB
64OQ8fHsZZXau2NSd8LSZPOxu+3j3fWpw+kVEQ8OnG3/N67B1p0CYs1XGMnXiDuERNRa5oFNvmQr
td9VR4v1jj/JiO1NhA6JveRnovLnEcu7kzrRYpAmyJ9ZKTxkToigBjEeKRzJ8WxVLHsLz/KviS30
WewuKjJejxLaZtoC3Tmtanzjzc2KwVe7a/IXM6MUUMajRG+tOG/YSjg0dPkVkyaLiD4hL+ndbHJ5
tGznM208w0l62LyaP1/syRrxnJCOjxW0ccFAJ9owOXozhaub/uE7cmnOvlJ3MbdFzC0Lc4fn4Ac6
3sbGpUshlP6eTtDu6T4/YnIRXJ16VuWka0ww9rk9gzCNSt4E83xebiQrFNVDq69Sj4jbw3YAv5kG
q+JZEcwVvgwf/w31ockJWdF4eskCWtIAucAgtEMRGFhY1vVNCU6GJ8x9nI+V2rTdo9zfuxbY0XJD
E04IkjscqEgXioXp6KbpV3twvMtOKaoVn3KNsp7JRd+GSfxbeGo4TIB5Mligd2fl+3S0x0Pxu453
qoAQHm5ND7J4noXnW1mYXsmB8mFXdXDuUr+sSnwJzRuEC/czjC8aRnvQiVBBSSzT4upEXp6e05rz
OBlbffYQkHCVdtma+Lqe1ZH22NUQeFbW6FXTy+iA3AM2QvAsLsZIx8p47iVHghK6/GkNgX9xHKZG
3NFF/FpMumq27/fBvhLbH5p5Y87/duY81eLzUJNxgVdW7r9caTXfnCE5wWR5+bQ4QW5aFKRPRLPA
/bVxsZivvacZzXGnEOSND5EJOc03Z1Xdl1xtkoND6ggwjpJvqKMEY+pu5T6R2exdA8bC/V7bo4r5
j/7d5qcdXsLGEI41T5RNrB48REQBrP/9fh97x/8Tb2TLLjY5RfAMvWh12U1mbQ7Uj/VZymBukMbw
trTfsbyWHRjMJ6dWphS/AHN1fZEAOkRLE4DJTFX5+4i5cvKixon9MzE7PMqzEF8JvoiVo9HDRN50
BZWTjaPOwoxpC+Rvc9BbZYkxE0RNKJO36pqN9OoxPQFt8qw6PhcBKunK33Lbv/NZk1v5BlJC6yrm
UHAoDTo/wEsCeSwCkQ3IpfUrGY0vAdQ6xrcX/S1kSxXTgnIV7+U9bi43n74CPcg9gzu7pgwT49en
CkxoeyIU2/WhsUpHjLYTeDqEMiOPy3lwls6AD1VMUZYiFzlVODFFIgylHGpeONbALxJkW2OKs/mA
Ui25eckEW4ScNisDYynlANhh/hPc4mK19atyZQE31GF6EihcNYeBJtZIRu1MRJ0iQJZiV53ohuwd
R8ufDqnowq+rUlTbEJZUDeP0a22n30gg7UjU90dGI9sQUGHx5ZUJwJFpHgXXaJ6QhINNXS2FPz8r
c8QF8QMOX2MBFID8HZKfFIISlPe2opKJUVkKDcDoyeKTtKi0qDtHGdLeDkWA3rf8DhrNe4xqR7UE
r+Y5GhSAoesQIi9SF3gjXj+c+f9QKTGvvsKXBNCBNZEtSdKMqoe4uCqxa60927llRaDIqsXdypJp
17a/6Py79pbHiSzKqtW5CH6DpFeIMkNdu5ZdoYGj092ycxC15ASHDG1y0WfAoRJr98QZEgB0M8fd
FSmfCfeZAj0FOHxHWFMWShZPWY6KUH8tfhAS4Qxq/r9stzmIvZN9f6Tc+j2d6pfNekBHAqppYK53
60W9e6XqBCGg/GAaRn0Eq+pDsoxMrdyxwmZwE96jws6eHJ0V/1Aqc5bUqHVxlpVN8tUow2QDADDy
Z5w+Fv5olBB9nQFCGPiiYYnm7mO2J3KroM95vChP3tA/3U6W7ac2oGY2AJwd+JxQu33SfFVFGVIp
C+h2gZEiQ4eym/3QUVTeremYOo7if4iAQVJjyyKbXdcqypGx+lBdZ/dZ9TmNMx7U61FxN4tNmlzT
oT3Bquha9xezIMOFJTt1UWinRtTxC/382uC3y6HTHWtQRwztQiEBtRgb1+sEhkOzMW5Y4wccRkUV
Hd+J2xZLPoRX6E+gKx3s/Qs56yb5eC7Jx8iuWAkZmx2kLf2zByOxB+Z2c5wCsvvebr6brotfyS5A
a5pGHUQ5A/Sxeeq65BPXEFeYUvJsia9MNncJ7inY+kGaS4tYju+A6xDXlCOjE4bq32a7RUh56V5J
WlPHdhrX+M9fspdljSaJDq8faqWwG1/c/vnoZ4mKBrexTvNXzquCqhn8xdcdUhskv/2EIW1FRt0H
uRn17PxDI3wYA9HZbBHuixNexE1oPQRHW3zhhGEfEGggYDrviQLnNL1MuCAWxF944x3+2GOUF4Pf
zzeQcihpPjXnC4xS/xcbM9gfA3n/YxadeYxrdixohBYuchbyYfZ6yY/D5htq3t36m+A9S/GT0uzA
V7Wb4TUcURH6UBS6aEkHNKG5bs0GxUhv6S3MMnDj8iagG2BfRshlCPWkxlA6OHc9ivwLINo09JEf
vRhenzOFvRW7M5B/LNzObT/7n/6ANrt9BJZQ8cFPoTEpUuwsED9gVXCCenV/ENx3zeJnu10KCuhk
Gdthv3/IKJhoXJFu74o+nis1XdjB7946hFNIORoAWJBK8rqzba0StMKkfg5weYCEbPgP1mImD/1S
xGPW/h/0rit0H0pVeItP50eIvSqZUFyFgmZsAcl2SHyBQ60/XlhgsDMyJiq5qoP6GO72j10bKTvj
H1aGZKWUEh6shncGrvw7gp1H1kKLBnHTqZpncr5D1hyh1diUKxiakeupa1ApN9CYf398/FFleeFz
q+xod7MC5/0+TPHKD542Kcjn3AB5JKybVju7Aj4hdQPLOfBCv44JLw2aE1vPoWOiw4KZPabUANwR
JJ07jfPXD8jWpcxXOrPVeMzk8xqeK2BBIqWqI0ETrv6ykv9xG9BTbRwLwuyVMXtGOuca4IRmtCF/
M4OgV5tGDh/0DnPNw8gqoEVz3EoCkGqkSc0fE0Ik47r5/usz6fboQbE13YuscZClSasHP6QoVT+E
M+AxcXlGI1Uhngj7cBzLIUf78kUaHHiaPV1xmYattjUufgSiQ67v3icIKQiyYVyhj5/ai4TMn9TR
mR9VYv1cNGdj/ghVQnD+Cn9FGR0ODxYfhOfgDnA/U8Tis3mk3iDmHUTNpl8gn9a6TfA12Bq7SNk0
+VglkvwzIVVIdvPC7Khbnh9wmPiwRBb/Eu0heDQ3VsOek06eTfwo5Qe5iN/vRcTrBzsr+t3XMGJM
TWUwt3IUTxNCSpn5ITDcK9gY6yzTDf5sy3Noiy6gOpwLDcMX2mXNJS9B0Lzfoqn0ERG8lYLoUY+C
EZDOfyTCy11uVFJ6TVeTC8bFbjm4sLKomzjEAajsg/x5QKDsaJ8fmJumut5HUMg3gFZRvPn0uLL9
/i7DRCXYy2TVwHGVQq8EykdZ4CLZpMJIZXCsCVonlwIi/JvaPYCeoNNGWDLqwiH4favSStVqYLz+
nrDk/WIuEFukfI0Oil/B5gkYS5O0rQ6Xyn8q9jCjFe+ikpdcH2wQcgJrZvAsp99sK/1c3j1eVpbI
f8nJCHzBdSy4p3yTA1+9hbKhbSAmhXlHspH5vOVrN5269jpwzHO6+uGaCLoBwWaJbqiBSAxzeUoq
yXrHJc4qQFOwQDwVCnOy9SA4c7crTjy2RWAuCubIEJ/YBgEAqMPuquDLmaYD2qBDhBNwTQyq1iCY
iVVoomHXRp3TZwfpVjPgmwCSC5g7eASnnAlQNQ2JN9xSxdjJ94l9oEOthh6epUaN0/Pg8djhmCXu
sgJyj1kuIohCC45nsBjbLErhLD+qEmto6VFYv6NenAPcjhUxAJkxrxFAOj2Jhtk0K2eaN5LrjjAR
91ANKVJGM4dCi6iUs8pY33XMOEijFwm1SF/FME71A1ruktevHxNbZwCoBxRxIOL4JxAHvp+xxqA9
EGkmARqmc5vkeskqCmyWXsHapw5FnKFuSrw8pE2S2dUvxDsmQMliMkggr+Xps+t4Vv7me8eN+EN8
3Uc2oBvA9P+JGqpqWoK9WM2hMbyJWjMzpKBsQ9qQeYVE7dlCJs9q65ibAy0OcxozDxbEb8JzgjeH
bewMVkYETPZK10hmjgwnBj7UxGBywCKvTUvJOHdCF07iZ4h9lKa1Ttefg2vwSQtriCYh9QZn4E8f
yiNidDYcAzsFjiDLR151aD9MSTEhc6nXaka12LA0bD972SkEEz9m4jpOoRo+VK3ECDRKG5azhgDI
4+GqFcoWe8yD8of46I8n8cTcVCoVyaQ3TCAyH67UFQ5/nPFKfU91eYIWooez0Bu5y2R8SQTXTAHF
COjlQLsDbL12C5LX/uwzefwfkVGRuvnluUfVZFuIV9kZB57rV2m85JapEhN1hQG3k0lcTSqeWk0M
E1Yerea9MLCG1+0EFUwZroqTO6QRmg4Envteedua5JbXJhWNlZGKG/epU/4KSeqnMrbPK0TYdFA7
5AJgW/x++Rn++zzLwKgbv9A0hUsKqVC4K4eKFdCvmj20VMIeAe5enMpbd2mldC328lrzJhZLTRqA
wlBnXMKYY1Rgjd0FMvN921fekcr+a5drDFM5rz4+SkGyqoh9zb/xCWRisGHPreiqlIgxuq8lCrh9
qValfLIgXmOyEyJJg+KETcLQoSA5IkZbHn6a9MMWSthrwBtWfcqa52vffZL/ULygpr7Uv1wBHY5F
3GFuNosUZHP4LGkZ1Hvcxn1blsJK2os/aoBNHuwapxqpOGv2dkTZ4mYtoDKK2s+3YRXPjwM1rR5W
0bzV3+/DRXQ7UsGduJo+KZGkSkvqPjWsHOyKluvdVdj1j4IsKQzsWjPAIbOWnX+5lpkbT0MUCcJe
MDOFl3JGxlG6u8Z+JkUeoB7T4u5OKn1sQOUm9COU/p65sMbYkKsRnRZHkOpXKW1EbXyO2/yk6zgB
dtLvWGzgRyw4/0k22BdZ+VRm/ctHFyHhU0OWJF4im+v/XniU3zQVNvD8WELGHd5inMI0GPQz2N63
0DLvsCXXhtwOfL/kW++V7z2bpJe5BbCTORr1hhKKt5n2h6pdTgnkJpEiM6rC6izoVHlf2FvzvJyR
QeSK5nMZUJAD1e7Wmp8TLMgpcJRKYHgLmPkcNglFQ+X2S7/E7v+iAsAaC5mJoh+VtOiQ2aKlYLxv
7oIW4gxcx6Bn42QfSQerVuP98943KnrXDeEW/aPLkPAFQN2KCbU5/SwbSJeOiL4m/pECIQAsQiBy
4HLrTP+XUc4vN41TgvDZ8R8s7NVLSaoR/FQsY9Na4Mc119J1VF10zXlWslmawpbd++Hg7I6NeeFh
zYVkn9SYt3kjHuy4drSsA/LyCWN7LORTbTpVcNtAQD0uGpHScUpKjXWWiZHkHhTehriNp2AEBKFD
OFyZ1Q6tK0JmqmuQIzdGQi9yH72iwnq2kYUEpzzunrYbPGIeOtQ5T20xGUspButBBLegvlfRwKBd
9NUdN+Y5cz18K41l8BFBQh9EMNGp6x8isWwAuhaQ6b19x4gfsFWBz0smOZVxM6CM5UL0iyoFdJmF
A34v0Q9xrwCno89VNX2+vkJbr/uvPBa2jPpLWChFczlE/7DyQpZ3zNm3Y/h/2hEMNGiRyIPJBv6w
5DnbtY23AskFwfoCPW75WDSRG05NrZzeBUCrIv9V4iQTbk/1UF/bmkHRjFgd6JvM67LK6emX0sm3
V8lnp+FFo6Sp5J9189259MRZ3IGMnwCBA4GySyD10sf+XmLiTUL72UNzwWrfQOrKRa/CI3hnzTEj
11l8kFk6gpm80HjztHKSXJJrfGSfcFAjDHBoltSPYLrWHoXN2PvfITuR1TaGzLUTRdTwdQPEBTMm
V7LYBv8OUxMNswiXTo3oqw6yHFBcAb/sjnUjVBq//o4tU+b4zwHSOl0QtBYzrHHiSAAyPD5zHX81
Q2ch6eL/w1Px7O73nxl1nMBDUDHujIJD5c7ZldnQHUK0GTXZ9uKWKeN7rXPAVmbFXqPoTDOs2PmV
A14REUScepFJ3A3RtnzNgtWQlsYsxRtcdxJsB2JNTZ63+Gmfg9H5r9ex4dD2kkRX3DM/7y/KLU+1
7yualzb7tdLfj9LhmvpALOD6MsoVnrK7QLXfuVkMS2lCTVFP3fjwWojssLEzX3MWgm1PqhLNR1ZG
SUTbFlfA6EKphmSh+ET2CI+xxbC9ge5ux2hacHWE+SY+E3TVks0tp0yp8Mpvs2dZVdtqT33zJZNO
IAV+kc/Uq/xPo47UXziyCIFb7OXUj85wJl7U3HL0kLQFy8dl2yKiDz9Hc38hHc7VIeaxs6tKegW7
upZu16m/p4U9zWrg1ltmnrQ+8PxTCg4iKbHNA884NP2/zWE8O5F7pzrbyU2i8CYe2J2URUo9UiW0
Dk3raR8r4QjtDmbley7pLlz0lDbgN0Fl9RdX2jSsRUVoh44QswctmGy5lyAr1RZzazGLOHqFgVfv
K2xXGWOqxHBKvlTdqLNKBoPt/mqb0t67TJCcVTbo16N6V34V8ijdI76SK9QDgR6H2KAquCiJ+EX5
Dj1p4n9DKjhRhwv2iBnXSANjWKZLLBxaWihcNJK5mQqh8maELeugWe2IUo87IE9OcdNE36NXPDek
ncLS/FOuN/6vaVVcJPaKQzWaeRoAQkI3wQUK3OLwUZnpKPyH8bwtySbqxLP1En275N0ZabU2vk6J
lDOrVCfXwRGd11mVybJURx7ZIbiM5CZj/tF7gS0FLJSQz1vl/ImiZi5PydEA32ACDE8ilkD1lAd6
HH1wEceemWnJhA1Tmgg7D88cj0elT8XBGfokd/z2iKVMZXfqAcp+FQK3ahjreNB8bIdXdt1Uxt9W
vdvw04rlB0DyqN263fZim7mx0DfcPiACcqhDfxd1InT3yFJ91/mS0PSPT5z7bayyFasIsBlNoJ+z
6CObCG3iVzteMVyqLhzdQzlN2soZ9dTxTTQ7I/v7JCwAfk7VCb+hpn7Jc1pKeSFj9rvxKZTeD8nb
i4ATxw0Uwm9FEzjrfLg6XAlNe2i+fO7dN6+G/Ao1h2ik0GZv8P+9e6U2EmLhmJ+WSTGbBp6JTtmN
qq2qUlcTOHrZpBZc5qYS2xiLp7r7kORHcfbtM/aYpPXlsGQf5dh14wC4uDt5/RAq8aNfGKlqUneH
20SqvcyomGixKxV0xNaBpnLuyV++A8OQRz5QieMPUEERwX8+zr73Z5IKl/+ZUqrQT/gKr1nrKYwW
in9YOp5GIV4Se5zIeOntzsrxh+Mwu3uYWNFaTAk9iD/BWcJwgbVmDj3Oq0zPQF98T5qmL2ddSWtl
XZze5k01+c+PXf2ol1snI/nxjDgb3DB6PLNwUdPbNl9PS5fn3a6UfbCIUpysiZMPOVada6zwZrKd
2Lgb8nzADrmSvY6fn7psyyKBBcbFfO+j7yNOsNSABQj7pa0EpB7g/0lXIUJeKrO5bypQpP7ecZwS
9KmGIUSxHhf+RTjC3MRI8YzqhAZqur5Dm5EuErtnUbvbz123gf72uO9ZxWEio4nbS7nniT63vIvp
HplvGbXQARqqOlVlGaniNCXz7r2dj/wXg6W3s3ubkEhxpQqOeYNdFh/3WkSN3wtTZx3ElUvUTuSa
wfXJLhnAbthS6MmygXccfEaACnifxGImzUV/vc/DEZEuKzLKl8hBFSITF+BhEpUkXL57VR83AA0u
NsEsLffBSw9d1d51kXuLBfgR6tQM7nll+op2rbLQAQ3H6NgaYrRtlR99ArYKNZrgimHIPJ9tlt90
FCg+ugvbMoKmU6gcVj+F/LQ31v07jqYVMmWajyc9oOBRz4hWd0YgGLS8hzt1DAqdhuNXU25P45ro
nAFaF2ThAjKyWkKalC7t3XpgJ5oivElgmTSfqoylF3176mfIZ/kh7mUS/BVBRFv23bJpS9cAd0we
V42MukYnKYDFxJ91WZm1zG5bcsH0ZwxFu7s0XAmIruZjx3hflT7tWnXLAqXtmuFaLLMtWQHmKASM
8J+t/21fVulERjn2mzHtlhzfunbH7HfBusui28PpRXktvjfTBZlOQaVy/sDe6KWcCWhlJpYeaI9K
eCPvVBA/Z/KNhLvMq7ZTr03srAs5DA8E0s4X8JFouC1yzYhEKJ9WsNphZBIk2wJx56MT4jfkF480
A8Jw22yV5EGIdUWMEoQ04PvRd88YkizRRXMwPHc+F8fdh9gSVcWuvwbh4jFuSymWe4ppFva45d6E
OIfM2q0x2Zd70zv2F/+7AXOH8OyCIlxna+vrv2J3nXjacKlgt7sx9HNG9kqi2hcWCh6XcEPcC6o1
s/QJ8MKrvNKeTxKs9+1aRu7d9GamaR7JKYfhvQO0X1GFz3nhfXBGHnl79jwBVRjKCyU1S/QsyiCg
Zg1CIXfL3qF5SbDWfiQFaYAYgNphwx6HvWXKirDKn9Zn1zT9juMWkGiBL02b8z3VhIoxc4qKfl/D
9BI3C2ZQ+GI9CKFqOpb8Y+XA4lYSimLmcMJhoWsUip0RSDDrvUc+TQ915rIzu/0xoSHWm8ojGQb0
AUpowbLqIL8L5OVDKSoF270r+3YOi1MbepGQNCl37SwC9Rq5atyDK8gQ70df12uQkn+gxDUnd+y1
mSpZrzOxXPbvglRrql1AFPG0cMTYqye4U09eSYWTLvXnOoGxrbV7o9PFZAEKej6GVA9NZ6XgcpoU
7JyzNjz/KC5MfgzXcJgCpyJ0QdTiqHlJLaq/hZEMnpTjwMmiz2R9KkZxUr5/dMT0m1BuFmBH8ZTm
6ulRz8Mkx+IK7V6TxgqACJPhLKK+9szNbpW6UGAI86RJw8bSJ2rixhcn8MExEbCYUj2IUVKgbS80
KPkktfdtWl8ELzit20C1RiO89AHctudoMjdgkqF2f5i/DO5mIs31Ef0OHmYYHMyJEyDZn3aZ2PZI
FjNl7Btao6Fxk8jY6ZrNRnirjS+8SvxiTsFpFQ33E7O8c3d3cMNYkSUjrX3TrHYODCzLrmZNG7qz
6lEq8JAjm8qP8LkRI9mQuhEL5oGNrdMy8las0bUWukvma48brZzrLPhzspJCyU7yuHn/5NdCktTS
4wdTOu1rlBdVH7gJWruLvuLmzDNmuYc/mM7bccKiw7zsObAgNIIJCMYCcWedAaKb/S2L7Bmkxhg7
U3z9vxXkg+kkvcC0iENJK1n9UqP8A8UKQJzAXEd0FALQEMXrQmnZV7Stv7FbtX8XsZDoXHKm7xCa
XFzLbGJW0f4Yd9lmXnsw8vjKbqFEZ+wPD092/CxjS30B4YHOnYTjw4LV1+C9F7/VpXYyZ9UER7Vx
3ZavicjnnAUgHPI69rFgXUK+bQu9tRO5r+YU3M9+xaHssZYT3mn+Y865sjRVIs+rB+f7Z5c1Iqot
BMmYHbT8k50lGNKO1HnrKPob5Ex3MqRBCmgC7hI4tPQtAa/lCr+w/KZAOqsml8vrpzlupDH9Flpj
INpFekO2n5bHPRKMRIGdGqwufbK/pM66XGl+eaVVjzicU18yvZwuKLgvND/pUf2tGN2XTg4R0nRj
z0sI6tl8cZLy02emd7DAGxZwN303DFKCyBQkUM9SZAe6aLxti7o40azUm7OZgfPNjjVV2obduj8v
Yb/0eoY1zuXOQz/5udmS5Yx1PgP4jLnCcYOIAxvUqRXUHcS3ZE0Etim5VGKDKR53/WJizA8o8fS2
ENbcWKy2T4Go0YJ1U5Sm3u3jq8JkUaOyJiSvnQz5wbmXNCaEUadB93gUTmgE99UUGZmXCkSBijZG
gvOFWIl0GY4pwMvBb2SvNBSDIgUopBeOIL3tBEkIV37YQCWb+1EgNS2VJemBQcTknEMZNqzhneXF
o6bNPl9yUz+f7YjvWfwOjmhU5VdKSbNTZ22rgtFX1KtJ8hrAV+eDzpAdLZFY1+kiBt+Gr+mFPAvk
Lc37irDdzFZnRPLE7RCPjOoBN7mUyrUnXNkjbIXPWEemr/q5mdRcVQcKUg/XYUiWCiYnxTudBy24
X9VymOt+1cNER6muhbQEXJ2eW5IXRmAVRVU6+wUGRsX3+vz7tyZGm0UVzsTa3SI72xKZkCst9WSN
EIjgrK2MtJiNnFxMjt84wwUT8RblFOwGQD5grY+arNwZUe6ciPz0SDvM5fVksWOiFJNtAskSo5rV
LfFG4+c6yPzY1jRdiwuAmf4Tc8YG3NB524tjhcWm4sJxm4xYMs6ogT/I1aYTTsx49KBrSBQ7nWHk
8sVVRr911rYcOCU9CGb3/U0WWg7mvq+MxTZtD/QBzae64IAEUExQBoJXVapQZ2NYo5x4g7rj3qHM
u3aX7at1AxSICZxUzIHh7bIncZ7A5zyyoVk/dTMMDaE7o/eFnpLwc1B8D+m7qwwasM+0XDKEolGq
JXjjn04lQX4YRtN9MZdeZ8EwQZ9azE1SgODvzTrGYD3BsbOGT9elaoryfIk7CYRdQmuK4CvhBgt9
y7SY5yZNkFxPJvm0rZ+d19zvXxH+t37Vq82HesOpxtlhbzSm/AY15V6sdEVgOE17XMGN82ONA0zq
uU/JT07SeiPTFV2syRAtTdDPxysYDb85FgBk0FOOwsQf7fDvaGNWC6Wb8Qxqxs3UqbZi3T+t2Thp
kl4/fgc5e/eEcGFtkx0rIC6Ylx3+M8yO4g9BOIxQIzMuWMsEJvuuVfg0fvSA0mavarC0AfK8mUkt
CLR+pMLOjnM9pxL4cd0CVPiz3nCqpNEWcS8VX4ggvmbxsXHums/0tWubCqJvpArw3cthdhyQwtM/
fK/LwN3Fu81ahS/C8F0eVv83LeP6AOuU99EV/4Lm01ItT12SKgN7v8jQ5+7wzLbxML2yR00BjXFE
mCioCBy/pj+zakTp88IAN77i2zwIUysefLlc51AN1mzNeVzF3Vd+36qiq3plWxhN26lvRBhbsn5v
06afIKMoA3TG2csuecDToRo0tRT2AA/baXbr+4JS1zbvwIBLNgW4sgglxPNUTRCv2rniuI3wm9dY
kPlh4GeBYQ7C/GqfeYhZ97zP6zWq96lz9Vb1AVMmGDmg9/CKJYY4IlCKC28j+qHcwsACZqLjrWhS
4ZGgZjsGOPT86rtz4bZdSoN+J77en2qlf2lYYHYfxNfi/T9FUjqiGiip9qGKQLvNHBsomK3yIwqf
36/Np0ojMkot9UlT4OBaMz+T4jvt3bpU3AZ7xGsFbD3Iun+qnuGdgGSMRXaTPrLWXjSPmt5insKs
KNkGB1x3Jv/0t6bBehl3wfE1BI+aF9Crlq6M2UG1mS8wNnp/ULwEhaUiPZe5nTci+TM/bp6miArI
lI4uv3hwu1GleDrRpSII9WuNWDDCeXn6fR1sRYNzgyP+Ra7GHNY0msaJNOP95IQM3Ko9nHKF05VS
diSb2jkgzIudxokpKlji/g33tSjNiqAe0eqFWoZIeVFOB59AIljapBj1XaFJwcTVWhCCSVUtNV+Z
cNI3VcIY66u4V1y2ME/ASvUOGBlcEZtY3Kk6zMQwH8jw9tPfFVV4XI19ziPrze17u6+UIXmIw73b
fnSXYmeUxOEmYmFmDiz0jv+WXuLnPSDLzwaIrCHMyxd0CfUpC+nnYgABj6IurSBoBcHGU3mmNEgV
WynwtgbNBBB9uol5r+dzEZcUhJHyQ8uowRVJ50pqVHp79qJ5CXspvyx/9SeUCY7SPeRNOLusnrZa
goOfjZNedf6BUPfrk1hIKh9URkOuzAim5Vz+cYLV7UGFGcEJDkanx1/42e79Nh4e2QwR+PZijJTT
s5GrpPpENkHyptDQn5t0M02TcUGF8V59iIP1UpLzkW15EFbJtJfA8o/itrRjXOnZy0EPkCxsxk3e
xuT6oB73fPlKETKQorQzdljFR+JrohlJ/k3YNsw7GjNiChOtYwktZsIAfzjZb5VBNuTdBAmvzNbU
p93pgRd0lqthwic83j2aAE+Rps1WP6CtTbtuZsAktQo0AG1fkFEfxABP+JdLiwrnrJK142IndF7y
6G0C5PxVt10P+bavgDAbOZZI4xtTFAsTu/emt/CFrLCdSnumFINk1LRV3JSFplidOX/0tYorKP4F
4nU2zGqK5snPp8VfM9IHZZpKGN/JeIaS2KGSTvckJbT3fafEnlh8Wak2rknEjm7FvJ15Axr7BSJH
Voz1HW8XBevUg5p7X9OEas5UwDPBBUFHqgP2UUxn1RwOpEtj8TcWogotNrT9UVqVA8yPci7qtdGn
ineyDKDzawbU6BgKAtFxnl//tVorm7UQETU4npCkt4SP3EgNIYNPfSBH9QSmxIrEYpdnASOUycVH
WHczfJcaOoOd7O1Rcn6nzGJ8Q7Yd7aSJE3s1oiSdy20mVx8R1FQZL2kIgmmixyvKHvHIJQJcyqlC
hiB36030KWtlG6SSMeNSbIjOXU39wYutk9dieu5/cA0vYdeEl1SvkNuDc+4f1SXZB2tu/H6P/WUe
ZGtG9/yKAyX43Da2jCqg9R6+HWXMoT31iDRsPG6oZn+NXY3WVJRlc2n12wnVIC9QJanF3aL+MgEj
6NemIXivd2S0jL6DalUFFhMSMB8+wzW5ghA+9BwxNu1t1gWmDbNQWgriEFMgXgsJHyrIoK+9dE9a
aFiwya62OhMuHuFLuAkpDPF7RWgtvbNHb9z2nF/ryWT23ZxKOtMxqyKx3aPp5lsSF0iDWimYebh3
kKHQjAUoVODrEqJ0J2oPCTVZHTW00zRzDZKr/wCSjjTtrZHRpkNjyphukXOOJop0X0gF7QTunwRk
FGKDGA/Z8Wd/S+SgJysHWAarQ4if9brbItzqCNoLFrmxyxRMSaTMdP4swIHpKZ1rC0aa3PIv0Qn6
CPN01zXGhE0BeJp3XGh4DW/fZiaarFvjmWCoAK8l1dnIjbME3gvvlZt1zOyiOFuzzrzQlCEudxpr
Re51cbPjvdoJuD6fxrRwYRQ38aAByj7R4728HTpLKnF4pAO8ByNnVnBgkDfsu6fv/IPLT7jYzPXi
Wllb2zxmOE+PGS0NLggtJ46kuN8wFpd7nKVw+NLONXAb/M1TY7HwNPeRkN854gk+JQtuPsnWGHZD
Z1iBhdNfnzqK/e9L+LOu2onGjfa45XuI4dqxn7oI8zlozDDdh4CeDnDa3JSofaWopQkcrx8OWrOV
2vil0uNccNNTqKlbKlt1Jm9cCO5PKpgOC7rAUmaYBi6Ayi9j3aINnu7jkSHiANKL7AWLHaOwSZAe
3cc19e7FMOyeqapHavhKxGQDBmZuNx0f8FHpQP77C1OkNwKSVKcfblbHEoNM4f1gyeIxEDIYVYKF
UFF2bbh7Vz/fNeQYHox5yTE2Rpdhs2t2QozQyCKr3YU75w1e8yMt03zQoMyupLKKPboPhUVTC2HP
pfp006UZfGp2km1JUYxPufLuU/7ZzCuYn4fESqTHM0SoeIERm3htF8psyYypn/4DqtD0TUzc3Eh3
LieSBZmbUukfX8+XtveATICQJy2ZGFnVxoDF/cIS17fvI5zZF8/NrwBk0t8Cqaz+y9VexzG6trBg
u603zGd5cPZX6nBwIJTJIU2WlYxd/P2QNz1+S1qsa7xQgdEcEDzA+hwpfioclGNOFF6xs9DKqs2M
MZJ+vwCoKt2sepZq/NoNZPhp+moVKFL/t/UVZNLUtEonYu++mpRQ/rueC/Kown1bbE5dRPqIgIbl
eWATRbCHJFUExEpZzTdRIf9gZ04FuRaO4J9Tk/KS+kzKePmTrnrk8T6avmGPvMOhW6JOgqbxDze3
jyS3jejZeNTKQw2onghRZVbDpBVy6xNnUnWsicBnIPEqJVPsBzxqHYmYKmgtT6JDjCrJ3hsLG7sQ
zG92Bhsedw3JfBKwA6ngPde3yBwU1BjNZYhsxKClpVNdG51XIYK90cMahGyklES2YCMTHFFw2NrZ
6j+T2cvdUwoFKilvP/f//kjEqGV1Cxh1CeElNs42qtB6E7YO4rV0RQ8Uhp2QkVBBCEXHwsrfw5VM
sU0j2fnRcQcUHPEyK2LkiFpVCZXJnhnpnnS7+7ITLFYeZwPL1rsb1CwE3X06CpMiLjkdnDAUEQRV
dyBFnqmWJFPNYfZEyAx3V+ffefU69ZntqaLaIzteciIbZ7b+mXn96r1FMbZCisSD/Cw4OdAEyQFG
PAK6Zojff2ruM0gMOuEVsG7crQ1Z6SXwx2nCsSrRDOIk8M6ZABSkmyu85r4sqFrX8on15DafkiYr
NjdqNLqJ8SnZyi5Lrm7yXlvtz+noFpg16YT+/S5voaGYWdpddQFSLZS0cFsyPewiaOZn7QKtnfDq
xU5tcChV4kTjXLdE/ZM6LLs5OdvQn1yShOQJwKLT9o2twrIQTX+iOmZr5xBhgY24yGLpkgv02QG4
dvYYyzJBsMr0BtR1qScb6v+l2WBV5WRYdJ4yEf1XS1T9I9K5DWSRO5Ekyxekn9DR2kZQ10HOHzE8
6N5kLTnaYNNC2LA3eaLudVUbt+IsBdq2NhOqpn626oFvdOH52Nchqgt0QZwOTmBUp0DRYKcD9Ada
BPBCI3SSHXxAeQcdoSfbhxF6VXpWGCZwFCP5SF+TOaDMRa2OOEK5KOTeG5+76JCLyAWHPrgFRFl4
I0TTh/eCdO/aXHBfR/xa9FISRbnS94UtvA38Q9XtaRz4jjb6BME07r7i3eXwsicaLikb7strquAz
rGjvtUMl3WCv1fkVFPTV6DQqOAI5Yddv6GzEBkNjM4bfHq+mSxhVL9bGdB12/4AHkmr942MqfOdI
yzqlyFuAYV+oM0/l/tLgwOCRq9i26kMImwnvyYxEP+RPMtZlKhKKEb7WTRcpfT8X+5w+I1MVVvnN
DU/oYqmpvcHa4iBvCels+wBBpK1JhTQiFDGdPGuoDRzvZGA/0V9OOGt2U5c5gIUN61A1fAZiSwC5
cV3xshdYeWWQuea9qiAjtN46tP0J//LfWA+lRfyBk8RXPlyvN4m73/l0ftDuKHftGdYENUCJy8jO
ZTDEu3CyznYi+RaHHoYKHUtu6BUktnbGc44aCFtUUGsImOB5JXXntuxMM+a1tUzFOWXNHj/m5Rlk
/oUFHiTPurxA/2164+q1dWFJTi6JS92Ta5D/tKbjrJQ9uY8jywY6mZWYWqDPy6f9YoXxrt09YMt0
2Mjj76Onn7kfUxeuTLfG8UpeY9XDELywgi3Jnwm0JDVH8AE6hDsUgJN/qNEcO/CeDY+7RaJNSkYy
J5bxDR/juvDeTDWUcGwmj7wRt0itanRwMl6MtYhY+JioJXrF30AdkjGagzVk+CW3abNbQqQmV9bk
vC9yd6exXNdlDb6IIF1Cn/VHi4+o7Z6faLPyFO5LdK5uMD52EhfzYXcyQGIZHxMDCVubbQ+bc4HQ
gJMReAk/k+fzYMxWCoUlsvUyCgYdnk9OLW5iMZFk4wSrDkmjjF+ZQ/iXMy/VRnNBUVkfTAlYj1mV
0gzWaT7oroPU9KVVQK6YWvJm4VjNgRohmiQrni9wgKss+ceW1Pm7/VW8e+mhbqIuXJ4E6ogSt+E0
UhB2AZUg5FQvooysc8YY4ApibtypLJAQd9BYKFOvRRfA0yvCtKIwOVl0Xizm8U6oXxnlJJoL5KPY
2IGo5tJUDVRu+YhwLdWr2yCoLZNFXQ5ju7wa6niA7R6bpzzRers6wAoBkfN1ASGZBGJ+NCY/YuE9
7uRLdE5Za+8RAjqi4bN4cFkjThlNY715XSBotMvofRBlN1QKd7vvc31lqAMjxF4lFkqdbM7C5JqN
pcJzSUTIE6mB0qImn2Zf1LVhrwrkqqz34YuCli5IMqJ7aBnQWyhxB/+P0PpMi9sO8apr/Rd2l5oV
lVYl2xvR6FCYWfoSZ04p/3C2ghVa/+LwcLawfQ0It+Gk4QWWam0tzridbT4c5uQCTiG1zuwAWB7i
CWBRYht88vKGsA33SSFOeAXw3ItzHjRqC+D34IDeLtR0uxQnOqGtT4dg9cpkyiT8ubF5uSGvUxqi
Aft72EjEFeCtfUEeMzkcUMSAfw6h4z99kqakXf1JsIJsMYvoJCcUJ4DMiAj2FOK7Sxom6akDOA1G
kDvVXpPdS7KVMhBaUzzy+NUaCpkCdFsAkOOi8pq5uhChKjYuoooxyZufUMUezn00DIHD1SH/IEBL
vJtEvGWIf9olN0FAhoNEEXgles+McXPqea5xlI83V3sDeX+m4pTrK1bVpJAipTTNGXmADGelnBSV
bdR9toSjdmWCthEjWcLOgd/TVuJrfRd+hFSsAsLBh84Cxwfigfmfz1Lu++o+fw4/BEIOSIp5F8XL
IzyPQAwOmo2+qF801TZPteYTc0klwD9JHoL5W6lmmtxPBPa3uCt2SdUT4gmR1bn4NbvftcY1Mzfb
c5OEgiKwMR1jREyMDh8liIYGM5ryQ18YgSOjpNCsFp/5B9rH3WcCbFAO4MqtuxxmSI929sfDnOKq
fXTIf55aRzIWefmi6JwZGjYf6xcv5LYdVABqRgsmsMZReeNtwu4vhyWdfcYHixKOTQBDVwTfPTOX
SsymH3wPCOLEK4f/E8pKwIh1/fblbpo7kEy7SRjP2TSOHhMyibPYLwVVQac3v92QPlP2HEJUJysP
/tx1mVGHpgZZ3GV/htrbGzoEWzcXFfeBjp3kdX1hiVGt7cW/Ic2G7eBLBYcHT9i8DreeOOWrlKNP
O9YjPhjWroDck4TOIwTAw2io7quYA1zAvQSMjqFeuIYEXrMY4AmU0U938kLDPgX3Ca7wsApFyiJk
PjHErq8zAHCNEEUfk/JhhYS7HCAKnBuGEcvpe9OAn/5YwR5iC3m4X/WIz9y990hZSVPHz/zDjufA
dwYFPHPjwdfYpPUId/Qn902gyDT9uLoxaQqqpLhGm7+y60GU7Scw8t9tRy/HfPmkZuI0mVFoH7yN
OJ7LSXtbSGfZNtVLLZTsJBdWglJIiTXKKbYksGubKB9+BS6S4CYZtLEL0EXUjjEoI8owBimf5tqM
Uxe0dKv5G5JH5Ly86B6g8vsKWFCt7SNRQDbV/+W3IYJy7PZvSIh6iICIwNm+913tgM8FFQ7VbUWR
6O2i7FvdBStFA77mM4ua0wuS5vxkou7XgKUzK3knsICwhmLLWRf0SNnt70KoEvbjGzeHYe8rDTb1
tCDzzn9Un9PSyrdUP3RoezkE0odhEVtjklnj7HS/o9ZZ+Xt4fdkjQemYhcJ29ipqEDCD0AUwckCB
0xrPH8RDmcyIcgP6XMkDDUt8VshqX2qvDAT9+gs5/Kny6/BrHAqH6qRpF4NZHGTyD+rZC1r8Z7QO
TWnL4oc3L0vIr6DFW1839JCoPsd1p6pD4yJnJx+mdihCwM/bxl88O/NsenSSv0iWJAZPi3N0ESfI
/sO2ceZDHNdd5aWIfZab/hS6Or5/+rG8I+yvlkhoywpzSOZ30zfKxDmpBORqAxungIbJG5Ep9VU9
1htuLqWiNsVXdRWESGHIqaz04nP0i40wMaJAFpaBuDk2rjRH2TETIQxA1SfjC0T+SL76JWHMZdZm
8Ycmcs0tjsQuqnDh0hE5QTO1iRtsbemOgSTvvO7rAOPFqaZBjcwEx/2T3OBqCKRVHQmnKkQlrAFe
zff+yjKRDzYDDygUIK5Y3T/lpXxj+gRWC0sTIInk74PmB3KW4t3sljYL3uj1LialNgRt41wSCCiL
VbYBFPkf95YZzhw56jlr6othy5fQ7/SsE3PnIjcKM9vtf4XG76cnnKtynFYGLGdNxBoUxdYK2cvj
tIacBVJj4o9CJVw2zVh6p6IWMOwJoXKCjWNAXGCNIu3Mn/FdfdEPwHnjuJNdIqcDX3KQe6oPtMPH
PlbM+X7WRG2F1ES8iVSsCTIScNmEPxLrdJILPRG42UQ+6CwsTkZZbq2zRkJZc9iUlZJluMNTtvV8
abeKgLJCixbQuqr0N6+H5EWEm0CCAIaqla9CfQmrlUtkIrfTH+orkrov+Jew9nv/v2zBT6rZn7LH
zXq29GhYYJFylk5E2n6iy676jEaxJCCqPVZWnhCjMl9RHxfKpNAkqUoUdhzP15sFLQdZyl0ricPv
GY+XF3AiSFweRYKh84iFOBPBRjjvC6S2BnQGmNJIl62cbRnuvOzv5asEAI2Mo2cPnpB1+1Z8X0sh
H6QxvgCeBcaDs7ql+OG+4ZYOnzMUvhDDvFX4pRH59bePiVMFbzAlZJjkQ+IY4Tfrk8ztkUSO2zaY
qDATvUHu1XYmkKzAdTk6a9h23l6DDH2571vhrR+DjDmkfT5+2Uw7GohVzIz2aopD3XruxzxwRQC3
/0NB+muoPwBc4ACIMoutdfOGSRD+ODwWJJTeup7j3ZCLMjLz8x9ogKvgApolP0GhYQrFPrx9uSUq
MXiH7h3Kmcfv092Tp/fuM2mZDfTZfQNWaYCn1I6eVl2YhrT0kcTh6HE/qk1MGyQn0hD7lO7yD46V
HhWQ1mvl102hiiTdD2PUaGaxGu8iIZnspzIEiIiuIM+EvNRbPsKP44rHFvrpPjrXy3XQVgubW7Vp
x+Phoe0bdVN6aTDZHwF2PhbM8R5zUD7Qr88zoszRU1epLGy9ee8zuhnixvulaGxQ3yqRgWxab93B
T152bTerlBnDqdQr4iF+hCJz2+qLgoZv3myn4CSVP+cihfTXuwg1hF8zmD/uoeMtKit7uWk0L/4c
T9NRz/XB0fmbWyIxNTPbOMbLI8yjgvx2ekUQqQYa/Yd23S1Zj6DBFT2cLzPKNrFogGSXMcqWzyY4
ryoNo2wkN/QueHJGbWHa72MEWsZf2hK5MUU8qJYZKmud01WogQd+pX75Fvg6CS1w8r8H2piO5fgq
k9Ay6s66feRwYXB/chLHAfq4+UgnP+rOfYC29E43d5gMgaP9HbYYT4+UC7tmrouuztannPXx2Buz
H6dzlAcdZnUoVJakWW2lts5finWjvWIpEyFdzNz+pyQOAIGUYs24MQ4p2vAj3Y3RStjHAdtPFI4S
9GuLIxCeh3aRrzwyB5j5/8iyQ2t/veGfJ3Nq2IFgiaIG2zIfw1WwaFP4Fu3wAAS5zTxJMM+tSXEp
QYwZnhQjA8M0QNf+4e+KfT3pWTfVMkGcwMGZVR0Ui/kWhgfb7U+E6Gzr0Yo1oI0fH64cwrIi4VWH
+f5BLkUGp7j78Uyw/YvTSYGsUmVjoYgLcfPlAic6p8j0nam5gFo2tJF35FCbli3hm71n8Dy1+Zyn
n6rkSjSBQSlWAHHFjarhusM8xvlHNI325rcz1HleyNf9aF+SgPQnpb7h4VEmAU6Om7j+VVKnTesj
bu/eUeTARJgoKvr0eeW6Qp6rlxydYe+KFe6blY3HScICrXBbRbDRIYuU2ADoshrW7ETh4W2BVgj7
Hv7k61FIwKgfd8Yn6o29/IcrGDhp6bA56gZEXR0NC3MU6v+eghJRzONNSdG8UB5arNu36kzWMtI3
NBVZOnbUNCJFw4Q7LT0iwftveQgQFTH4pJAfl0iVFnq9xV09mf5B3RK3N8C+4LRE570074noQfi6
TqRmBKuVP7+raRuaQQtL5I5EkvCt76Y9i8hdMDf28f9y88LvaAKv0ZQZ9YX9ea4k0TMA0r8zbX1H
qxkvtJnF+ihwUW1W7hX3dxq2jrblOVjol0DA7CRR5QMDQcaepQFy+NPtYskV2nXaE2OERZos52wT
MQ3Xwx+xmPtdZQY8NpTiGs9AvGFZ2n9XKAXIBuQ4utFyOQOA+BcdAfs8d4TCpP43BW6B/u4+PGMe
1YFncCi8Ulu59CADS4ObV8xxO5BHT0N3NJoc8zcrG/LNPwc7yicDfi0JuKHULTPVaTFDw/SUi252
OvbT72Ao+tT9MvYs5hraze0b5ZJ6E4aBEKcfZPe3wRBTcpN1KuUxDwvJ+66nUEm7RcWsEJdfqM9X
Po+rFa1jTHRwvvv7sLZxOSJWdRjZIlFpP9ovMHsYPwBWeoEpw+sTvFutxawX/QSvLTYpv/DMEN7R
e2sThrpnL2EO8q3Du99sbZHceo/iyFz4cL/9hpvqG5q4lq+JXpS+K0NBW7OM+zCBlTQVp/1s45Pp
5J/sbAamJvascXUfEYgCVw9wmpM7xVAq4js/ffBfyzvwE3R0PVQUr11MVbMohYuh4WItbUXCyHlt
x3Ipv15xWvceCXbViIT1Zy7HApPPPiFRK7M+Nodu7pak6DxIGNFkpOBxrc1gU1PvahgbIGLaSUBd
APuHaGzU2hVgTtDRiFlA1xZuUMo2f7BtiTmBS7cpU26fHuX3z+BQXbGfAl1b7O2dmOUBdFJWjFhG
eRzqJFlTeYc5tdshwm+L48kFetJf9hPk+21hSZ+nfiNk8n5n+c11nkS0r9r8quqmGVvaVk0UR5tD
r2AzkdoI9I7OdsH/MRvxcnbesOikinAHDmw5TPyOpCEuk7za9k+whkLLqaUisTZY81EMSpYckIyL
MTxlnpHUlplxrabjyv7yCkeYM8IJ2/o7ogkUNTdX1XQqDPBT+KPFmpUyOFy/ENbNZG3YP24nJ0Wi
451g/4AiId55nZBJkmnHDWPQejITvem8eQzBUIe3V3vzK/TtnsnseFHe+4KZtFT1YRKo31tWvo34
D2C/yiu4kHS1aiRUnAGvVgOeVTtZD6hOfVuFDPIz3aof6q9nTN8OcRJB9PfsXemss5P64BCPdYPQ
snPDGHUi2FiScy8LybGECJwGmWrkWbcTatWjoCdrSJTUVflAXaSKcrTqFZE0R1QOAMEUkrP8sG7F
30lmHPuzyglJH53K3LsHh0DRMorhVPSOIt8cvq5xkC/BMYYkNG0VVLA9FHaAgIEeXptZWNlN/xdf
8iOFp9WGWzHhO6JFe3zzLarAjujnQauQ79q2gHnFWlOD2zHO8gAMGH0sSA5BWPmtfhohEjgogB0e
axzVyyCsMhe9WQe6aG5J+QMWkAECGSNWTYjlMvgH+VZj9TZvRt6X3geOE6+bwMRdvrWIhefsJrB9
pRfbeGF6D76dTtYyr2Oxv/hp+JTglyOjSHZ3XVxR2/N4Vyb5HHRpXSWsU7p8WNa50R3cjOvFju8N
jWm3lDeCNiDK0vQhZ9IieRSyK27/f5C4n8XBaxrztPf8goVRaDFCPAd8aa7e1/R1Kx8aEhl52S/o
bdxGxCzM5mvlzrSSHQJ7mk5klF5Ln1PglPuIW4LwYZbEcGJG8zaoV7vokPVx/DbQjeODJ80f5Hzo
KMZjoQ6wN9FMSU6GzYhx2Jp30rGYCu7WeFdUYAiNpYuzB5ymrCStp0wL55oMXngwnDFsp2ScPv7S
EwtUa7HEhvCg6+VNviLeCEqo4P4A6dNvKe3IH/6Ntm74VK0JBizcfm1abOb0ulVKlDX5RgVJfN0A
JWUIYGopEDWUQkIwTZc43KW6TGcafnQNK22FxtrwP+6ICchKJHbJv9bXoiJWyys0RYiTsZH5PzUk
CCXIMcmzdXLOXkLb25pmB4klRvvTVDFrbn8byMPxqoUCWJ9Z+2eGM+p8EfQA+6XW+0KgxNO2sdYR
JjjnwnRaDWt+L/rh6xersNwXXx+UKE4y9wZAU3Qu/mRRUSLrXPdWFUFxHnwV2v5bsRjT+mryrNON
4B+3u0aGiRtVrjutbLCj1IGhNPCxCttlRLOfi4M0yJW1T4CcMb8OGuDjJxH7CN4j/J6nupCBEQrq
YtS4neuNEFUF9sVj0gTa7cbWA3pE/IOIn6GkTVlgKKJI2p4W+5knl+wOSKVKkwAA3ByX50rB8972
mxgkzQvCo3ANshsq2BdqX8taydZAxwBK/5DzaHmAnkRJgKX4eLo7S1Z6LtWve/7/EJVNWKSfL0Jj
EAMaEou/sM2ppX+U372MJtRlykSbUNxibTuI9xqNg0iz+EOkJ1SZWb79zljTcGHXaMBDhDDmwkw8
Yz7WSE1LlYt72z2a5lLp14KECt1X+UEiiguXH/4y5Nmg6yEwPx1ouA7loSYJIQFYGB+oSq6bFdHI
9aVg7Lrw5egpBYrsbFY2dpwmVsdLqoPTmpe7AJopcSwxyZW1DFaPpHuLWAVa1SpATr3dlwx7eDtg
2K8wQhnXpN6f5LUjoQ0ia5swQhzIIjyJDeWZ3Q4urZK9HoBZjHC66HU9DBwUq16cbtrpWEm3GNo0
gvmumnd3xatsRgxelpOUhQxqPIgQ1+IRB3xDuINZFFaqQqq6jcFYWCgIW1bPBITG9evwK+Hpa2D2
LJ416PneY5XAYoIwBxb5Yt0jxCGk02Eq/lSe+A8VS5+sk0uR40bnbzKOCWuUojshgypWXf95QnO4
rMQMymKjRNTAbYmWmBxL+kA5MwV5tapcxfn9gk2vzS2gkh9o9oTaPzOxTVLeuVCIiPU2rSxHlU8j
cJZ57guuJTUZMA1Kb2BHeC5EoOxW8Ln+Ynsof4Ho6O5FXawwhAbIB5hG9EHXLDALEPHGTh6iIgbi
3pEbpwG6pk1UMIbpObMQ3u5xM00zVyCVPGR9r3peIXXBnY4vrDSwZr5XbLxgwYd1nRCs4z3B7RG4
BcgyIW6dq6zBr+4EvX9cStJhnWV1gXkXmGHtpcXYVaJd+GY1QFG/KswgwnX2tSNEnKOgYCA5x54F
X3DALLcbHG1iC1OOvQ18yuUDFDRYzZNu5YaPvgzXXd+l2WPBMVjlg/BiuGGqXmf4y6/OILNlbBvc
1FnOY9ySr1MnLLDvD+5UcIo9stzzM1u1QWbt2g7NuqIkLCnjTqz0uZQ9nWvXGbk0UZZgpjBwJdiZ
EkQ6YDt6XcU++GcR0TRVorMYb46KUOQR3Iccn81O10cKR/xEXKJbTnOOVjgEXDak+gh7CQh4UBip
vR+d0CP/Cg7e2RPZ0h3PTvzU6rq0/KifxsGEccb1RP5oHW/wymSN9gjdWCzSTtlTbPe7DRvwu7JG
kBcPJzNsNUfi+2cRrUG0qIlIZrb4+FyKXwe4eY6E/rZzx6CiRvxrOC8T4XSSpnwwUWC4Px/qFQ9I
9mPHnmvR6nJtJCtUKd2hmccZQYaPr94iq1AH89E7r8v71e+Ekeud1okg/KAYVtbsYSR6WxPlroqW
VHWN4k1l0QTKhO2E98iAiv9lwsLEvd63P9CHbu8hz0ZQ2k8K5ezvi2H6yVvyLbPYO0vwbnjqyEef
7oB7kZh6Pjt4OnMvri6+QXG2tM+nPwQ6oWAxqvOGFTfjw/xnCL6KhArgO8fpkqdGpJTeZbxdiH/m
DSIpi05F1onSOW2RxNHWSOo7JX2BV7hxtOBABfKVM8GD+BuR5+SiRXG+xnTlJM7VIEsEwbpp2iPM
3Zxdt1DwLIlIBGJYrn3o0HK5SMv56Bvd+PK51hh0mr8RqfMSQLMySkMQT1sAzWbsSeTYj2lf3Xn9
h/QxvEg9mtgNUNNdZxwe05aLAD6goL3h4qN41EX6x+/IlnVfZcWKeiBjJPj/JePcKLqf/vTamB0j
+cGaeF1cU/dJuZb7B3oeoMzJds1fbE03qw2zl8AlTlW0oER30+XfHfIuACYAlwMlcCJrNuGu0qCu
RTKFIRf6efis2d5zBI9rDM8+xA7LYjpKx+SuUCaOai+wv6noQ6N/FI0RU4u71lUjCC+UHMDUNfiI
7BdIp4aCxKIkmBWS5FGfWgwND3nFS4CRnRzC40RrlzOW33pU1bXh7LQvqsZmgD1ZdlOqMhsDGXXP
z9lBylCkLeOUc2pNmEVYZr3w3/zV3h6Q8ayualKcJDusS7jfOZaoZpCzNEHkDJD7B9zHHKDkaejU
0Bu6g0qF9KjwIBaNnV7lMQN6EE3HvmSNqJr+r5iCjYAd17GN133JddnhcSHogMqjaVed1rECpc1W
j0y533N1MaRN9WtyFFBlyO8HhnLFOLyTqp145ao2FduFd7bId7EW9AlhjQUFJ4FWIGaa966Afnzt
115oB63/DpQ8Uxa7d4I1lE+FbrFuZA9URGFowed9ee4Y4AtEY2Tzas3GwbAPgIufdwh4Y98iyLbC
4mCFjMthUMbSM3WDnap+CTWhfyXZ+9YJgEGzoLXBSqY/zfReuBLhSRUiyEAbLLjgAEorWNTWeWGW
9UGtiTNdZIQRkPccYcKkWRLSpBBoJoIeTPeGAJVNvO1f9DYLAJr91NwlDiwkvXpwlUiiDwFIe6g5
9+c1jAkrrmw8g4ubra5x4amLumnjfM0Z2nAvrkJlLeHDm9qexMIRXILwU/tVXs1BB1OQ8enD4QRI
/SLdwLFnZN3760kL64LFGevPvZQdn4RCYBcTT/uya/7UyfMdjOFxK1khqYYrMLRFT0U8YXeTpS0k
wuVZSiaF3hmGmU859ubu/zv8JfWqWkfSCvPb6zkujCqAdKYNr/+BNWW5oj1f6oB9QmMLSG8yP7Mi
yalEOiGr7JZauYqpxp40Hlw66wXeO0kRi6441oHoWkbnsuRfD8hjMUGZ8QJawLKE5wbX/DUh4TEF
mL3Xi240XyCaj5dHZSjL7lw7vCdq+PgwqIt3fEx2Ost/JlpguDPbDu2Qp/PLgR/mzgxMsykONDnG
qKGadiZIu2AW4eoDPwugBLFnnVY3F6UJvnnl+1r0FdnjnamsFN2riegToUGTByJGkvAGxjwjA1Jr
xCCujT0YkfF8DzZ4ktR82pGlH6BkHk/3brADywjbUaIB7QgOCPFB3/n0nS+NK4Y3KSWjT8nXmyMR
g+JB6vN0axQt+Jpd+JKC1Yhh2JyTdg9hnI0e2znCksQWqW/rNQzrYYXKrvGiM6MrA0Kk3SvfxodV
Jt/PjZsPBmPyz/niKNeFRNzQvJrh7179ivVLrygcCGC978MkSTDqsolob4kBlPqK1Ge7G0gs0s6d
IubWh0TbTVxmf9XvbfryFHEMaMBNjKuDO2Js0mpHJd+baHPONo71Kz9Lf5Nk+UHDtCTh1TbqxrA6
vvBkVk8oyomfT0SGMXZzfJv30kxUrKXJUSbIXFo5A183f8lu2pS7A61RBCcPXPOw8kBHFGl05vAj
oLubGwbXaU8Ppwrh7XTb26HOW251kxALetvVGE5MwL7IqtJDot0SADw329kSd+J3Z+7dQEgf44sh
KbWQGnJUB7Z89zWyIkWQ1foIKsz2AJWHmogqT/hMgZPsy3oz8SBcWobC22ATicAvQmv7PR7Uv2Nf
O2+Z5n6EWvWmXPNp/G3OZsOViKj6lmmyoTb0AddF50LvMpFLENfzMCZ4s8qW/h3c8oxloLBW0+az
hEj2g4o/0GbYXArzh6xmA5tjG0LgnD91nQojrkhFNYnS9MpHcoIg43PEsxhwhKxQc6kj5vQ5Gus2
p95ViNrqVy28qwJ2gYMNyINNFyyzAOFM8eDZWIKF4DF+hntyTALoSSRMgDuJEH+oE3ejQjtVaPOs
95TL4pFCTMXlfVm0UpwBk5TCeE64joxoGEHcVfvQ2mw6adSVCOXMBrkOeYcVM3Pazwta7R/ctYZy
8NlvYowTSQlQpGjToGbTkTmnMddSWcH7rTV71Wy8NAytSKnbmzDIS0UKckPMYcFUCJFk8cbxrZxI
4W6WLw9u1cKlTj4dP/lUHUvUAoFen54JCVWci8AfWaqJGuMxuOcpMbdtyC7O8kSU35/s+UtQrGll
ZGPEiTHGxWKCzRBesHY5RVmpMuO9ecyTizfggR5Znavx9U8NSlwWFIpb4d7a/bZb793eEPjwJyxi
dMIaPZsy8FdCa9pIRvmZi9SgUL0zs5/8G4aIkueAZwvWXQUQA1Pb51jdmPyUbApHXFukopJjaTPw
No+n0Fuw2yWyT5Uggi+Cos1MsHO8YoxIvk8yyU0Gj9w5+FM4p2HftSz5zqUsuLv2qn511T/6GvO7
j+Nxq8p1DY3EgppnIz9ECUS1fEky6REm3M7zt2gyIItySsSYT2QITwVEr8gXfWZpsWGXo8NSC9sN
S/SsDpXA2Bnxeh10lpqODzpjxG+kTPUXsPinbX5/VLbYMiVv9OTwmVOhvmEvU7g2ng5XoGtQRzW9
A4Fb5BDEklFVQLy3iCdHZSRWmUoOOt7yr21OPp/HNwuVj11rx581AmpLtstRe9u/EG/8H1n70Yar
hTpcK/lzKEGzAPFegr3/DzQOqIUy/wHNS3h/+zhUJmemdmgrfO0nHJPwFx6cnONl5j7Jwbcbry0J
67fowZDAV1SQrv21fWjE4lkPzIKWqm3ImhvdEmU9gRSkIKPRM9bVUiHJqXTaoTnTknOOZaVZjUbM
DE2+3su+RmSsYdiBlSxVPj5Pr34PGoWqaMCUhk34ao8y4FgQjAkmD/vAi1GxPjJlyAxBv7Sp4rOE
pw7fONheT0Qrp8vpDWZm/Q7UsTMJ9pFxH6KBF2K95oa/VhUFlLDwv+f2hj/fVDwyv0puBIKWJw8B
Hk4F762PDGiIvPVGTloJW2H5vZMhEH9ubE++6hMcSsNCyzapbv+xBK6lfHfP+m4JaZyBrvL1wkPa
/8Lxh9HcHSjQVcV0BBXGD6CZmjczf11bEnZz7OvR5e0qM7w1mwkQS3U2mXr1gXjWYkIsly7jaleC
qdRQ32sbkD7rThnsuTkXd51pbZcIl3HWkA1KsXMH3ubnn5BTDrCTlgLDKQjL2ynvFBfVFjx+tbIs
CUTUxF01ew12QnGTyxHwp4xYsFsgY9BPTdvHDbiTSJGzZpH5w/an5hUR9KBRDob1eG7Dq0oaGE/m
EttHpZYgGvOGoKeRnk/LddeTxdsFa39nMW0u30R5qwAx7Atdig0DXJeahXPnvt+0eYcqgohGD1Gp
+x0umbzP0vdYMIirAvJCx6wee4CRnOzSHb/mAJ1RVV87gh6c1ntueXT1R31zjl7TlumyoXk11ICC
eF2Ph3429jpdmKLH09MjK9U9/C05FoZJDZAr6slBX2ZWVGVf86mdhzcAViTihpQ2ZCeA6w/e0kIA
VlPs1GOqv4VetNW+4GO9RqYMb257XWkU8GOlHrB6ufo7Kyl+jWGBo5BvZLrcBvrM3MQ9c6yT/PNY
59dHOCPIP3Lt9j5M9V1ERXQ0w2IV+bYkS+U4TtpwvD9zGrhzB5zxNz2pIxxgJKD2qTWXpeiITGvD
wZFHhLcLjg57CQ/fdMFf/6DGVNiAD16aMWIwhgWAs7SqsDpMNVam2vhV6JxyydJLcov7IXm7XL9m
KUNbFnBVnpHjySuoiQLv+XOQu5EWs9vtaOxtQzp50fS7W1t3Q64mEvg/CbLwXsqX8N9cKC1C6dPB
AE5m/np3F9lU6NU0a9I/lZl+EC1HXwO605kYvnFhjChzsGU613wvZJXtOPQPJ5GzWVTSleyU0qIK
fLmblgkRMJsK6SHfgEq7vXOUZ3yPvdzb6KR6fv9ylhmsL3VbO4FPMllW7fUwY+wu6Zb5DhJjoT5x
p4mlpKQppGN9C+vv4kHrIfZ/lYj9Og1pgP8t4CHKmnDfPewMT9VrAAd3pASxvhbh/vHN3lR7tIH1
gJf8P4Cim4qhO8vgH8Rol/dS0tq1GpcyLTjfElP8T4W9V4IDUjZh5Ts+ZUHc4DvOJj+sqOg/AAW4
X/+VpLB6U2d2tXye2OSA7VsCO//QMd7BPCidprUG6OsWqTqZR+qwVwzZGPEiSVrhKT7dtxM+6MU4
7+N5S7t/e/MXTfVtsO8Lz6kSfqgOQKNUIQNdMQ0r3eNSMPwwqlx2j6SEcV3ex51uhOB4XPuXa8Z6
qUmJDLNjzYBLWVEhmRT69Jj3X9r0o7qK7CjPdky+qp/cF6rseJNE0vARdroPLOPH2GtiA2eNCMXQ
drJaXDFXgZG3vOGH+5ZAf5BrRQJEY+URD2tZHf7UFhLYc6DIABViU17MEpByQjRBamNYeRiI9LSW
Deej3ut5+mqIpiZvdwzCMDd+3A19Z0GgZxDDENjSwxvra/8QTZs/XtGBYB8YD0BKYi+3Q/aCKkQ2
F96zr/VV0S1CgS9N29sf5dDcf62iHQy+8nTa19Xzlyg4uPe/0efIDNxs13keQOHlvJVh42A2oFk4
28BuweX6I13WP9c8ebvxxIYIZ83DPYqDXW6MHB9zgsC0/jEHtHwfLwIQWa5b9hbwfiMatYQmmdcQ
YxXJlEKkxG5WeK1add21NmpfUR/zK1hexvYVT7xK0pccYGSVQ+1HVAN1Cd9b9BT4XOsVXYxyzqk1
D6zpF6NgtLjpPHgLfreJsmcZJcP2Zcw8+yoZxLCH/SOzze/mGg5+JqCZqgeF/4NsVRvGl4UiMfms
qvj62YuSjFlEQvnCXwhx2u3QkOEDMajCjQnDJp04haEuS8eQRYVH4g5P+MuvMt3mnAWx3ZfQV+c2
MN1gE0GR7OM+iRBgThkwlyaPqPhWnXN3xWW8PBY/l/ohSXxFCEFqzmMvAF4hiAhtIvbzSzicM/dI
FXtOouKPBhqVxupP+AMOE+fTT52qUW0eWKa4BZzcxzggUJTc7TdwB1W6t/oIkDl6hGbtXBBH8zbC
fdFGL4ogSONYdPVvfL8n8wvq9sRx1P97bMd7V9+jxXQ2Q//FJVZwNyp1mPv6UJwzaDLcgISrYp1M
xBIzQoIg6iSG405P8pK8w5tsR7uEA5YLf2ynYSDBVHTFnXQDru1RG8ji0scKtETT9Vq3Zcgk7x7P
UToGUaugMEVdeB7gDbPb6ljwWwT6YlDjfcMQx1zDZmwNx5+4/Dk/btdGxgnVD992OpKs2KyS1hsN
YnAOW/AV9KSX3nIt2pZZCcWnGpOnkJ3vaOGX4ZbracPzP5wtXKksd/P5xwXoO2qHHOK/jnEdPs3x
RRfRQQjr7irBrRRHwMX9gaa1v7m8FP9psbDS91+3y8xGeQmUAORe6b9/A7xbHHTV2BcC54t6/Avi
xujpKyFqjJg6xk1EFP48AqZ45Mw5XS3/lsirXwXdCIis+QsSPRwBnOp1OibYtxFe9QafNzkmZaps
eQ/h/qWh2/cRXQzEuVcqBgcEjfW1WxWRJukI0qoHaRcCknI4oe+CZrNh1q5LtwMqbaU23rTmsz8M
IpcAN5MpTmRZHCrGpIEEWOxQWjH+KMnuivSg4wRvDG7s3Gv7eGQ0sHahQC1lHgjv6ZJxEYJDRJ4g
VzHtBExJDSOde9/kE8J9spGj16VPoDGjzN+LOJ2DxPZ05a7uv/aj+bdhqDXy8TVIW2i9c/u1KLZB
HOlP12GM9PjPSzkcWVdqooQ017tTAXKJLUGPj6cMrRBzPQBqGwsEERrVCt26LIU4iciJxMv4B/be
RUfa1L9Uwz/21/oOFn7+7dg4fKj1mKF32jC2zNyJbIU7I20FHm8zQvKjjr0G5X1iSm66v9k0VAhY
h5fAZBKSAx6+NIz4a8IXu6Q+JTlBaNF0ynkzlA3+A93ykpW1gPeJI7BMynXcw5x5lCzxE8C06VT0
fhOKd87YAcKYg3gC8Eq/8HoNqt1/HWgZFYCHF/X31067E7nJWf2Y+ilLvIIABfdDIxubC6zTaP8s
y5Y6K1FP7eElNd5UDVUz8DJAZqkPRYiH2NwYDDodXI2/wsQi8mX9kd/n66ZobbYsymZTsNhj3d/s
RQA5mT52Rx5LT98G/HIzMsQY4IGB8YI+PffGnFjo5w/17exJ9h/HdlLrJ/Oybm1QOj27FpLkrAB2
vTPFOWzAq8Dqpaf90rZhQFnO7htlAWWrilXyOsojMDEM5EtmIVPMZixLAJXorISw2wlZW8nXwUbS
XcEPBIw6wBMWIO18gmCrHbg+n57FCYk8f8RUT4ERhK36RTt+2MIURqkovXtQYTY/8v0f0qH50oBF
CmABp6qh1Vy6D4ok6gBNST8fe8I9uhsFKBQ+Iv3QH4YbJUtQI1DoENI6bZKGiL5YOiXjzU5z//yC
fz101u3gmQK3dehI+UnA94+J2N6gKnK7IUjpDN4SU+cfsegL8jDN2gyAuodJpf/qd1WBCS7S7ddC
J4CHLmmfM4m5llPuqPeOQdl29P+RMcg6fgocNXR1xeoeO5zCgbOGFaCzI1vMR4TWSX5Ay8RB3GuC
kSiwATvENxI4g4AqAQ1OVSqdgKNoARjpr9wBBFvIXv2Q4AJoYkVh4OZ9GI8C3aREJLw3Br/xl2Il
lineT04cTlRBeWTpZnkI1Xqr0nqc8pvpAXrBRnI6pI1mXdmeD3YSj791vXTnPK1+5ga5X7YsSfKx
qL2CAqyXL3aV+rznZiY5c1Fw2eosAR2c1DuESrdvCtQrUPOMWkQpctZ7U8eqf/4ZmDSNUk8uWt6C
2BrhvrQp1rzG2dXzLsZkP3zgwjygY/3+IOyUswj5YjmuDYfFaIko1UcnyQ7S9djiVGQc2bCMF3CY
STENxuQ/Ro0abHMan8x0ljz+SfGjqmBDf70t53l0OOit2onLw3H8xQidTsM4G1sXX7SC3oLAjN5T
ZEHSOp7/qHoJuVeiV0fUwx6EQ/9eBtdNNnPlJWNvJj3LsmDjYUehmNUjvBuCOS//RoV09mjhbO7+
oVJS+JZO9o/EhvCgYKqLW6+BCWMwRzqZniEOl7USN0R4f/rKY/pz1IqUQCwxOXDJ3H26bpkWuFRL
HYNKOHUx471VzOO7uFPHy6BrGsFbt1kC0lmC9RlNtQOgQX80+OgK6qFdPXf0tpfcidO1YHZsYgcN
TDcQFTZkisqgkCys37tHtck31cj1w6sabS97Ka9bX0KoCkpmJh+Q+cXzi7WU12AbDeYH4exxO/Tc
day/82Va0VfJDWJiESTbwmU8Mam3vaaPaji+Qnd/OHBTvICTNYNECezB9WFzvqttiKn8zHkqOgKg
PxOKKk13lOJ6ZDgxEYocecs9ZFsbkEwj8cSAEWL9XKgfAj+BRJUUsZAMBT+BI6dwSXb4g7wYcwdq
TOH4hSfMWnG9yWFmPmEw5lVLn6yLp7jbgOpH9xAPIXt6OdwkLZ2WE2r2eJn7+P8nHf97l0xa08Sr
rI4V0CLMSuY3iLfKHGBma4zvEqDo7mMDdbhGHmO1nQO7DvGDWYzTaJoDkBF0fNKHAAhk6rVG5a8c
IFsrSil8waQqEawOQJjDPm8pzRt6sUKRK3xdmCccQiYzIFOgc+pnijiOEe7mcUa9T+pRxuquskPP
iiFdo+6RdY+C5Q6i9n9bX0tlZRaKf3uuRBARvhchVIa6IK/0UZutuuMcB9kl6+WOir/OC+cRe4E2
5JpQRQt6XQeUldYhtLb/yoDnckGiiaKq3Olh0bQQdRw2m9BN8ivD/n61Pf5Y2UamACpKzTGW3rY6
wka23jd/TEffEFaTNGXEDeiRwWv+JUNYN7+FyPpwx4KZxZfQbrPffMggtirGdGE3BOeQMVeWDdec
QzBJmy4YNIkuy6HGWaE6408CZ47O4YFupA8BOTuIzYT98GUPBZjbtXogY1GV8ovXpQMTFlqT/sQd
SHixotPAhFwg9JJ9T2h1oGll2Lwcp+8DEnEcel1a2LbH/GAnJo6oBSZDRiXOvTiCxoX/fW8iHfbu
HNW3eTlk4b3/7BzN2Xv1jimqU2YknbVCplvhSE1T5/7kWOmobsB/i8DG2K+klE+HqWLyLddHdlDJ
7L3oZwN1jyIjp3tNgHMNMvJY42j0//L0+YLbrWGU/oqPebPutF3uzXuwDpM0semIBYovx7x6XOJL
l9jbJbJpRvliu56AHiBpauG1EwfgvcSDwboc/0LM4e0Lw3TYjTFLkVFaqvD0POWUdzh4CaJnJg7/
P9/flkUDOCr4+eOt9dMl2+NhEAH2yVZePhKV/wF1veeEYrOnPG9xpPlLIxROiqjuokXsgdGLnFpm
bHuNzywSYsJsOCxkfRZDbrYb1PDrT1sx9mfskXo+U03uggU0Yz7wCmoKTZO7bzO18LpZ1X93aDI3
HKjbj83SJmjdhjFh+RLul7+ShXkonF6YIyNy/lGdoui//VO65Pqkstu9lHWv+Fjlv0lYZATwb7E/
fqIxwo/PymGCDEW9xGiiqTeOsKzoUJd6Zaiw27UWzkni1EwrddRqv0uIibjG9OxapGi8dSbqON+K
4MJflP9e237T1a0MG8P52Ulc7OR5ajsjYhJ4nwazhMGoFH+Pkfll0XnfWNljlAqFwsxoLzXJIolX
zflBORTq7+LVF94BuNzKe9xoxpwqkzjYeotKkZ6asdVttwgnRjrEP/drek4d9nAjIvWJA6+M9ahD
WKu5N/qHsqLMdsLd7YqPEb3htCWT9hY9NJr4sEe6kdFq9LIib0+aKfc5mGbroNMy6XWmu8pTB4uZ
BLUZo00+6SBIe5tNwp8JMM+dV79X0bUS3E2+9Hg5BUJerPZGWD8Eb/tSKMp5DyuOmjo7dOXr2Ran
Mt1Jz/CPYU80uXvpgOCqo9CJiMlvBnqDphu3oyJWkJLbrAwbQ+X24vUjTbzcM9xYaeZIG66L/8Bc
TL28DnMA+TmpfKXMIR5GRromhhb8P368mSejOvdu6JMoIukS9NdsooMTXKzDC5Lng7vjWqGLdjn5
XZcO3GL7DUhyEWpkRNVizfG6J3xBPVPdWzPMWh1qd42GFjdAd5sCHfgdhEVAGE3189aKS1suE8MP
PKToxjcRPVrd9qCdOdcnS4hK+T27EWMN8j5mqcd0RJSEnWtWHyY0xiF6ulQZ4/zy15gTGTsKEGVi
NJdHR0hbYhQZaJUQnfkAs1cTxwvqy2QXgdFdxNP6K6YhtsBsXkBKz3T0crGhB5AZzjxjDBODbGyl
wiHxCIUI4QMC1zvGPom79uAmGcOyVpsho6AW7W5HXoDeXITSSKMZLfjelsm6tHAgo30lXvbNxrFs
GoCC7lPfMrxNTsn/MRbiHEtQtV96ehITKpEZXnnruMWeFJHwTfKv+0wOTpSO8uYWGJ6B8G3prxZg
HJxlUqK28EbOKms0VoUd7BxGF0713NfjTe+rnJB1NJG8O7aR3gHHHyoAxTCS7e6kfHXVzAxWI6Zn
5EZvNfKphI9ATAYWM5UW90cZ4EHcKFutPD5xcXBQnlbf9b06alrPcvDN2n4MUxIydeT2RVA1fnWg
OKuqf1ApWY91KI6NPZR1+xFbn7kUIdBtCqL259jrFHiSyonOdOSYLsWJUE83yx7GpQ4CNFVLC5gl
+Dr45D7wZ48uhsnyixB9hwau4rlA0Mj78bH3K+oRUDLSa7X2lx86h9LHVgpRZEWmr9+spBt0cdVr
MUoRz3H3P0j3yjMHWxqGauQUq1yzDmthiF/jd9jnMAApLLeLoH0tGUq4AfrcbJ4gxlh3Bl3DyL9V
2/FSSc+eYKosLOJ0iLXYKqGwNsWMSN9K8b8wfXAXDspx47Sj2woL/KUSkWeRBGJEcI0uNpKnnIAZ
V44wARURwqwfkk7DQSlHGWH3zQw6suAnvbfHulUCQsm4gDUFp7P5CE0zRmAgatX5B4Jd5g5eRlqP
7EjySrM3qH6kUryFof/rwSATBBLVNTtknrU5D3IX1nJC1s54FNhJIAXoCGbH1LkAYkSJ2pcO76tT
E/phDQcZC3tp1Bq+Kil+hnD9Ifk8L7VR/28kb07uzE82m2B2GfVcl3UCOPWiiKq66n+IsxHRJTDH
Q/G1X+6eZy3mRL5TTJVcmYsSFiLdC3V0dnm49GgXSpdlPdO9J50zBqM3FH/dx1TKdRqH3OB/77Ux
SkI9C4otvt3ZL4geTXmJ5QrfKiC3btlzfnpnv3p0e5mq7dGc4YU8eIgBru61uGDYRismL+7zqSKf
dIRyrqjeuWwCvR4b7JcTfmQfOt6hERSVCNDSXwG930PgwWbLSmqFLE5/HAFdZHZARz/peAaVp5OU
r2PJJrIOhKt8c9zEOXfbY3CNnKXGrKaTQg3O2ei4K9y9qSHhW4z6tXbycCZGTn3XB4O8d156vJMN
8NnDCDvdGyOTA710K5Seh5/Xes2fJsK7rUG5bVbJb2poTOZBFZWnzrjZc9SI5vQcM4xm/2ofkKG1
vGrliHY2SMgjaJLtkJ+5C9M7JcYLRr1zYIQqdeFtkcrabbFn1NK9s5BGO95VlrTIRNv6BxwVjBuZ
OZwYShsdP7WA5xIKqQct13Dk6c+ZhpOLVWfrA3I5Bp/c2KSnqUnJR+3qcXq/5ddjt8adIRoipoTA
eRA6aeOX5Q+UVc1fQm32F69XdZaRVOpDizb1/HdkyJL3NjK2+Gwre7TJHRmc5RZoRro7JlAwzIkE
g2l+SwZfr+khY9lKQ7rR4GGRwOAJpQrNVp131zrusehrXOI7yk9v7JHLWUFIVVollB8cZP941slO
zyv9bSRlm/G9QKn3+9GvCGIcjONOW5a6e41Wx1Px7ONzSGG9h4Nhg3jlJERTrxOmf8hYMPiKt5kF
ikMplbv/I3jrgjB2RyfoT6/HPSpFKtOWuxrMu3MHRHc0pW8tYJsgxzeox8EdVZYjoYZfe/Y6KErK
wCZKrctc/EaxT1cXepF8ymQ8svikNJdkCWFJTpzvKwby4zTtVabCJ6k431tiNEyO0Sgw3iihI/Ga
ULl3BiTAwFvX/rs8WhV3SBEKFxxweqxhMiwEFSLQld7lSDKGW7x5pg8b78BHrzrA7+27MYxrHU+I
ceA5tu9qb9qIXjFYeMRmDT0RTM/pj/sU3zlXeC6GA4fhVLe9tLOfGeumI7KuRT5aK/eV87nPtryE
wDeaCBNv85bypsk+i8sgBrrxeYmMbsesCKRiMKiXY9DBi8HcO12Wh8MKuQVy4QbrHx7Zj7Kiwcsq
XaogLjzsSVt9r9jrk6rz5fjcjiCeMVj89RUl3kUWUjU3nImmQ2KmuMqZ4rIqlv31iERDl7/B2b5U
oHU2/ddvtTsAjR0dwCFQ9Ql5wErCu7oaOpsisq8ymzgt5V0Yu1OKYk4sB0WcaJ3iKeiVn0P7Q7VR
LsOxxtexkSA7fvtI436yuUokaU1NgjB9C5ZjwAuCbadsrBjdrV/P2mFk+MO+wZSuAu9FmLaXQNyD
xi37KSgOko0jlaozfaBbp4W4oQps1BY94cdpPXWQBNkimRUBwIZI4AuC/DPpprCwi9oeI20RpKJz
exuMWgcmRaa19CIuWelizq6/SIi7ezxaTghgXFZDzGAN/Nl11qnQO6MKYDnrGUtkzBuZ7LrcabkF
BHx+ZYKyFa0B73ry0TvVFNAiO/rYCXlgIN0OU/B4P0bwJRQ5wHkq1Sv6Sqp+Kr25h1BGJVKgNkhL
4g/zWekVmTiZCNtrNVyLiKSVlaWL13yKSMhml8ouFpoSIJf4d+n9PJ0jU93w3043/xEOEtCOByj1
XHCBwnXgKYMvA7e3+LF15iLnxEzTs6AblN3brLCJl3MK9q3yVX2zbxpwquttPB2nz1Wjn+VY2Osk
zopTM6IArFnqC5/7x0QuOAxn7fv79/+rqKfxn38OcR2SMH39KFu/womRb79vXzPs7r6PHddCwLU/
aQSCM/jjt+w9I0mtPtluTYzaJif9NgIkPxIW5d693vJinLY+Y1MZ8XaGlKCgYJ47QYq50g64EEPo
4r7sF5dHQ2yfPqbMLuOljJMM9BWg29irlyI4JnyK5CLUr0ZQ981uYx16VeqUYbuIiNkqsrMmHbP4
zdWkQd/B6akiXUk+w7YtwiliXjW3UqjYh5fliwHKdLstRifOIdIAU2m7ze6yR+8wgZ91aXt7Tseg
TpH8U8N2D+iisQ+i/OlMj6O72BcnZz/aplvv/N0bQPXn6mOOvzYYqu8vhNCM1f7ToMqQcT4qDDou
y03WNqlgMx33p3p1mIzmwS2EAZNSsMsunrnEF2YwEPBPidzI5/nbHfyQMT9zlSTFM1cZ2h0DQniX
13kLzVlToPGD8UxnaLmLt9yFUclJoAVwKAJBbBCu6Ar8w28ltlg6q6xy9c7QgQr2PWjAgkBU66wl
jUgayXF0Q/WoKdPqLfMZHYe49eXSb339C+T3/JcunypOuYfJeqPgOkMdlN1i15w16W0gXtSdaP/b
lKBeVFK8yOlADkTSpT91s2zOXlqavRqzLp0uO54fQZQkpZn9cRU9EZpH2xGvlsGPDTgXKDcN2hL2
ocXqYxslPrTKhROgV3H/53/LKzjB9Q3dgmKpS7KZ/GpKKlfdagEzk8XsdJfJF/BqwyYpZ5iBa830
svnKgytx1XAEaAOvSIVGVGY0Ch8rybdU7hvshw6KE4HA6NzfbtgTfXsXi9Tup9av/V6poPJpruSV
J0i7znrThOiKzdQhsjBCmQWu5P880Ecq1bsTboOVuVx/tM2Mn2RlDEVL/yGiHVkA+rBPdYOCsN04
LZe4ee12AKfUC6qGIQD8fP0Un7tO1e3S6SPWWgmYcmJ0NenV71+Fenr6mP1YPwPGNNksXvuYm0eF
QK5X6FFGMTJezf3djO1gO+kHk2TlvaqAp3f6ENLDplH9KA7JgMv1jiX17btw52/67UGkgnbyGYON
OIQzr9zd1l8hHFPTFHK82oXnh/yhhJ6HpouXXqAOIAlzB3Ld42ctB7MqRj2Bk5YJ54znCBhrNaDV
BiiOPyKBh1gW/FhsNZoXrvP1+p4VdQjrvODqXABnsc5PTbAPyjajQtff/cmXAqNfe+1c60t4il3f
BDjsSBHtGiZ1jV/Z5++JpyNz4JxzkLP6LZdfXSbGCEOamDYsdrX4lYcc2CGV9S47UlDqgTl2xXGv
tZqVm0BaXnxUShhyFQJDKxj8h+8Od5G0JjYwX91iSlbEEf/6rWKEJrFrAlzvt4cY2w32ZL7t3rVp
cbbyKrWnoU8eRnyu/hPJ4Y7IXkf6F4HpWNv2rUK8jcUQXOLZOyl8iJpEyOcxkfCUZ5S1iBwvpZsv
jLLv9xVSSDwIoMSzJQVHJj24JSGnlVyMQNquOAR++4rCEz+3u8t37OyQ3Ge8PzeT2Akk6W0jP/re
lGVolYsCe68EIfuT1XNzhAUb8bl7OtMAcBMvVRveROM2Zn1J6NV2euB08Nmjefidgdp8Q0SgJ5w9
FQEFZ3Ipy7iG1mObk2MIjN5PRI17U9+x6CGr9BWeJN8v9ig0OU0UADmoaqLaU7+hqFOo6F6fPYVU
+qAOOxg/fuWlluUf94tlnYobyRl5qFYOyMjy7FcA+Pr5hglj/EnOhqBBiPbI4VexL1SrqgeICp/+
6Huvvdp1S0wYVEPhVsxhO80I3wsfegEQ8jFzz7GwTQ93Hd2FsC1ICMM1loH/qh/0z1WlTj3cYN5k
cB1Ho57VG6tG10/wg6lzv7dz8sRj8eNCmAVSCu8cXSRRy45xCtvBtGCm8+dyFt+tMzbpVsY5d9hf
6iHTG1TERZ2pBV0ofpeJqX79bN5XWfYZv7+vpDclPV6LEfwCrgG+3Cm64OlpQyodSt8mxjAxfk1o
rUd0xR7TfkUHHzgbJJ6EPrVnnfLkSGBfKuwBTPPHfPSIbNmhv4cMsSsbF1+g2D3kRVunX+5g3vYY
5HrvD+1dUMNvXCLUkRrf7Bb7UL38+3kGAQaqwzxBcWYsrA7+9al3MCzkGm2x2KK6AVZs/gTmWREh
4Hb7NZwQ/ogi0F7Ogau+WeR1Px4CqqaS5809U8oJR2D43h8DhI2F5xLynmO3dFsfLI+ufvKQGQu6
XASLF5SiFJd6MW9PxBYIAXph9KiRVwiVh4yOHGR9fxyR6BQYCT2hUuQA5nsjzcVPUdd9vWir/g7q
/j9rDNA15kQiOEhbZyHakgdQH2zegO1yfcbUO/PXB8fWOSfydeY1UpLgVw+n/9w5JW5Mg3dkxIk1
+J+ZTQ52JKdOikoRbvg0tmMP5ZKCbRwR1zyNZQuF9CNRQkp4AKjmWALKHDA+gKIkE9dvf1Qv3+o1
yz84cmo0nK/T20ZNl0elWYxGL882/jF/jVOzpk0+qhZdGTerAPsoToyq6RQuU5LQasbJtFXzRFFa
6ysheGm42czgltDJFqd7RPZ25nOB1DuJJRdL1v6NsUdL3UFjLV3yEb0cNo8PvAXxpLCdsofzGfMj
kkErA8FjxFL5U7cPmNQzfVjh9nHbMNAsZEOK5B/rJ4shOpf8JKItaQM3YnzbAYPTk2bgxpoGStDX
lTVaCLOb5rWf1yebOKiXvquE0KuzasUOyoOrqjM8CZUvchBGpSqXsRg3ei6vZzgb0RvpDshScAxj
aBs1ZfkebIA1ZyEkhs/GcIfl8BJaq2iEdP1hDBaqu4DKRRqgvs+5v9SbKoCKx/3i8+SP3IFuwVBX
V8U5xCZ1CYpULtZC2WfhVlGjBoHfZdvvlx3oWuEXohGWI6rzJQkmWv0AZf4qizf2tY7vR8XYgYsW
OGi3nCJ08ZcTJo107t8m+H4Y9HToToKTkL8UhvdWXcEkhZibXrYnOhkYJZYy3OOyJG51/2fDoJUB
mNlCHa1PZ3WnbZztbQGC8wQTAQz+J9dAC4nulxwjGmcrBV4dQSsfTxJdLvWWTx/ukqnw4IY1mEVM
jOt3iv1t5kT1ZoUhxFncHEw8Pn1GcD5L1aJSWckelvo7d4lh6ZxQ83EwBSMGc4/F/7y8klDNnB1i
PcOQ1TN1C8VvddZBUdAyXLvRLXF1kj6qPD+Votd6DkJFMdTikmM8KP5zeUkEe9uF+ygtHrgEqa8v
beqrpDyKrdz4fZZQQZgG/NSFfz3tMVPf5EusIg03WeQJ2mABPGdIQtnoUWCfESGxKGs7dtyYcK/A
kEA0h68/26BqjcsJJ0IrDfNuW+4ikvhTBmxjiG7mWrJNjd46rWdtNoZvqIj7EayTgy+Dy+r+gNqZ
oCLyDhBlLy27zscztt6hYhvhuU0nvmvYyCLlZney5aXJQy895HiV5SwLnk5kQ9pteCYsOvx3Mz7f
PaE6etwvAS0LKxJn84cjiYLG0LALB188OXKyR6K3/83/aQbYOzDctXClzMjEoLP5cu/WFrxYHbvr
A//Vrp7xWxRWBJ9x1l2xb57znwBsltTnNuX28L+5xFgHHbGLlJmF8n/OJb2jk+axuslBEGx5HDUf
TuMc6VUfEoZAPwjh3oglIDI/YwM9Fys3MiHniFAlXBqq8ZGzfIUQNd3L2tJNL4nyU/Xo+/hqrASu
dAuzc3YHXkmykWMF2cstJmBUQtC6Di9lqD4BpOCm8PYwnPpNIfyEmop2UNF7eldKQmmdAFS0ISAZ
WbvWHZ6uWx7cULdtMh+0lBBumcA0ifC6G0a5hl0ZxVIL62CGf5U6G9TeuEOpkK/LhoZ2OIz2VbX4
omZ7YuMy2cm6rixuyc/CspSCYQy+5kl77UVMwCntYYa6xyiShM7hxLxZdxtnn7qqYFLuYlMHsiZt
z4CjjkATsauCPL40b6C/LxZkjIF2snGIF4sDFmG6E2qWE6++Usc6QwELIKPk0K3y3k0zQL60viYi
xbRaM/tQSprEtOyYNKoLMElGHiKvlIHOisdmoFP6lpHEZ3VZ+kfooIK/LnjrT7kDGeDCYC3eBV7l
BOQyO8XfzgXfbT++WBtpdNxIPHhbKeWnqutoAba0Odzx56mVtsNjV70hqdM2oVN40/6QyZ/4Nygq
wIRXcKneMZUBNJxwLuvbCljEo8lz/RIsWKOJ3FkvkRj7cf+lJnvDibXq7YEPfa3tJeHGsi8bzSw8
63Ts7jyHIQa3FSX+Y/JKMC3aYdRN67fGXjbQCxK6MOFq/WYGqyJdnAzFKF/loIW1xX50hwxV0soy
CHgIb11ViC7wFzguA3WdxOvypOwNAj90k1qJuowS9e7/0NLuADIHXYLvshc8N1LV+MjHAifoWlrP
QRgVpywIcaTjyhZPnZXCg0epCe3OSgROe4kyZ5Pm13RE4dzGtnLh1Npe5sREWO9s2b49l1LndnRh
Yh1WwW86NoOB6FyIoRnTzWQsNv0ZUBR5Ux6y0pHXeSDyE8h3WNzpTWJ0oGIj+KFYaownQL+ongl8
JtKSsqYolS5OP2ea3xkYaBQyWQorG+UL7lnS/y6SrYsXUstxVHx6/z5tDekQ7FICzWiADLPPKwsR
phkbcKxuFx/Ey8kYJWzbHHfaP2a1JNGT15uqJBiZq5/Mpot9TvxsoPkvxhzXoYh6wqbGDN5Ypi5x
t/CcFxKfvPtZWf7Hjtz8LpRYeeJlJd7V3Wokbs275/JQUgIrFr5/iEHEU6lNX8zI3x8Kn5f62Hjq
Hs4tBpA/wclMAUVlpJOtVmBnlIsRI4nMdQkME4mXnLsPYEotnvHihCoMG/3dHFMvgLsg5J/jnj4u
l61k46I6GX4BCwVqbHl8hQBlttVKkuvHCkwyLytL5Fclz6ZipTr1CemVnN9Y7DjbCBcTcUfcG2nz
Tve7Nk3dFyPqFYEI5ncGj5jZs3pObVdtxF2e5geMvztda3vfq5IFtMkrnRBlk44+RV+EDc5GIAvi
CcIQbWqDHYxTZL1oOPsQ9PZGGVIfH2PCne/z0c6bmzKQAISenIhNSUNo7sTUp9uWsnurV4e8Ud6J
q9bvzDdUOAiKdW1a15Gwpmw8dYctXtm5ob1XCZA3D3R70dhdKR/63UavELM7EA5ATHhFaKYtswmr
WjQYRC2hXGH4IaWjfSkXg6qKfyB1haWeUQeMgRV7K9gLhmxpIZFzVJeTN5/0nlVJK9x+rbQ+cNNd
RYlTDyFzuaJvpY0dIslwE1K17kIxXy/D62ODtXtYqowPlcxjozLpnjjg5JK/B04RHtzRUSkqbgSa
5PKnCvCJFFvZPdt++5quBO7Z03x0wk7x3nmrKqEO1FZ7WNgtn78Wiy05wHZZWa6xN0VWsNlrpouw
+wW83bzo85FPpl/dEJrOZ0LFmofOc/9++Ppwke+J5x6oe6xm0t0pWRUP87CE8CnHd3yK3RgzaWd+
fsRf/kKoOYzMOXYcagHVti5Je4mPV8unJwYq684H7D7hwWWuX1ecrFQUF9QuswgdnS3Gdta/rB98
46hEVZkCyR3YbKE8qcwpePmx9ukTUP81DxXmAwFFbQB11dO1I5RVlWjP4aS/o95kaDzLhjA/OiYQ
Gv7WbojOsif0thh6UB4oWfUr4k7oE7oZSde8TQcepbaOewdxuH9VIQi3IQ501sDwEZ0VH+CfrN/B
Few+wFUYZWXvd86prMQZOpgowv6XybcaKcnvRDVWPBDwA4gfnbSvq3XvgpzENlcoJLIlRoB+GTDK
9MCovHo3U7XaU8wpZJgQbql1bhxLuGoLwr+9WQe9huG/LCKqmmosyJh9fRocXMzC7/j7GDnZjSVW
G7Dm2n5WtPpwY0CZMpmlzAWhtGV+ynRzdFiyBC85LKgAwuDYuvN2J+o9kt/0iy2M8Tev64ioOFU0
Hb11abS1EkQofm1KZWO+2/mWq+BRQl8JmENurQMui4IacQrVzekrbHmP0V2oFut7dpH54ymIl9T0
pDq1AK+LJT+tQb/z0C4uSQODf2g0j10sHnivIpUxbgXybobLhsXFz6rszxsvIzat6rvbcaq9h+wO
vMsUKmnaB8R2S6s6/ZXYF+9IYO6Weu0u8VyJtbyRxow9EOEurUET8K6mh/VojYPDa9TQN4zmDal6
XTJxp8apgJac8MSBWT1A80Rx0c/F2VD0exd7MRVsuKGEltPD4xtPjwQGBHBORrIZD51S8tLRN8K6
QyhwXPT82LtY/TLvss56JyhNzLenx6fXZUYyKXUrdMvCWUkpzz0eHz83Tt3/+2Iz3UBOfoNfbzOq
I3r/9YpRiTGKz0C/Owadr+OgDfoya4W9/Qu/v7EVc4E+xZZTbdFUymSIY2S+satDCe4ZWR3pvzrn
CueZAJhzM08fVI5j2Z0mSAIzOOwtkyCoh0Ko95aMpMFAtGQ/e7M7q7xVCnO15FPkq/H3vUz+Awzj
M1lt6Uxa+qiYF38odtmasB+GIFLba8WgkqEtZHS59lQLw5ksLPx5OMRC0mZvcDjIdlEi2i0vsIFZ
IMOXBeLI+uyaxNkUb4Avdek3kJXXjplmeG9Ot7wzQt7calu42J7Uq7v3jjXQw9SLMabNfYZKxKmH
FNxmU/Y/7EZeCtSeiT6+sKt3B1lmD2Fi7kVJG9gGJpsqUnisNGMSo7PM7gf0pmty++0qjjlJ/DI4
IZlxktVp6lF8yUFJCdQNrY5fpAM1/XkXd5UKcljC3izAra4tP5tF1IB51abAU+722KjhqoqeeSoR
FdUeuvRQkXIqLYRP5WX8umtef5P4jCWOuyT1sUI4Rlv+kiInpts8b6uKfooGWivx5V/z3obcF6bG
2XqhHgcEfxE9Jglsfz6eLSo1nOidgudyOkz9tCP/EvrpPTOwBGw+XlmBRVicyDKw8LxbWm6MeS+W
QpvF2+puMTlTikRyraxUfVWtX3S9pmNoHibCiIIAI09L0Tbc7uEaYCDtHvyhbpLfHrlwuhBsAXuV
UmwOp9ZS3/LyVouvVLAekb7KzE2K4sfBa/W+xnkkInhq9VulSGvQRpCAzKbQIxbwcC/Io2a+aVQq
znOY9bI7N9i7+AKTZzIQ1AFGo5tRMjQhZlJx7GR52eKWUOdMLxSH8ZgRDrqedJVZsnqQp8+sgPvl
asHEsw+W5/250ZhTQIdWR3zvewAlJZrSEhbb9O3nr6FKb9STGm0Du4thl477WSpbfUzYUlvnck0R
+US8Ze5Wugha5sbrR3zaalrc9v3qlbffh2P6XU8Q0XT3yvP3v+PFZhhDUY1xcteVHdQh+YGPT1mB
ShKgJDRyaQO9qa2usyFX1dPvjOTkwDc3hz2TDFaBxOZKhX1C+Y99eus8SuuVbUCKPyt7WA9ybc1r
JCPAqde+C898AqCyYx5zqkyegtbVqVSnKDodcjRyFxoPM8poK0FpAp0TW5pRMDPH1ootmlyFB7FM
xQXD5YDcSdX0ZjUy+vq5+wBYVQnZNm1pQmNLJ/EezHOHpAaVow4vyDxAZaYIG9mB64q45dtPxetv
NM2Jj5a2wVTNc/o8tW1SHANN1EzG0TRi5+CC0pFA3cuUbW1+lp5eV2iZKxanpFr90q6qRKPBgz98
nwptAWh4XJ5/Uyb19gx+Dx0//9cY99cGkytRgdogWtpmkm+yDokurktXjWZig7DwnXPneccBjfrS
gxEXSZRjFF/+B8L3XZDEpYUaMzl1QnzAWP7nBDqip1aMHCm2SZNPJzgi+Wqf4jymHsprJmGualz7
zM5pxSMiC/ra5nPSWGAQvp7Igi28iajYOBPN4+ZLRnCfeGH2SfYSAU8tCjc3joh/WRAViO88W+Kk
wZRNeYGc+HQ7bZYfgewPrd8VWZ70RnBOQewrYyLYzx7146lLOwFB4DyZpDP3FDr4iTfyITZkVHqX
w3K6OQumjN6ifgEW4FCyviEz0udXeO4H9XHKRT1e6V2UbNlVIUHrTJnONQSBw4cmBLg5sGTjoTH3
ZA02LNwLzuGlKBMphVXyV8lEywU803wX5NJLc4ra1dBZbBEXEY9YzShV6K5qLIhwnX22fwfZ35p6
xOhnsL8XqMCVAd+n9MplfyzFD2LXy8eQ4iV+Pi3Wjuv+qEGTX/BERxd7GSGpWrqwNdROSln/C4q2
eySAOIcXYQBTl/cuB+IDc176Ju01uIG68xomF4Uw+rniHh2W64msvISj/sbaCoEYXcCEMiJe/YUo
m1FJhHdxQyl3VLvtat6a1SKpl2fXpPksb7HtQNySkgqZOiU/k8o/KQSjFE8IVZg8R74ZDc579qmS
Z4bOFFyAlCIwY0eXlXEYG0hCQ73ISoRba+CW2RCWhA5A3sS3ia8MXrPIXVhd05Lguw7+IImhzbhJ
4nyyeo+v+QPQv46Sw6RaHkfX7/ToLaR/TrnMPp3C5y6o/jtx66gLWRXFXuxYGQvGJANARifl7rW0
NHOeMjkpRGIomJH0H2CCnykC2E9Xf/OrFHNztQQPkSjmTJPpQHdDnsTfi2wI5M5reHFdodQTfWpj
dfZ1PmIqHSQlIpMRSArNgyQGPCes4IosgxCCa7slucukq+PCWJ0wrch6aLwsbjDQY0Orcksb9xDE
btBIALGERP5lz7RfIK6S43Q6BCMoSFjFnzQZfUBOPOA49bPUuarxYa49S794XHoYuTNsG7VtdXOs
xcX5ifEnJGg9gaegl4dNBNGNxwDcDmL2cbyB8b4F8EArGHm2M2nxkZH9rMuM+tf1DrnsDoxhy337
mU0g03v8LKQfWp3/JhPkAedZVqfwPSPcQyaY0FfR2mjeBT8ZrmC9sZXspcnuZny1razSE9wBcJ3m
jCBUE/xMyiUW1cQtdEWS34MS8lpbnffylEja13aHYqbESUgpj3za9WOriwdZDgFtVR+RNt9IN4yw
UCG6w4adyvJ0Wyx7UJIl/eydo4DK7NPFIFGXDMYpZGFimo3L0JmilqGBNIsLYcdLtPEtMQiPL8Km
bTFYRoqDOKLQdzFbRUVIldGkXy5H8aez4u+ZTi75im2gIlEZCYUD/CW/oveiB+Dw44SFifTmytmj
PSXKGhMn7rsImmdIz3swv1jxfL8LjeW26j0JXzmQgyo/oXbgvI/GtKnDYVzQCv2J/K1cVeZzt6b/
7Y+um7mSgLUDS4wh7AYvpeZO9XGvhVnM1P/zcyaJocUvM2FXTUiqoOXJ5163c6KyVRfpfZ+OmWaF
W3sOsVXxVybUMmEOUwN5QhiUtsEuGDkp9yc57QdvCbTr5dzMkvR7C9cTuYWtzO6TVC9BjS+76WqL
MOs+QjFWFlt1xi+5xtEaPX8tJ2RVtdVkL09vZIMemSHo3Sc6UWgaecfPBIYu+b6ELswiVhDwuSh0
UHrfRAffj7ZXZhsUNc8XQb1l6huKqoE+yTzDP6uc4niusqjjf3BlHRBJr9HJi5bAOiFL8gF//Buc
meLw3NoEDJRQvWILeQKmXQJlPfo6Q703XocHT9MSUkc8MEPX7QUH5CagW2kyWvF8o93cfvwTTv4v
w6jjSMcsHUf6M3m4SQQE4hhNSUiu4BSv5dXzvKiwyYLm0menWHBm35pdoMU7FRvpuA2To9nN3U8h
iOtE28uJpytlJ+xJ86KGIluvkloB7117Ivl53H2gS+m8AILaZAdCyjYud47HMWk2ZScTr3GRmlmo
/x4ZCEA7GdndMItu6PWuMSsPvDKkw5RxzTwANFPfmytxH50CPN29XZr2NNJDHNwi4UM8jm0syI1N
tAqiVYw378+nktcM7UZjJzMzyTNpHspymhqu/5mNvVmz90slKUC7LugYnvxzAUE1yZllXATbCqks
TRI4fE3usoMyYtnOsg+7KgN2Qb3CH1KWXqBccMo7hPfXTwb2WLeato0aHzS7suANnnFAwFY19r0V
Eh6RKbgUTnFatn677BW5VHqmICUFWIJJQvVqImXgFcfKE/7DQorXJGJny/JlBpF9mIx2eP9R4Gfl
F6pE6z6fU343INraTqtzQC4T7h4Tjd6hK91tGsZ092OfOWiZJcthJSxaPfayuvDuA8CjE8y6bj86
KbUpEp/B1xpK+gcn3Uq+UbGuu1AL66GKTaLD/Zv7y29nVCtZZqXNRugeZDUyPI4JrdB/swQc4VYI
UwMSw3F+5rNgZALg2xCRj2+7OxRP2IohqkJXZxAiTop17a751BO7GWh5wbnlyAtgDOMKLCItiiei
QLWrQZ8/SlUhd0OEUFjvZTnEqRp/LKcw2mQ4sBefOow1U4fXhw7s9+aunkda+g7kxM3fiqG9jZwH
NnTy02v51w53N35pe4FMbxRQObgeV+psCdCC8gSpIyDfD4SgV5dZTfOAyt2jE1Z/C6HvCowEpzXb
PIb5sKmzpxr7sxpR5m3D9x94paQwOiVAVNQVmzefkDmdZ8O7aet9YwTEvMihm2hhVVWEPMgmEguH
EXkqpdXS9ro3C7/NwpY1wbt1udKSRdy+SF0T1qiT8upvk5Yvped8jSGndwnKu3iSEEE3ABlZ8MCX
/V0hBDaK/j4DxxlUJaNFi3lUgfmtc3PVXaJqX2BOXNDuWWaqqZr4/gGWYg4A/6Gzl8i7qONWktxa
TgRH6NBRK87ZGhkA+LjoIHt+T5x6cmwgb2/vDI/YGt91TbWTbw83mjkz6YEqQ/nIWn6wrSKqfdfe
Vgz3fEnK6KGTFDYk10KO37HgrV71hOZalTrbp9VgBuPeiTugxliQ3a1jF+QBDhGJXIdJ1CeAQaTn
yQcPGqc0f9PDFBDh8JhcOZcwyXTulgaTPzPlkiXrHPsgIy55lqyFQ1/ef5OyBxhyO0xqyEVMs2Jw
AYa77N0LfvUpmLwgnX4ZDPrZoVbPL4zayAH26dRvcBkwsf1NwGbIgCTc6lxwr9/ObUho9ikCnhHL
I15lFB5Z/qr6YynlPOVz6P77p22d8z62Wly7Kw5Owof5+KAA4B4zbpzyBX6HSgCUDap36GPfz4KM
Zn5uRtEt7aO5cFK8T3aBbuUya+aLPl3L1NLkpvEKImS2pNR9SCCebxZT5uS24Xi7O01o/7xqREYR
mqQWepHIpnCj0UqvTMKCJF6/t5RRE2w+ZSyE0nxj3XCNyDpBoSCker/IQamfYLfsSZ24LY/zHfA1
mxHbYnitolB+o0s71G+snEUYFxKBX0mIWqR6+MIO+vtCXF6c/WlF44SVZkOL/vVWpbJSncQJW81B
N3WKeWHqQDQzeCkrfG4WkPECrkX5pgICb8fr6deujiiE9M5/J0JEyo40GXcVfnizk59JZ9WdBf9O
j7E0uwsDYSLTIWm2AEuKbD+wGXBZZYaw2U9ef4jLWHqP4GTCTp2cx6e7KvqfF6/8aPYNhbuLWJ+S
qucu+QyNd0ylAEtGTaUJxAzjTckofqunu+h2fHqg3qtgJ0arjdu9NUyIbYfjZlVaJgPO0PBX6BKG
oEYai0EQ721tMfyokC2HAemtr0ft2mJgDzriYQvxROHxY0gFTBacz4oW5hQDGOktfOs/jN1WHa9/
UK+t+pIXky2RFV3NciChKTOkyXDTHjAKIfx0TcY2rTKW98PJ4jjc4I62fIonDUchTeJSJVTg/Ecr
QJGSEoZiPoV43vn/kE9sxidKCvIo+tSetSxPtcKJMBc/OWaXdy7GkdF3UHAgL0juY0iC27JcFAeC
woN4CBI9QjImgZlB6SUK53oggMIpX+FCnKuvZxD9vJTp/QnzTUcp4CQlpa0HKntSg3N6TgsBzVsJ
lH2HkSRPe+CbmoQcCAivRb6E99SR2B5Ajhvkx9C7eBOot+C8uaffG6/+NXq7rx3sTreuwNB4xsyh
swQDrmAAAjqQEGtt/3aFiSS4SNrQXqJ+IuEP+16w+5KVrG/MRbNMa7sfZUKCLbdTtre4m0CAKfne
c7tmiHAYCqfFdLoCEmeNI9RDhGA2UNbf9QanEFQS8POygQquzmbosXbzc6FeH7HtiCPRssvhm08H
HWfE7vN8pfHRNzS56dDETuEttgKMLS7zReMGMwU19blZkOKq0y5Uol/98W0owWJFGtDroCPYfJxK
MmhZL4VRvmHSuPy9cvL/P32j9qGwnqMAaHcP1FYUl2XMP7kUaxB8g0YQx6+TAZaBa8oTpTyX6Rkg
N8bK/3x4rY/pf7NlhTeSuF9c+4n2o/wW4WvfB3YCyM8sWJ96qCPzSET448xWzGEf2421UaB/x2IL
gEmgmu0kboSx6P5l9m6y7k7cn0Y9VR3KvN1nw7w77O6K0arVsLmcbVJUOYfmkhsXHppaKYYbUUC8
ql/zzEQlgCOy89pWSf7jdRgNttCEApROwa1/OvxiF4JOYdghkyS7oYOgOMPYK2LSkIRS7I8JvoBp
z0tNP6JdNXuJX6UHC0HWKISNSIeIXoFynqjYA4ZSnSraieGVBxXoJA7vCtq2rSt5gSwDsbaigZI6
V9B5gX+xXNncNX7Fuaw9p8C4dmZWDO7iCTgKJWvTV9p+b95+qLwhFx0qsmu5rhB+Vq+zEDPzYIUt
ue7PHiqtxRn64kmIPptAYyxCzdDrVntbAfue1ihEboPyo8rizalYmvc36CCRdf/YWWLmvDx86+J4
y9zGKC62jgbgfbz1+xCC5b/DffZzI/7zei0IdypTHCvB4CM0SNHlwibxuJJHA30SzBO3lLOP1PcL
gkgNqpKIrD2BBoji2D7O1qXVWtYxut5ZND7+CaLuwlpKa3TvPRzRIjRWeSFJo/Zr9q1kUPdAwA9e
zCxlMc0IL42C2V6fbwhrEW8ynpKq63qO3+ZpdsYeNDY8oZHrubEWJY6yMurcih8TXfiysTvA1pXg
n5eH8lTVtIMOn6iCpjJ6qGuZ7G9Y9dFNO+oBYS23pk/ApacnUC0VVf6AX27LwJy8vDNxjj1m1vth
7cmZcOXwfX5uBZPpi3wjHTmsn3FV9hwuL9jkPPezPVHeu3mQzS1J4EBvVVed74H51/4Pz6aoGKz3
YoQ75BuKXX34oer5ar/XPL5iwIe7TW/TZNZ8YJZ2k2ACFUFB3sryUYmq9z+S/GeWtblz6fwyum/Y
bzh86CY6/2t5cdlz6XeQA3/nfGGr2vTQY/3IiZ2FL31mRj8j7SJCrfHYDUlBg2CkH/wNmw/dzYOL
q6h8UibddCxZx64DPQMTy/HlOjxfFqPvYvEMejb+ndBv5g5ig7J2V48yDjbSekf+oFkuCcphYb/l
/+B7qc1cpHULB6KT/mlKoM2WyID95DjKG1KtjKK3Fwv6uAy2GKZdr4vcxjFxpMY/HN4FA2ItXybL
CRpgFFgpsFCOs6+kcpag72leG0AN3d4byH2hzXO4oD/nZ8CW2zZcU7q5AQQYQ7cBN5Z1Aa3xw+Bq
wQlP/p78mLhy+ZsyHEggn98Gp3v7Sz6XAbpABWlEREINlIcLvplnrGs04xZcslEtE9mG+xoKuAsr
52m9CD7cQIG5XaHRdTWfJ9EhV3y4vtb4BBpRJEDIltJ8Autdet5dJnkxA+c1exdr9CYW/XeTQuYd
ohYlKsvU3sDqgY4qgPOnDWZLQgwdaNu/U3GjK+H5QJtoFfKAVQtjeFZmW6QoYWsoZOFYsMCXdW7T
8hJvQG162FZR8Z86JD+Qi8C+O3mslFB++8BEG4nVb6L4L9qiOmH55Fm+TDGSCG6L4mBhwbn95eXV
VaUD9iyHNsHUg7qBIzYsytuMMH7BmnRA1VkOrggm5Z07Hcna+KWyDREVQBVVkJyRt29ZSJpxP28C
/KlOz2xpCwNyVnjIA/jAQ8g+iuAjLkDm8m4oMsox7nt1Z0Geh+XGc2qJB8zUbBE/KWhL24Pm1msy
BE++pHVigqxeehLSWTuaXAvjgFVLfCsDiVl9Ug82CBEa++RWH/ahm3SF4gZW/XpLSSiqpLIqF83S
p34ohFehIy9b/AXiBIQbPTAdrhbVExUh+wwi+PUSk8OtuaaqI+5QQknkGKhiK7wrxIoudQQoYpCo
HLsGHYuOq2yhYEaVtocZZUFqZD7+jewyFKQSvR0cOHqODTV9/qw+VGmJbYCgpzFazE2K9bpBgNS+
iL48jXryt/qqWYLLQs55SdFwGY8p06UoTRxOT+NQsQ3p3mSD4YQ25xO8lwKX0eRG5Ok+QYiQ/Ce0
Tbmu4P2rqE+yNHzDEil1pm9K94mdPT8HumiDF8ZefkC3N1XY5FW5FbO6s8BwcgvXFVzy1sXODmov
klQGG57Ybtwwmdn83SOGwS8+NGnaVnB4axLpRLFcxccl2GAep7qO1OicDtnEhev+gT8TlFT+UFD7
ogN8egBK3uw9LBkMS6xBxndT8nvzAglZkTEGuTUBgI0mQTZmj761Fvc3A7sgvW1VHsdQ6jKqDdvO
WYJOXICa9O1LUHL7Lc4+dLvsA7KWrfJZJ+NVN6QRIEMB8hbSyDYfZoCcu4p1LrteGMsDUegQucDU
aTkkpWuKf6q2JoxI7AEOR80bRrGy2bz8XeUdtF08LtoH+hHKXjdE9sQLcMNVT/FZyKt3cFpKo8RL
5XPqB0uOst5lSxKij1q4cr5iOc1jeLoNCAtOwJkV07XuP4vPvDYvGu+OByU3SgDwsdkA3h2tgF7y
JH++sejnDiMs5lBClqSvSnBMbPckcIwZR1Wby0tdwSKN/Ydi9r0KYlQmZjdl6r4wZGMkZuOG/V9l
I5lqQYQdOGxD8yoTmTRMEAeytT3f90rJTQSxnuHjtJ4aPDrTXC9IIxu9rFWBdO1MyUCHj359Q9pO
imawXfviNI0kCLleuxRqIwwGYPortSF0LjrzpHvMMRkNQXVad6q8PPp2lNetP1CHHDk9J0fP3tVq
clOklwQV035niVwGeRVJXmCnwXO8EQM6IB0Gc2DDQVS/vzMwEcThX4WjDmz1elGn579r4p8t7FvD
JiplniCok4/XBOHOEr6dx26hIQgJIAaqqQsUWtAh60EpJ/mQTqwQ0PVk5aztDNAZsRX559mWPC+8
hxLFOkWw4wNvBO3IFbJ6OV5jUBFU79Ey8HKOXMQDs/KE+6+Qv3AgL4/rHfZvoshl/5GIKM4loEs+
QdJLSWlVhEHAaICmxMEXMuG6UBjw9aenjLB6Rh0FNBQeJueq+4jg0VNLtF+FwV+CIA3mChpAptJ3
GO2XrjXZkDATUsxMpZm+EOKcM3PGrq1bYvZtQOF9Aiu+0jl8SKoIAJcsj35u6DtF3z9lahL60x8c
orD7F+coIXcFZOWz9GSxbGuqRoYyk03FkeOkwZAp1gpZf+CsbbrTYqL9oix6AyyN045BbuEWMv4A
aIvyfR82uucrSzTGpuQB8BYCqEY1Bf8tU9TBB8JZZJ4Jz6UFtNKYlkIZRsKWiBUiPDdlQPr0F7lf
kaRVIt/jjyypZt93x6jT6fxIANHmD5HQALHp1EZk2JaZhsU+Zcf+qs4vStBVrlMV6l+EsGqmrmBp
v5DoAiDOtmfXIXzrgcvUSJzdUNm9IF5sA+fTjYBFq7LrSMkqYxVWGc+K+YEWiR5f8ur+Z15IScft
nJjbBjN8/6YBTVEQ11oWTJUUhs+PF7O+2yaFmEtIiKqcYn7beSP28s7quLOg7Xds/CGj1CSUqidB
+dV2z4ylHrTQuV+ucrWL1J+dVJ1L5Sbz6BxGYUHwibW9NtJxIGWtg8mg0JxnSoFBKcR/LoHO+I6f
F1nOEWzGUr1gKw6Bb9NLvInJZd1xANFIGuqNQSdg1b1gpZ19aI5EWCFZUZdQb1GI1htxQf0sNo9y
uODHz2udcANKiOQO5J73xZ0rz8seqjJYkd0/Z2F9KaA9saAg2ltZtysV351S5Dc3WqY+m3NyFoVY
4DAorg1q+AP2s4JeJ8XjS/LXsnewExQO1e0JQlKrESqOOR3mOqwh/+f/PnrV5mmcCV+rz4Rnh3dF
iQTE2ljFf4pCs5seWBqTjk4Dl1c2H8LfxayDAh2k707CJJeZ8JX/3UEUaG2pSZofS8j5+jLYpNPZ
zVEmZWMNOVX2WuQIaT/+2uboFrbWzqgZsNOyoPfA9NMjRGFCeV5Fpo++l2SgnsMIVp+Q8pROLsWm
U8HR7+XRqrqCt2iGsCMZb+i8WHbbM6UZl2NdU1cUjgwI5186tTfCMqbqnq9LdPU9frfOfsNnJYSV
6GyTivSXy0YlQ5r+guF3Y3rbAzWbFqTpU8rZX5YSKfZ0ehar+9J96jCZn1RJkTWEnZqgViwOZKa6
5nIRczfqnlngxQK9KjC4Lrf8FUCHWRwJUofL2boAQRiJwGPXUry2LcDSdMC62hKUkYwMVD+X8brO
nTdeAt7mXRpM599GbAMBUN0PZqgWuSRyEicRI3kgkZiPD8xtJs25LADsftUfacZaZsLGA0tGBUow
Kn7nGyY6tm3W0pqlDQJjifUlXZM1NmYfF5L+pFSOjjezeAhCCTy5KU1hH/j6EnHJI/CEffUUe9NR
BiDy6OQXwtpF2t27rU+/iKTohHvoRgrmKcSsDPzOpWsiGZ+uHE5l+TByeKWJMH+OhWvaq45QvRJj
olZSO9Ac/dxbt6JkevAUVd+PD4BTL/PoS5v7a3bvl/LeDGLqteEUxRZ/Q1LzGdPhMlOoTPR5ome1
x5fjZ8VFKwI8W/tU7pUwI/wJ21qsCo0l6d4KVo8ASCZE++pQ1ccUeakuYB6k4UgtsjuUak/rxtFi
QJL/SxITI5HjcG+C8iLH9s5RMgUWB/IOhBUAbcK6A+VsZkDcg2n/sU8RSvQJ45JsoQs7howMelzS
WK8cKQQOa8YuEi2krepvpczk2oOSGth21spEz2SBw/JBEGcf/xEpn8vVdIXBaoH+55O49ZY7bzUm
Icw5LmQt/Tg8O/r9tiXQGQbJFX2c9fV7LFlbObnf4ccZRjjQDFzFuyUQEdQPANgzF5CqqzJdd8Ur
rPEfQq9INsTCePLBIR82Qe1Zc0n6aHsp/L32G7HjiKjYidRRr3KzRFHGmblbqP2BcGMI7iymUVf9
x9Yh+w8eCGPpyUl30PqhozdOJRhTcN7sO5uYz9Tao030bNjV4BWgj56Ta7IFiqU0Z8xwKlplq1Ca
h96mNh8FfsAs4Qs5ybxMb72/XtPmnhh9HepGRzmqH2hwlmJ78VtZUljTiw2SCrFh/nM4ljhG6FM1
Xxd5RDcJomXrUyK5ucnXIY5rJGutj+FyEGl8oN+a7cMsK8qUpZTXQ0ZZU/a4lHCk7++mFR4yXI3z
QmtKfz78++sXnbl4gvJoJukE9b5OHRHZswLGy042pq8JEISxEGn1rcFY5QKrA2g92uEP93/3Qjix
94se8cEtH6C8bF26/IvB12QPIMh0ff2G1QvzAoYx/UVcUQXSYHYj9GnMwfPi6F6UTaXA/eBSNKkF
EoZQPRupaMFZc+FDfWZ5An3TqGhhMPj77/Ma9acOkUKg/HnXsrvtANFdSLyw5U9D5m1yhU6IL6QA
3C0NC1nPG7QjTElmQEa05/Qv/VwcwI+L4Qsj++V9CaijIhPIA09R0zM6PadMq+eiZ9shiDYGu3Ru
bUb3oPlzAKwWETktx5BbICccaO2pBe8XghOJBNkDAdpq8NZrQSL7nakq5cydZPWm2lrQgiEe4HT2
L8FnQ2XVJLwBIYLP1YlmTaUqJqJT0QLVPHNjM9sC8VtzZ4l9l+yfd8EyvLoSXwBu+DCUjuuYrtgW
0Je2+aaH5bhedNaMQ13HpKVkudESwMbGAdmEGnU62+iwPMA1tU761IS3LP9nDLjWrHkEtISgTwCo
PfGJHmLRceA4E3VO9SGKdCFp2HEtVRQBM+twZF/GoRTFeuzMoh95IADHrFZBV5c1xhIgt+h8ycwo
5swL4GUAeUvdnVLOkxbyMf7ImoS+/e/d8BHR5UjXRP09rpSPABNcPaphTvGSBt0vzNqZ0kFCqj45
tezi+9TCu+Rh+G4KNcVvr2SY2DOO8fUhA+FITWMh5ufzbCHXc6Cc/tXQvD/aGCQDED6UUon+ABG3
EWuz7AHXnKoYJA/e1s5Poy5Iiomq5n0v4/NQ2s9OK9qUBn937VZ7cv+AKmjT5sNv6nC4l1PQF2t5
sbs5AwQKT4RvnNjzyw8Nv1GThtWLt+tRjTdv3UdTBQpizUj/uMH0ayP8AmycHqnHpPz6DlHdBNom
KJSUsj7lhSC24xM8mKkE7rrguBmTMznWF9cF3autsi74DNPUA8oPrb+IpQVATpYiLphQrrjTyHcy
Li9rKRyfhvOfsaASy3Hjxm9m0INibzbF3msFbi0I9qM7+DKBwLy61BgFGhdZFdc/weAOn7aRR19S
Q6aXyfem+uonyiAkF5fEbHMB1/dIotEVjlox0ihdDXDCClGzPbALR/YU6dBmtAi573PAPYtXimBb
rnbrO3M/m9ERpxgSnzVCLf5n8UQuQtXO5ZkXHzqLeODp+3VuPUDlhWnXrvJ970VdJT0wqcw8aEd5
+a1V9B42jNFUr6ZknyKN0Dc0DMoCNaJMTM81rH+CaPZ4gdtODgGNg0Swj9PbdjU35udiEQZR5AEE
u6OtDXsQ9BKYAKFR6EiKy4yFfSXA0HeyUJNlL9MyklhZMZU1n3oLjEFWVePrQBAYq30E5iIPH4V+
ooDp1AcYmReOri/+hjys2fLtOug6IYgRiNhCN9c7q4fCPoYzIGTkdZpgW9d6ycCU5C9IH1ci1MXS
NPF++EM1u6kqAhlAmJlTZdrIyZwcJ0Xk3v+Mu2DxwG0/+DD6x/b1i8O4a2eYSedVf8CHdbWxO3Qw
6Lz43xwld94KI0o8m0og/Sk5b52ffJrq72uysPx8ZnKHqt1ebvpVYSN+uAK9WRz8Qdftt485YDBu
i5bxbiZzzdMHJpn5TO2KsolasErtZNSqqzLI030HIW+ytIzaHyteJXASJbia7d5AqbcXRhaxfHYL
zGMXoKHWYhDClU5L0XCJs5NlorZIUft2D5GnK8q41n8FRvkx1YXhICcZVwdxvZuIQmMjShgps5qJ
ppSxP13KKwpFmB1UXdTzHmiW1jGuIIeezS9R+JLGAqZqxCUMQgj5FXUWRNuqC/i7Dzrugu4rT1x4
sbUW87loGg5OgpmrOARrmbcDptfF6NJP+eU4rBgzZ1M4r+B1Gwxvozyhf5HTCHeXHENs7pAeA4vk
X50ZvUAJmvS2/2VXD9vBjSv11VSd8Qv7wXpHOftiqKTbqqH27xlzK5NmTFhARZstuUbI3W53ym7L
D7aWM/byLFlUQhNZ0JEiclhwHjLxAwNkp7PK05VmsinVSqgfev490UPnjfGOI+ES+xSI8n6/bvd2
mzxNv56AKXDTiiJunv2bixpoRica1uE0u3SrW+gJja3lk1fS19YEp45csOUJkuRkEWiD4JCBCfpA
HoYUCRIyZz5edY/1k3Yv/FAVNbl+UkEbn9aScikGbXwRb1yehDAWyyAeSKrQ+HAF34jB4sXV+kHW
5QeMw9KMTDtNMLGYHd6krRTzYwWFjjFmZbcr4ZI22Tt4NB2djIWW/KBc74a+xKzlihG4DMD33NbX
6E7P9SjSBtcbUi/j6uijBBhBWvWBA7JmcNDfjlhBguJoLkp2ru24Db3XUXILw/RFhceTQkfJTehV
aQJUPfalAbjgYtXRl5q5YsAkga73hj2Ffh643oX+g0owE30mNXpI8kfErvnD9VP7RFr4HijfzHFh
fypUT4Xs/l9Ks507xghDabxB7aEYPxV4HIqSQ6fRX7Lql/FOe4FkO6RD5wdOxl/vIN3qhlSLowOR
dXmD0OzRGDyGDkXzQayU4P1wN2VZtKXQJ3FkkuNs2I1G5C1Nw4aqVL1t36SeY2VTgB+voLUZdw89
bWf3NDBh//zVixt7wj3tkajjbuQ8fpzqnr23vSO9JtiK8u2nDkmnTE/eF8a62sfWMLlAlIv+sR/b
ZxAeF7VssFQu3H65Wap3AAj+iUawT9aMP9JgXtPKlmpUYFo949t/JM/Py2nQlADSWyoPF6MiNLG5
Khb3MtIXLMVIRvuvoAOnB3YK3KA0ksbF4ijGOnNIhzjIbguqGlkTRmSpThQgySqcWWkNeeljOUlM
+C3KS0531Ucuh06N38UGzMlMVP6Q8gxRQDKOYsFSymbn7w3FHRgwkLARWhuOxRQIZXxw696EuD5v
kuf+8CJHmmlFINYYxyq2D4wXbMwCvBuIteJY20K5FS6pnV++jCq2KjiKIBTBLDvEdLbklZlwe7yG
ooDQo8wigaBN6wMriKOSpSu/lfaUg2wCJ/HNP1Y6QPTAa8AkLp8Eb7viI+QYCkx4untq68xWI4Ik
b/GwFMPZeEqOcLOlsVmnjC9ucFn+GYKx5LPgR4f8hNae7vxO8u6mkLi/Qc1+osfJ4Mqhq3uUzGkE
hU5O+a1uwfyl56VqSBTMRsoAE3Mr0t3wuFzIC8pPKM1igrXao8SEiTknds+66sHtz97RsETA+QLs
hWvKU6jBfYkQoDk3bNFl4SMRNFU1VGJtmQB17o6XFrDsUGZuQKIT/v/uIrPHSuZMOQdtzeIToW+o
591gpe3LLp+U9j90FRnaUf92wFsgbM08VuYuI41xDDycWiyRTszd09/xwkwi3KeTJ3rkADTBd6/v
BFANVHmBkO+gCNv0wXdnAyWTqRA7ddI0VEey4fM//6XmL/B7JokhTQe2asBog8e+Co1jGmRv2l1j
xF1QCuvn7xYmU0Ndle0zH0P/FCp6Ae1f/y/GfJU28fKNZHfPAkb6Tk26ln7G3AgUGO3TcYFYLL5a
rl4qxunY2z/j1vc9IrJ9BP5gyywBsdZkyh3+VitHglh/DjvSy/bZvuAh8CqbXXdc49RdxTKtXS0L
0TGbLpAbD3YBEA68DSKdeOB8AJgVvivhcBkbItgFOpxuG/d3KNV/XfCSZoh/ds7dY1p7imJ2Tyfp
D8xdTlyu+YvS3rqXzAE5TZV9RngtprVO+CMfrKUCznVj0m7puRpqaHI0YwdzzvklQy7wMeLyy1gZ
35ktHj3Vn4aTky61RnkP/gHHzQ/losr8XIC8yBX0yQCuJAHWOcZWeilJjud8bjZY1eeQmd152psC
74UzloDb0nsS5i8i2vnt7r3Yci5GaYOoHPaq9By5FdzwrnICYhFRdav1IS5h+t+nTy9TXhnH9ErR
Vgy/lGom/Qw+c2I2naP++q+jWzEStt+AXjGiwQbEzxmfgTmwfmQV5gUkgbID+CG6pEHVS/hjj72U
j2vkAEQcrmLs12l2NEUyHqg1OR2E9YAP783slpieZeJbQ1BizEDnWeeZW/ESjm3y7MgA/8n/lObS
bNh89tx+IKGKfaCtVuOsDosIv22pPzwft2hx+V1oAblEZ8KpqriqebtZ5KTGbn/Ed1x+HJQNt2IR
4CuXSzjMKGOx72MNuKUvcBjhLovMjlRYNBtZDVh+aLumXTDaq9pWtml/5anbst85SWGfMk/G0Jd4
gubvyoOpNB/cjRhNQ6yaXqonAkqsBbaT+JqvkKVxYZ1tO+P73+xXeHiXNgX8ivwz08bHH6iAxpOi
NhJQdKAMLKu1dfviz0JJuJFB2vWQA7NislI+TA13pU4C0A2gMtsG9x4Sr99S2tV7YhFbzG67YYiV
18tD0KyWzvoLI2jGARvCxCKPHweDCTX41GnwREkAk5HMxMXWueAk+l92m+bacOhnncw2jyV4Izeu
1cnMxL0EZ2unPj8cVHCZJ/Rm9yTQV5GnbBstDZhYnA+g02QKqvV44UHiKr7EwVvq/Fk9fXoe1o7+
5Gc7VJjbXI0q1R0fT9Wc1Uk9KRVkcitzYKN7DzP3tvy9fXDXKX1Q7sVp8AV2b5ZHjtzJfU/Po0Sa
ji1INZvfQTsKZP4rboAsMM0xx9tcKUZOH96IsH30m9m8ee/YeMBCKLcY6jqjPtqLhhmlg1EJMVbo
Rv46FmNADtT5ho0Z5znTbPVuFMS2aheZxTeejZ/iUsskkl0StxBpm8lT9+FO6X61jTCFLZdO70uC
6wS1vKVLHt4v1LYvwHDZ4ZXvlCzH5IvmMYT6lIG8qoo/mDPCk4med4iaA0jcwuC6Juktydg0UP80
MGoxuuHps62R/38r9+OXBeGJME7FsyUVjxKMz/SASxFGWFXutioljANvy1pHll3OPS74M7pqf2zH
c7Ix1zkyR+0aTvIyikShgIYbMJxL5mdOuD1+imBV8ZAYluWtTXWNS4jl/1Vl32jrA8f1EpAMEOV4
rBHQYNajowkUDw8OA2a066bcdrfF4Kror2+r04toaNGDwWzHnAcov5oCXWtfePJ9Tkd22k14MS1b
f4/wJXgnga7CBK4rAaswj6fcd1vTHuDFJtsOWDkDXtIULzR72obKp6x8OG8k1EE7SaNWVa8M/d+a
ZtCUowdaO++oE/yn44xer3rAnTiyl58kHpx1gGhI/QHYCIMTyGS6JmJDyjhF2NNiFfwmonmXkV53
ds3Rn6HRZk70vOPLvEES2F30PTd5MjMSt+Y4Ujn+CFv0IDj1HvAXTDROcOCdVzKtBIhax0H5YJ8/
3+sPNLee18kjMdSnXrgEiROQPUiPUQzx+QCf+eGE0HZcff6I3AiYirNzgMvzLMjNe3Ycb5eMFbpB
rNr1vL/J85J98QqIlbU08P/W4EIJUQSDJOGSAmBR616ru79ka378p26xRx73XCZkGjMJ9kQjEF+T
UQkCnmD6+B56gOmWKiodF919Vv90RH9xYccs/RK/zG1aNYop7XkQ39eVr4uu0p1/e3sFlDViacT1
fDG3TBTadm+tGcdpUt5+6mLYwcUtfuFdq0PSVVTVqtXOVOWtUuVLsYTe8ysK+GNh5AVy1+pxSIFh
r6CzSyyJ+bQkxToWHU05Mc6uFUqATHyOs89nUaQGmDKC5XYMVlZDgVe/G3RaJ6ksusXdsd9ah2hc
stm7CsmPXptqgvLDhaeYVMuNdgmR/6VPLcWDzuGVgbsfzxdWomUMvUS37Fzp/DoryhjMyk6JnRaW
bjJHJ2bnClq6+Zfo+xvt/ulOFmG7wMuJkW4dwpCQEtO+O9rtcSxce42B/X+iwt1kIdeOLq0w6BET
laPv1IBCAzVKNlqYGjmhCVFfT6LyG2pqqSlRLOySQvC5k/emn0DdQrVI0CB0ENwf26QDoaabjXhv
rTjklf84u5R/oBvpSDJpzUwk2VVAONHs83BrtYn78ryeoFmthh6SB0Mb4Z4hvy62pRAxsl6GsxYI
uPdmAk/UgV/sKqId5dYBbIAsgMBN1bO8QxgXChM8IFjHJyqA0/vk0fxZEvtFWDAY9eKYHY+4YHxi
XJDfviJieDJmfex70D4WvCCdf8cRCfUIrUgBZhB24znpnIu8PCUlhD9Lm+E0uA4GzrOQGQJ5wcZf
Uq2kJxv3rcES6FYtgRBAFMT3vzG4m4pLXVhOCTxI6UCcbxZ8GAVayPCrQ3UZHud1U16JvzwOvfmq
/nXA2iNTiIt9NKYBM8BRxqBq8rRa40vbzXwqXe5Ib3CUp41B8t0fk5x6HkNERLYsf+YckuggqNbk
6MGNtX3Sggpk2JijjVjwW/WqtXcLSpoLGWSGnfIufm+dC4H9tJDP3fDDLdNW00d2DTcjW7cMy8Vw
xmjg3o1CgSQ+OvIwOW2IC+P7vXidZCkk1h+9wvUa6TmSDhsawTKQy6XwMkkxuqAQIu1L0P/yjGDW
lYZjtgujs/AKTM7lCTqW7VjKB6XU/WbL94uj7CCB1U14I7Scd7tqfqHEr8jN+oYFygDlQC/OfJfP
Rj6ybtSVEMXdVXpT9uQc04wIsHJYbk4waVL5Wb2mCKAFUGn2Se6PSJ2/ZlBFs9k94OgWl0Q6OXEE
1/zvBQSJdYahKN1Z1zLHgcGC8YSpD85DbCRtDIyc6w1d5aSa0AAo+VK0/N6knmlyeo+Uh0pW8cbM
0o7RAGvYQaiznr9VbfOq1Hiet2MRFeQ63aTsXB4kssrDrgyR6ZZ+d/mlaoDO7XRoO9OCB3+Dbrwb
PfE3R7n1VXuCiiWbgSg3ERI997gbUqg5aQsj7rMdt4su4ZakScN7PkYn2cv1+LdxsSsEGO8Jsy6D
tdU7K86WBhEXURLR9ZrogAu7veHuQG6mVTSIvHkoHRPDRUF8cSx2u+dv63621oRHreGb6ZtdWU6P
uCggJjDm/obYBMft0YN4CJOnnScDT6IDYaAbSSkQSJjuOloquRe1MskDTpjka6WzkXOoffyIqRpo
Uq+Hs3emW5iCqWtM3SzRNhcIip8qlGbXZ8pm6lTeOXWKegFIFYa/yzPxHme2vbLYHc/6PdYMuc06
3rB92jDjVNhiQ6E1XDx9wYFjMlf93JJsIpbpK3+alWhS2Hz4OZzwxeoOx1/uk8HzF1Vxd1eLqERw
d6C4/mmxYeWXiI2WuP4Oow6CTw/Nhc8m7vpmr1hA6U+ED9F+ABAX1FByPwbmcLrCUBQqvsViHcyp
O0sXyDHG+a/7izdZd0niMhZumzz20MldiKiUNvvwQ63esrDp/r0zfS0J0DhNwh71s/d5Hgo5KgcT
fsoveu3b6o2URHEdv4v4x+0faFMH8uXB8ZA50S4drOjnKwhHpVmqJgqZl9Gcla69eKFteKlUbhiW
1xOnDh0jedchDrxafeNT/+WnWYM7SxM8I40hGFFmUgTjM+a5LKGaOneplSlyZnutrGHgGF5HbC77
TEvznEBUzorWGNx8JeO0Ij83skO12Jhwfu7GR2tGBFVC4uMWMocIqLNYd9JyUelAz8hwKVs3pyv+
fB5X+8RT0L/UJfFIWNfzsQgZodx2O3S2SBOfV21rO249+ksLw2/g+pHCohyFGH1V/rF+Cd8v8a4y
ruZ+FxzE8/B7xVnIwv46ryCqHtfhO4urgeXKkJWV369p10X1AJivc/PQ+q7p5o1fEGzfGs3xmXmW
amRcYeXlAfbaomPK+n2St9N3l0iOHl5R7MBlkRH0AXOj9/Bv4sjhz/L0jS2VWq1Wz/6I4c4ygpwv
g24+AFbgtel+od0Us2x8yHCzN31vzIKlIIm6ngl5G5XNn5HPcMKIEqYUJARB4ZIJLo8eKWravkMo
vdn4YCSEL1p8H05csqe2uGKPd9RbaDio1eGv9E5slAmLshC2qOHdaCr7kW1tj8SoKynw2P23LCxI
Ow5VOR6XqZj7k+Wgd+Y9exiT2EmipUtVZv0Tstot20zN9ok4UK5/bazf4JirEqgiO3S+A5JVwNJo
LPOE5FHnK3u0GmhrXwdFowHgEAg8tBz5cZGlIEWoEgXzBXBL3V7n2CDbCIhKMnm1sd+OFxQqSkh9
37QiCStY4htDyPrbx7ZlOxO69FxZuGosUrrGQn7aTpRGpQ1+WSQM0Rpse9DbEJdEur1yycQrZaNK
zdCJVg9yZzXRMqvrMvzkKiRknG2miPDWjgdCrfNfGX75UC3f3DnBSF+NUnCWi+4rAXKne+eMy2T4
8htYyQUE4S1if30h0iG9ReGJV6K0lC+sgZMz+CEXnI444JFnhMEe769Wusjr5z5jrBIFooxJ5syX
Za3kZxq7T5YyNkQsO0YPReQe6NU00I29hAemFa2U5hdiuaY3tJnGR2B7EfZ2xX6VgqiAKJSh+Zgr
YvH/fDOSkMLX8xctrTDPdU7i7cRQmDsOZDeEf1liDe5gJS+jY1uEMJKCKzPQuLLM6qkvXPKYQGuN
Ir28Oj6KF3ah+LM/V0AM6QOW4LhwnMMyq6JxbvIPOkC1q267DNBEc0/Kmnp8wwTHhxPQk2W0pnPE
pYgVH0LV/YJR5bsG4zSRN9T9BAyGycGiRzGA/oOQ5NbzcuuAEeiVjeAr5rHlyaAktODdR+i/B59O
Y3UDe5RX66UghEJEyiY/yXvZXuiaGEKNkH4pmmAqyA54D60s5XDAM4T3NVUxjl0o7Y+dGcfHxdCC
xvTMfnnc8Fh9fczfEJHJmtyKIFJEk592YHPXn2yaLEFCjkeXW85IQoGr1iV2RyH815T4DfEsF9h8
h1S3IbEBeDbMDlWTRoEJ+LGzzRvX+E5Ui4qVt50PW1+q7uG/D+ibvATVSZlo3hDLxSNT0V4DeJHu
wTbpUdjUulR+MDdxdm61wOjlv+Fc+4VNIm7j/zaqSFoa45KZ6oe1nQNWFAITfgQL98PdGKeKQmGT
L4q7GWpMckPNEAhKNeaUAfPy/EjZKT51GZL1tchFiyTZvQzaHjTkVDBrNS5vewUaUTriVuCrhU7u
8COQ+3z07yMT7M/w/0LioB7OMbrjOtWwgSGKf+3j0stcm2/XsdWLIGXRE9F2JTC6YDhpLWPDpY3L
1OsgoSz52NKmLgdGyo89WMyhQ5iCZCeF4mzMaLNBh35IyFg7IIGNOa5y9FO2wPMqLm6dkakas6rC
Y/3u09xYucLmM6bDOyQN22q+Aqbgpb2DntbxZHrCqbS53mR30CWqI3L64jT06WUllEVtG0CKnVbg
OHFk6+7pgk8elcsDJe7OhD0dGA3R2cT34D9MtqwZx0xRrpu4bSYvpXYMELffmPY16IHVujwzqzje
dwjdvwu7YltdpOJZE6cxRoU2zb8Q3a0DF1eI4onsDc45nzK5+S/4erIsE3aF2Hk4RHpYbniY+6hd
rhYZzwvIUDss6p3CTzqJu8lwqetOe1eHruu+655JtNodee9HBxwZn+DKqptyaFki5tK0nD0yjifQ
S6PWRqCtFwjWlrvNz+tLgc9JmzY0g3EpD/3oO+YmTujBppLKPuePABn6GlUrTn37oG5etu8/3m+2
R3DCf6lWCwT2qb+0FkzWrxzu6+7ohGSlsUf4VBeXLcA1dhdP2hjPhg7Np7yDFq947LDTip4Xue5f
oAqIl771vcpQYbwSMY92Z+DYv+EsMnZLhGys1Z3b1HiuUIfn+Thmqu7BerlGzUcJFgj52WBE1UWJ
ZGAFlMgtKWBFw3DbqFgjrn/6etWlbp4mPzr4ezuJg/OyZlqxBa57UIyujGPOgvL1iaboE69qiaNf
XiUgrpAQzCwmAiF8Vs24VsxbmR+stGhivGfdjdiFXZ10QyUmST7e9gkZjnbtOfoz4hzpAr2ZRKFx
yqhYUwSvynC29YO74ndwL+sRAaG2vLSok9bYs6ZHjRJg/RG0VUW5qRMeQc32rA6ryS8fmMhAugzP
td0XE8D7J42F9J3HwpKSVf36TTlaADC34BKfr/Um16lwx/4D069+04n/UGijWijkOe69eNg3KvBe
eRZtqkFcZNt1gMcCZM1SaezsJygRmERdMjosAXtZwZjl5wPqmomV3KuueHW9/MKEB90VEJuQY0dt
/CTyoifP/hp7YsJHgl1ROcC3lXjP9UQQRHW+7pTxkxOjchJULUtYqhKgQTzQCm3l1g+iDjWxDcX0
6pmcwVHNy5CJqpU/YKwrWRj1MDpKy4SB3o+bQzQ8euw6CwCjAfgQ5h+0L+ZfbM9amLpqHRTJBUDF
zBHQoEOl89QQ2OEvMifjK8Ybc0TX9tQ7woKlcl0yjFf/2+2GYDCX52ZCQaZzfLiLdffX87r7HvWn
sL8E5nAJmPxz4oAWHvGDEHCtk5y3wqaayZAKkWd1sWq35roMfBxshnV08kh4GfF5E2X0hrHKS13M
san+Bt9ZpeW6O0AOFwpwYHwLq3zZyf046jtnuQ3HeA65HXm/butFJ7v4OOWsCPUn+tM7+ClfdbY4
uzcMCzxq1pdFeaUnRIfC0uNRSW8Nb1Cq/iBQZ7PvvC2sUdJP4/RK/t8mNpGOO5aSYLjxNzJO55S3
heCupMDxpsA7sXhsbr3l8wXP7ImM+ujo5AvGtZ3uyQWbGJ5ovNtDG6fD5/6i0ajzSkMPItv6EiIn
dAft1/JbZcVzToUgd1mdZcazhkhVnCt4g94GzifMO1XV5WtyDShEBLaoxrwr7Bz1XStclTDwNGtg
EDi072Pp1ACW8S6Cd/HsnC7urSjRZi8iVLf8AeWlMBQfmS6qNic/S52dNHwmeQwUjzIs9iPmxFZd
8cJPdpECnXqHNvRBkXZI3tNeCedKqQQHv3SLFDo7KluiGlKMsSARPCnFNstIs8LFj0ewAlnfN/xf
1Xx5cQz4qmjYSe80Sz7o2+0mB6kvFofML7IMVtjDAIgAgl654cjiMpM0pITYKA3r+jhT9KJSJx93
PD+mP7SujeTrkfnZ7VTbzBoReVSD0LaUhnB+ITGUEL+hgjnNAiPJGtzNijsmrEfTeOoZexVa3rQ3
ER0nQK9jFYGR1ViilvfD009xEmLzk08hQ8Mfxtw/uXoZ/PYsWGdMJc4EURxFcnU9jw3rWgHRDRls
es9NbN/S8YwCRYSqPauIOgkpV5jqse99Kry+32nZCT9Risc/9+rW08aebwgPpHjfKJVw9WSIx5BD
69tkwiMveWFq53bYtNqRE56LpxpEBGxqiPltALBt54Sx1MmcvCYlOULbz7J/NyITiukhO59nAw3Q
tnKfmKUTBo1MbcZgyfoQCThHz6m9n9OICNXL6UBrN+uaQifWcjQ71Fgek6Mv/BGvFU/AnA4rzxq/
jBgeFfPHGzlnYhRKQcznuXtmqmycVume+0W+mXW1LZXbTj+tfahj4yOo/pC1sgNyk0R98Fs6Ay7b
Qb3ope3xSRdVSDMgcjiuv6MFWnWDUvXIVU5R3OzOWkwMPVzfG7ETlYRXBo5HpsfyPNTwJYVihNdu
t/RRUBKBa3xn9e7m8A6+EogvxzxEUfje+sJeCGoUb9k/+ZrxuLGWyx/SwKvdOC3MTa6yHJ0sR9UD
/WnppLslTZP2LpK6OIY45Chsn060cWkOVbWYRIyyPZWi8PzHjagNuGFJ8XqUPIiKNYgo1TjoxgxI
CHYpu96wFRz23nKeF+9Xngn2KVuUFmgsZv+Y8Y7F8GSkfDXuoeDsOkrnXKl/ez63W1xDasNP69aA
3PfqnHeBaIggDg9FohDR9PJ5VzK4skw5hg6d+Ux0zTbasmc8Gi5M5mBHgGuPH0iGGTWA8L89rnTo
3VK0wLB5fQKImVAQWuyv1QkdvTXmJddNtOg5BEQ/l3fxZgbiuE+3lGz6tB5nU71npV7pP8bjKVsP
rjy4S9eADKmxnOXS2RHxsi4OMxV8zKkhKdXPsfY8IUuz7dNJChYS78v/xgGYjbFZCCc4h5RWJyGk
lZ+nCkm/M1rhSntp2rMlZIrfBF3x0RPsvMGqMRZT85LdzL2c1KB/x8XTRRRtq7yZA0KOOZ8q3+mu
6v2djUWg2LLLgCmtf9IehFDGS27D+fkH12HkW3xoHeeMAV6vroYQnCtXFKwX3RM7+rlhH71mCO8D
4zqlFNSxq3aCeNkZXBDQ783NR599T0LoDaVu79YFnVAny0uN7Y77RGtB48AGwlR2ug3UolUnNa60
TixvRFN0o5phu2K4TkuegqfWU1vmo79lWKFCTjt06gfSbF2TRqh9X90hKGZLXUaO77yy0Lk/Klaj
U9N6a1dFEM7Whjk9btDOIUsEq1dZ6AVjBrojN7zHJa7vhudUWbCQenYrVGZm+UIBo++rnvXhyFKz
c04u7dx1zmR2AcEFhLrDc1+gKJvenGqMv2PM98FZzBFlOya2BdTYpFm3JAPCMfJhKIHl5zftyCBK
ZbemPUrnrq8iFGgu7xtFZwfBE0Xm0+xsfmuzr4ygIAv43qpxtVHbHaVfoJT/l2rgaaZFnPSorAjg
LAecghEq3GNaFfgt38/CjJ8Hxo6dMOmhHeND8DA+88PWO68MLsw7Vr7zZkmdag+x2Y5lJjVZQUi/
btoxLdMRRr/IQr9A/5Hf8tIJJvmggwfBhNBYp5T0z3BtmgWkRxIOpoTSBU+yfyLIB9qzrKZdzVcO
TE5e/UXTU+wjbJdOmaEBsC5tK+LvW3qowMDa8CNZex9SeKw6TSxmXPdOICEwQ+ZcSZCAWlk54ZV6
J4k4+t3weWti9QbLOH46qW74DdxeOGPyc+xk0kdq6AgE+LYcnOGWpalKQl6XR7p1Tgf7+bc/lk8a
+NcMQuQiq/tGeLQTk2IebOX7LaQFblEdAjTG8VVhipX5sFXB1+HESYNPb3bRwxjiKiZ1a8SFCANp
1McJzsBdyDrgb8QsSsJ/uRJXZh1roN1Tg9sEIcV5IRUXHQR6UjskiJCF92Nfxv2VZnoSNbp/a3dv
PlsqCLUQ0dJuoDKOkr0o+75UCakUwihmMkSShkY+j34pOLKpomL5wnOCwh81yZ17ynk8Ifddxm/0
Epw+JYTi596NEDTrp+wJu4eIfFGnJpvPpW+k3OeoTyy+KhJMsF7ghHUOmLn2AmhrmWwmrbEhReok
WTkomSczKlJu4AKswNXtKy5azV+2FGCLQCxOR1dNUyc018w/Z3l4Qzr+t99EgZVIkv0QEPHqLBgT
xc91DpjXY9WloFpCpUyrGwjjsszRuPC6yRGwnqqfoAhIDod9lmNCWQ4CHTdiHeflB1ul9VUg9fCz
zsJX0EXZtdF7VMg9nDwvbdu9crzBs8ajvODpIZK74Qqt4skWHwz/T0ZbEoHo3UZOkRrOFlAE8th5
y38XIIv4W7g7h8x7MPOALhhdxFSHtDAO6txTYHxYHPLUFAwiqTC3WcEiIWvUgLEFKH4PMJg/PobU
m7NMttRt4y8FnygQZyaCloB5DGlgkPn/XmV/uwmHBkEWhCuRi5GLaOWq0qsu5sKBOp96G5QfzifC
vJTSLfQuEAfzNAAt3Frmtu0ZrO9Lyz6Y5+ujvd+/qK4qPIOpmKrEWgv1FRfwkAC8e0+FjLasUOm3
WS6UaNWnG9HhFoI9vqG3NQuva/YSgASlhZGIststTnPynJt2MrGZkFYaZ93GkRu+tCwGaPcV5T2H
WL6d6N4cN8PXRC+DsoNiwpNF7ea4XmmkuxSCYuTy1muG66zMbXTX00Chv0kWZKJZLZL/1D8C+UsZ
sjBv/uzjNBserNPXcOgaPxk96dz0w6QDUQ6uULQE/OxcMcc1vEK9i7Dx/nFZPkNc7TyaSxTts6An
6GVSt7m5O6zrF4dmm/h4/LyEu2gNetUMcyrclndChkbr0Cr6LKrYsF66BRMPg5xeSsbHO4QpiYFf
gywp1p6WKqQBatB68W/OEj112NbTCvTMRC+JpTBauC4CoNaPJOLtZj9SsLo7wYnaelHLiS8M7sL0
Tgui+0A70GTKgE3oRrKl26OGcLaRNykYmLNVAWVJYEECU36g9l/mGjWLTrYgbCDZ3NNlwIzYWFDU
5M5N5qp2pqaDq4eM6niUNqBPYTiKnPgAWEhOZKMJk4geY090vZzGaug85+TuN+oZTcBEaDV0Yo+f
G7r/nb/6YMCsX7uaodEQbXa4B62305RoJ4ta0MnXeBVFJBhCim6ka7Zc56QoOM+e4ZPxutsu3sDO
N7rtrdmKz+OElP3VYhA+OVNtq3zUku5Uuy6KdtXlDRIcXNAjm19F1VVfaR+R6A7Mr3oZu7lMob0s
4QgphsWhOEOVSIceySA0BLV3UaBqOXCpZSGW2lRlW8SLl2SbruQeWJNuK4oyqhn2z127vQfWRETO
botJnAD633rrPchNkPDEOfLRpWbZk5AqxjvFb9yyapnlWqpOttx0Jn8JbE2+R+AzVufnv5sI4q3y
4+oBlFZyckajgCmM5ijskYIp3z1BCu0+UaG5QgDKlKssHYoPGVPhqYNmu260htoZBUwbk12GgSM4
pKPW2bZ10nVQvCsmvUgx8zNvaNwUnWUBeGah48JkbS5EXskTGSG6z5/tnbk9e6HIIwf3/uGcosOp
Hr2AFNYMEBIrytwoTG/041AJmUbkNAHgBckKZRWYzMz7y3ZGLKDsXC1t5cIzO8U5/0Yxyg1FlCc+
n/0p/Zs6AnH7+tzZZVLEMkcslhHNy9mHPQCBxNa+azKNY10Us0emtAbRnvsqvMWlkVnkhU2bsr+c
1YnsbvV/uQROS9Dw6dF+KUqberbjmkJPpVJD4wS5D+iaX3+7v6pzqN7O1SMEY1eO5fn6BPscsHpK
5L/qxxRwUVitiqLbTotRCT+u9iksQdLkoAzSwXh23n1JAc+BUZCI2GFHhB+gh2p0CrbNYjagO8Kf
OJhIgRevKRBZpQJybrRCL29Lcv5qpDoNkadw65pJvUDaJPlzcZyK5K2CMda83f1TJTi2RvG76WvP
ryCB3bBw2eUjOE3rGZXOdTGfoXYJNRKSxjPMBSX5VIgQFpBEbpQhjTpuTkHtHLOQaFRDPzgVcul6
Fcjuls+hbOIYFO5QgSRxMMDA70oETRPFWH8XThxqUS4M8L32tDtdn88AIVOHg3fDoR6hBtAcfP/4
339LCV1LiGjw9BUBXrjtkayq25rom5wFObPptacg2N8bMjqYACwDW9B1pfdoeagFcMb6x2rp4q+q
bHc5iC8G1wNVy193pe5YnqgJpkU0mE4J+g82kiopL/qHOCJbTqyPIdASPJaO6FQkt/FFPHA03NM7
n19kRZV8B8FIRqLuIO1Gl/23KMtKC+dyQm3j3bXt0wkl/G4qBDbOHST29+eewta9VannOP9yW8g3
e+ZEhn0gjW4oRWUHVwoAen1M41ABpyB1i9jGFYIlIGdzQMP906iudJLZyjRIs6FpQDjyVNeErfdN
CR/YCMG6zsmOq0m4+RC61zFbTFclHLWUS4DncBTl+d/RkesDr3BlfoytNzkuoaeHq2vj3ZkOgTPo
0TTAHhUrJjVMfOiY844JRSY5N84uNJPVK+yPjC76292Qhs4E5gWF77cDGEdoQeK6sDPc4C+4DySx
CqLYi4iQbYHGw1JTmFoThZ75QPQsE5b/z1t/6hzSA72Q1OxzaSj8YNct7IUz4qXOyIylGPtYCvJY
0YtMwC+rdnJlAwtXkioOmICzJO/dA5NT7Any7R5ESigI6UkiFhxkkfC7CkGCwP0dL/AIR4gRptk4
BkqgOIIBRWuj+hQPvIdrA0B8MFnHNPG28hApBoLSNDdIeXi9bnLQxFKuMmHn2ILCaFwGbxtB0Sty
fFKoe8CIz02h+TBu61hDSnuyLsJ0tadDNc5YQ4n53viKzfNn+eXTKQKTHboIZKTOyOj21wSL9ccH
JsRm1myaQn6rJKinWKkmJ7w2zgZeep/ROIIavdQHIaRRf3K7WO24wQc7gWNXfBMQJMdZyG9nFukS
7lxsp+qsv5gE5S53YVsd0OOfCDIwmoo24VCoZQS4MyehF6/DcuIoihbeERfcisDVAvHK0vjTAgcY
IN1eMmEaTjDxV5wnOgezF+S+xro+/cHW2v3yshzYahu3M0PZumN9p6/p7zK6OCdDyFfQnIHtAHms
1wHzFl7JD/bcHvHpVOCLA3pf61lKChUfgWaMt9nPSR+kyNE7QkAQTyExZLNO9tOXNeMbEUOrwbOg
dzKXjE+f8ERgmFAP6AN1fTMJ1dOfqoWCved/dtQS6sXcFi5ADvO91D0JcxpFSBPA3Klc/0euUvMV
rxCHdpdIYrnmWHP8oaK8CQUVtMJXtjES9Wl8IZ8SGlJXHs/94YFI6ZGQQeslB8aapBmP8uIFvPnR
rv4dwTic/nXPAyQ+WBMgqnI3aok9AK+L9g2qYZJBRf2BIIwo6P3t2CnRmxQopqYt06/xZwf00EDE
fYtP4ZBmQ+cHtxLY+2EDTPiKiBwcldqKSZDkOD9NdsA+RW0tRiwGp3iGOornkg7voqRWmtkw3wxc
0AMgF7ZMS3xWPWNMzYs2WjgOTZBgWs63DxIs9X68IhvMH60FRtS1+o08LiYa38KZgP5BvaYBX0KC
bi0rsjzUHCZrX4D1Nur6S3sQST6S4qiuE9RUqVbKlfP35A0pt4Jpuu82ZyddIngJaHbEeQbFCR+o
OsINBTbExoXitGDNNu8i+7MUDqaer9v+1Iz1yZX3Uow1sNMZhzgsfA+ahu6TKWT+oKWXWp9HWAmt
HBsQpOOjBTnM2NqVIUzkSK27FlxI6ujVGXJ6tbFTuKxeW98eRPSxdrmrBXYaep3KO+TmDX2t3HLi
uGJ2XwqCJiGt5CoZ0WWpBE0/SpGDn8etlrIk59TCe6RMgPfhkyDjCYZLNTiO8G60NFyHPyPH74Lo
ZNXu1cBtcFU7DvfpyxEOFgJwhccr5eroQoDPljCQZDpeFTrKHZWvvgIcz2LhNt6tfh27VJH5cURn
VMXEYXO8nNiUJ08YEkyXC+14hsri+Q7pvCrJZXCVBBi5oZICR+WOIUADvylbT4VmwUNqY8J/1XB2
ExWPN+9UnOgI0QhA4NYkPDzNwgavZ+7NkRRiNpntNqnXrEowKRbNyx1YqxvA9aCUyumxBtOjhoM8
lt424YJQ7LJlf/qGtCcEllZJvRPo4FpZxJEeTzYtqpu1GIqn97sAF2mC/p+OdBpFLHr66Lx0HMmV
Xs4VPISlJVW7SyrbjKDQO/uJLTzcqwxVMTgsmRFboS2yjM5EWTLK7uDIs/3VBIUfhClg/xNe32R4
fbWUq2qF9ov6KAibsNiO00FXGtu8QrF3vH2dzdpQfkjsXceapDDnz2Kw5wtFHU1APH4K/wnW4Fmh
VEJImR3xxoHxhMSLLENMHpoi65M03PYVeBLhsPujyaizF6sofKFC4Co3hl20OoUc6UKcwA3WTLQf
kNNXjQlUW4Bpccg3pv/RVv3pZTSKg+9QsbsesYOjbRHb+PjZquRIgQTQY+aQ5qfwEDQmmhzMU6gT
oQUqhiuCkf1WQ21j09NmG5ynu62DhYgNBZPt6FZdT16fC9/rP+yyQgpoRaCSc7prXB56O+zfMIgB
zJGynlJcrMxdVTWtbqwDFdeGuJlxOvR1YIe9qr3jxCFTht0P/tjvJZ1H6d4zqE62Mqj9m+KKohNz
JxF9b939HmoAcfHFjlSr19LC8yxe/6ocGJOzCrjcWwkUkzEXEb9ev8OkhBCcDnGFWxmjSPgj3Nzb
SLZYAJCF3wAQ0QvzHjn9mR/81Ab7pJls0Pzrt2WIGaaf38VwVFCceGDXYgRLPYaPoAlafTc8/urH
OYgvubT2/qq4G2L/j+9cqbHqplKNKsTaGTA1uv05pY9Tm+NeyDQyQ5ETwctMdyPl6E7lFshKOhQp
ZtR9YGZx1rggYPO1SN5HRq0pIJBpon2TF4FsvLJhp9ME8eeY6SPTGbIlNrYMuBFVOV+p+jDXrn2b
T29lNaLLC98YNfh163/ttZQMOtXly++pqxdJmLkPrI6JomkBgndLFmpbDXazO5L0rIGiA8RZljCg
4mFr2czDdjSXC2aYXbVGDQ5FvXKamwsdxEdNNCwkdTnc8BT9ovTgynQPJ4SaGIeNyWnPW6AJswOo
saCUMNEEJvaOCOpg6btNxZxZaUz3sfoHKRpY5IsCMJTToAg2Cv7thzzRNSu3WffY28Cqt9O2vHEZ
melEboB1ZB0uY22TPAIEt3RzC40iaReSIWaU5Vh8OycVaFpoGU//ulBYGTQyvljdwVLrkmuINqm5
UJN6ZQ0GXeFFS3Vadwm5G09ZSl3lS+r1kfPtAC8+dK3haPLpwiG+mAlEBZgJYYcqb4FJJiBmWfQ6
8hH1ODO8RSwF4L/Do+cdO7NTMmF6gKIo0BqR6Lia04eL0CjES+dUd4hxI98fP6AwMZH/9eJaa3BX
oymSG3VD1IxA7Pt3XU5hYfKcrFF1Sgtizo7vhY6k0niK3kzsO9aGtoC9eumy/UiQ1Tbuv27WzYBr
CbHNCphUJECYrS0xVG/G4MTQwKxJK0bKMzqyu9zEbRNmi1vezoVZ/dFr8eZ0JTpFaJlORWN0fCw7
VuVLe9JMol+nA5VKBvfvQt4rXPuHhsULVsZ3/8DFaswm3dkwScStyD5gig9Zol/4N9ooKk/tlBQJ
8ZYrs2AvcIf8Hx3t8zIxQNG5PC/CdvZhkB6MkGq1fEPVdYzYhtFhLgCJSaP5iIOc6SJD5wMNU/oi
XjKASfHAHUHtB/11YvTFIrxBazz+GrBhDrKiat4B1XAAfIwj2r3ieepPYQ5yrZy3qeOjUokx7aux
0D9Jprp7ZzYbd00slECPOfkuxC+ooCL7c6d+7XyCzrITSmaiVuOn0Pec1fbpmvEIkznZNcu+PhA0
HQRPb3VwDAPUTGlMS3cqJg8lT+V/oJlRL3E5XWuv/zK2OiD+ctbwQWaGulANisWIbdngCnsCyUDJ
OyXp4NzZQNlIwrfO5fYMjuOXrCJni4m1Q0zIOSYV2uXJRrGyTGOM5LVEm8FfudlLH0ZqgXMopnA7
HbTlyUOOuoKwE0ZPxd5OcENY9+yrWghA1QBfls/ly3E2PRq75LZC/RcEklDVik9Uu6EB+7uMxcgq
GW07xt35AQg1tQdntWuU3HoM6IA4FoKr1K2fl3BNfLBf7abdaQt8m/ZcgIZkB+nTr4ZhWdKfe1mS
GbjWeWK0c6Y/7l2pyggX7otLuoE0DhGNIvwgcOuAnFXIiAgix+tp0bS7cnstjTySrcgNz/+lPjDK
MxYHQnuymQ+NVIQVzqhgnabUqXtsuTFW4Le8z2LERq9JK81EEaamcQO/skOkv9nMAA92FQMbr+3G
mH8powoXhBlM5rASY6zw9Ry3btzjCdOTYhstWvFDVP80+fyH0rhIVS6jQ1HfpXQVo0Gfe5A6/U42
oHuDvwI3H+rKFW9OIl0jk2D/bJAuix6IbzUHOvfCkBwWJnrnJx6+8921DVF/KgL/i85f4wMxf8x9
Q0gajr3jv0vnMZ4Sr4OXCTtb1cL5d06MgJL/Tfl//PyvDzSGni76nZveRnUfunVlgasncCETwcUB
xTtzuE/HMevp01wsAHwJTTJGbAhWmMis0qn0ll54z2IfdwsD5hGMJC/tnpW/uNfowFiYgyJ7efIV
rrH7ZHa38KoXLUziaonwg3WCRelCCEE5kOyWQQ8237Z//saWWDHmKfrahBJuJEhpundZ0unvH6Qm
m/XSaeaD03GRWUkv9D/7vjUshcEidK1W8wo6ZYEKqsr0hxR2IFwpRVISd9oCiEHQX/9JYtTvL55s
FgnhGgevmUgJ3tVbzWZEmOCltM6kgqsdwYqz3689wdDAM/yBSMElVaU+VU8F8JVNvAJdQIne0Cki
G8hAnqcZXbCZRXj2cu1CDM8tjWRJIGQX4+DlOCvyKrSFGNT2+BEjnd6+Sbw/bTDnN7geUM75+2Eg
pccL7JagZz2yZxbXib+OL83e2xp7KYWSIx8RKjw3X3QoUarLJSEVGWCLB76Zn+tg4XS30gMOhIfi
KIY8VTIiv70HEx3M/vjBJb978Q+r4d+nHh4sLpU/uwUdYSQi25lNc/Kvms127cThuz5mpjrwO3gx
Ww7szt+Ups12fNjTTSNg1IZ7O7WDM0ULy4J8St67dFujfLQ1OuVQxi+7j77+duZTrk9kFpIGMpZW
1HRkDGBdUHg57OF7G+7mdWrzvWgQtTvAtCAaq2LZJQXJvUNA7mG3+MqnIrUPttirqrhOfpxoJQA4
gIl2B95E6Ntjuq+e2Xpo37VaoUcuoCGF0P6oNQCUvZtFbt8LgqdPIXhoMQ5yx4WBMDQ78vD1CKlZ
UDsihMJKF/shzvkSFNu6gzuWUO8r2ZIhT//gOZ1MX9giVTQh7lbyTknqoUNE/qipjAV8H4lbsGNK
3XJNJ2gApr7I6pZDhGDDezhTs7MvAuDmDk1DWmNrDvVFwGOAaCJiCoqSjpo93O9X7/A9yz7sQ+Lo
qiz4Us8feEk7ivuBBSUY4aM8VFT3Rgq6rNyv9voVwMhFVo6PxGVyowVvdSHNxaSqHM22/1n4Qhv6
8meIqbzvKaL5EeGYclnHZORVw8ol2Us7i4ts/wKpiO6e+kUZsyl0ra2Q0AyqeivozTjjoJAyOnS0
a6IPDEO5hZIEz6CPlRSDRzduUeKclApApvFVgLyWYp9Y6ipQnqa7d9hMvPomkXvuP9lTpvtX+Nzh
gzMvXqyeRZvd/ubVUUeWQuT2NszE5iSz8xDRvwooiG6AnY0kd2B2vJt8kG3Ipp4nzEHg2MQNl4rn
hHuI0QgCX2yP4erVtmCVLVHTU3WJzewggltmyH8+Yfk1fwlzBxIt6EFrBQxCx6MUdmY2Ov4rKYMQ
B6/a3r+N9D9hQOJNN8RRzVa8xMUj+khPUzrUACPn77OVP1ePpbF8c6lQllznHu5D22NmHhzNPHL0
93fOrmjd0CTc8OJ5h8U7qnXo3B4leG7aCUA+b5Ik3w4E1d8Ut30J4KeYhWxTkIgnkxL04MZuxHgp
Q4E018Er1CM7boQo6RLP2dEJ1LsSpk5ZlMaAN0UMMU8pIwFd2352wD6gogulYBqZMbArnCqFvKOi
AmW63I2b9veU4pEnJ1RNgXIouPHO4oqNs9Xk+dSbDANem/IORvLxLwxxfIbApZMbK2fhO4AG+q+4
JEY1QHai39s8I8doXkhs/Kxbn98vLj9dS6UAbzt5w2V9i67AwtCT+tQtQd7el8LSA6E0Z/RZMTUo
pGWttBdob792goh0dKItqPcK8Bw3EtIZ5PQHbMIG9f/aWGwbEfAm2Z/Gn99VnoEDSprra68YDXD4
U3IXXZ89BT52GIwlaQKybhi+nrY6zQvep/XGbnArHcAumvnnsUUxkY0i4JucQbDhHyZmjEXwkCx+
YOwdjlouFiIGMznXXaOnynwrCdrHrhvcVek7R5ZH6LsMjT1Cc/mLNXzYCs6noS5aJaKC/3hrZWQU
O9j9MuRNLSN06NUnwsHX00cv1RxoGRRfmLP3PUY+vHP5OyJHXKRutwdzU8LWmIBkoeyYnvpIX6UA
XBaQ9GvmNIWkQxvPhu+YLs+wL0XDyNBdU5kzQ/7MGVspSvqqVIkG/CKEj84Sk2VbLS8tStMv6cBw
MAH9sVwp3GB3qCnna4eaxapqm+VvoKRfVz9ViSFDB+KdzVLwI8lxuYALmhlapIFNUTmqV1jArvYb
CTC/K5JpzdhUydgQIHTigpgUf0erG46MyHP7o4U2w43Y83XHLY0+eFeyaPZbieodAnWJEqA7Fh9t
rET470NO52Gnpibki43K2PjbCjfZjqV6xmnBo3Z4MIMBmCXkxvZHfQxQU0GRJCg5f9aoegm1M/f8
wUImL72OAzZkimUNMI5ahvqxIgsSqKOXmbDwMXIAZpEra9ZaMC5FhVuKLSw7ifPCsnEgY7gGFig6
hcKM78y4vGOe914sbDsNEuqyuPSx84V3Imz0dY2ub932mEg3juiHLoUfnrP1mHq+K8NBZFg7bsQF
MEtFkNeuDWO/EAGSzn6/bkbvZ0HLSC48kyNVVqyka3QqkvdjCUoHnBtz36bx+NdqHy2NqXbPIAKz
xol9KwwdeqxLmhJXYnOhFVSCZ2rHsrMIkKTkEgBtR9nnZawBnlNEV8uRKUtw3TJlhzkeP0UJy4nX
2HFwsd8W6i3i/ZwHtPSz37aeZu9VeM88Ym/PXofgcjg6OThPA7DFyJWfEOT7m1gl/+iVhU1DMOOR
VC1MZoJ2qbn1yTOjQ4edWobxcwZ/ey5mwiAy9JaN+Zrudkzd8pQKHSO/M0POP56UMmK4GqIW5Tno
zKilEiOrWrS7m7/tVqYGeP+h+/sxkNVD/b9IDbtIP1D9/6vil+I8c3sahsS1UcQqHmZWotoEBv2s
VDjtTRdTktONePKtM3Tl1yTjHIa54XGmw8B5t1p7cMaDoV33oZF3iM+aa/niIuy7T7sFi87HOyvc
DVl+QANqN/Bhn9KsTkibhYsUFAY44a0BHCqNwG6ndep6jZZaY3IAIeXo3hC9+KSvmL0ixHyp4KCG
n4vssmpgyesiiAzOg/+W2QfMYR3cMqI/oUEPnDnyKSDSMjHzxPTpbgdJwl1qrKmWj+vAYOJK6PsV
mfrvJnHNagMOyjbZBUSuZwRJ17SS22F+aBQFT9FtkNHnYU31y6sOVFSRd/dpb8xdPKXaz1+9Mkdc
aaNDylYSyUkeISfZABh8p1NxUUl3hq1u6Qzaqk1qmiWyLWJj92dzWudTo60kW2MBhOrgmvHOoffn
CBT0Xhb/Mj9QiPPdi+mB3xJ2IKlFu5K+GksIz3Z7DuB3yYYH567+52a+C/baJeofCxC5cmMr2JDR
BaUe6vZsSksxxIUqE2J6LtRpVscV6+Kwz1any7rf1w8FrJ8mbREZ6/XP/s0cPLyMYujVYEg9IOA7
21iVEPS0rE7uBSArsrNr4Zjcz4nmwI0faoarZQ3lWnVt9sPBPJHG+eeL7LvJ1DU8T9QA3CBwX7pa
FpCX9ZuZrzPTUNkIrQqujNCIfK/IG8IozQLE5KRCZ4sCfx2q/sGr5i/imYQZ+lt2VH+RPeCsZFMi
L23DR61YiC9EIDR+eNSeosasgXu45ZxP4JvFkzZtSLibJVSNke0/UXVZ1DP8+n6w5rklGSHKuc1r
lnfvJUN2J4NcsoanWwlp9dEtXionzu4Pt9I6R0TO72HjiT4cisVp9SwYOjHm75ufou7YxSrZbpW8
M5fBEuvbElIuGZ/UBDHn59f29TDiQhwUme6bglHAjGvBXDSzaSVZd6hsR+6F2dkMRMxHbuxExPuH
UiEYfS/PajWCr7hDrBCHg2cyrVU3DPOnzy6O+gGgMJ6xHimFyadCXFhGcig/5yxkO9yU53li2x87
aRh11wuak/bzR3CUeowDf2e+OW8kfYjAzYrm1cfB7N+weQhpZG8ck5J6EI5tuu9qdDVcdYTyCKSa
Zg4sLIQc3oYwJUlnil3ULPg30WFH3SgK4u9ydwDsKDHQ5aCPQa/PXa0DGxgWHG2AeKjhqhhW5cVL
2Tg9v+LOWdpEqRX88IohjC0tPBNQzntW9m+mDh3VshdAULTXpw37WHAJP95fipQouImMQoDcKunt
bNYlF0iOA6MmqismnIufK+CBTWcE7Q+OtnyZV7vZ+2F1J39XkGaajcGoc+g2WF66yNagtmXwMb6v
/2AqtKFlYnjOceFnlEKbxW9TXrM7a7dczvvjdGDQDCzofGY8RfZV2K2SCOkaqqlUfU2TwCOp15fb
s3B0Fp9bQUUPDIN7nDK1DfK5HNQPGOp7v4+e86rJgf9bmz33sZW2oO2fV/kGQgihwzzxwr1NnTK1
x6yCeZs8PoTzGINGzJWo8WpBgIyVx5dCSSRjLt/z31P5LQh0idYdzG/sqgNn6DcTbVVw+oXkQsEO
8wQezzy92tIjryRoLk4YgYKVWlggjZDg9bPnlqEpaA7M0FcmCer9JM02Tlc+apXAnGv6jiIJbdNb
Axi48DV9Qp+Vn7j9xpW6C1j1cwXSDWRaVQZUjxfR6ZspO25XgXke2O4HQaFJQKCCNFCGA0uN0ktn
krM9l6sEhzPYgMG7f457UAXFT976rvIUSG0jBq9MSLPPNHM1ht2swk9v75pnubCERW4ExhuEbXiD
cNmUKYnAt4OnHkGOiiqbME87BQkZXtF4zDDN2uPjmivg/g0xkU2hy0KEFZDbwQ0572Wr7ztjbeSQ
4fFOx/MpgvWB7gLQUqE4YlP0CunSa36ZeSuU5x8AX+mBExJyXEKw4AVsof6W77R4imrbJW7LmDiz
7m78TFfsVQ0/YrjOO1Dff1hGlcfc8gAdQ+/ji6Lw6okIpRBrZoaYI5lTQCoexjT4Gwqef0qcKWy7
yPjhGG3ONW3gdynq17OiEPs0UJKKJnGm1wI37S7NeKvPSw4FSfGQJmijMO2QbUWPzbD6MlOPjv5Z
S/cU+ObI9P8J/xJ2vMeKzP+iEb598iy/mPsFC5oOClYNsAIWFmkPMFbEa4gho/ECKWyc5Nmoj5Jo
oTXBk5hLu3Pl5hWPdxPgDksbUMdenUyuipoqzmtHg4mBpHfXNkPvv+gOqjFZvKuEHqT9PRZqkyf3
I5S0yBpF87PNT9LOpiNg1Q6vOAjJDWA0VMmvnrRTP0xm/+kj2iL2jUrIFZmqoCp6epK7EQ8eYnxO
CiA7KMqFJ3TStLlIjfZi7hshDoS1pmWG0fcOftM9lfuKsqe4PAgg7HQkPvE0yIJmd4ySPLGcZA7t
VmPzhUWtxeQLi0Vjg3X/wXaBWTSCAFnbSzH9EzT1idCpyULxjU4cTjad0uqCKo8RQ2wiRrJWAL3q
wi/uJ6XpGvcihab9xo5oWQ+HPXbVo00Hd5hVaQjCS9GDR+1OqRwR89NX/cjYDBZCXOe+dXtwNOY7
77EFP8dWTufwYjuQ1nuw8utgNEIQ0DJk6ATQy/V2yRkXMlZK7z1Qww0F8nxO0M1BR9qL6M84A/6Q
JOPpDhAd6eIJcjEoaRyEcAj6MpsA+HinqBR9gIMIvkqh79IJknAp9X2u9WAEJ8ktZXN+QRzc7qje
RVpn21wqiiA2dVfwbnqtdJpnDG+48lEpGU5V93YgBi963e9sUEXFteGP6XDzX+2UZySbtgxXjlK1
M1vENoDJecdeP8TnJPoYzXNwOIVAoUfLcGEjYSc3GVsxmmpolKdgWdR4TGe8X7gljJUcpW9Ka2iO
MnQvxbR0ESqqZYeqrMCBYuYBL3OM22T2e/UiL5E0fyobO/JuGwNBStCvINKXKhQqgoC1M+2JJMJ6
QKPcyQY/8i3vUsYM/49UMhocZYTrKAMM2BxZO7g2NiYXoSEI7YPIlEDbmGupsQzHVXddLTtMZDE7
sofMJZ4O/G6X/Qas80nSR0CDyCKuADV76psclp1YBT4w+DAv1jDXBhKzeBrf+bnDQp6/XI7iA9lP
3AyyXa9XGVOv8wgfYQRxESaFypmB+KMeOzaaZq7TtvfdJxip/91//mXDC4FutOGVoo+iJlU+HgO4
FInmv6hlEyMr+D8uTF91lwWEtmiBVlGSBlySdgl5DDXSAzhFsBXtwXbIxn6/9LQhLFHHPc5D6rB2
45VTv59Lq7WG/Gz2Am+W1/xmXMmFf9NY0EXoeiHHpAS+tRnmEBB5e3+GJSw8g5uNrvBHb8h2esXn
uIo79pieodwb8XTytgUGIYa1C90zd9s4W1gHWzyt2wpKTRLm28hpU5L8/eto/8nvs0YMItn5WjSf
faR9mmCMucev6V93q1LPI3kDWmfNMWG0Vbu8Xmuv/w/z6vvBlDH8hd2l3kvxtbGU9t2ivpAJmEQ8
fO+Z29Lk2ouQijrnLF3BFl9kR8vRb68LQlvma/7dS31VnfT9pkAZyWEYGNfS4BDLbLUKGSt1q3N/
0K9FvfxH3spG8BENyPCF9yFyXcDw0Xm+yxtKBdyEOSINROh2Edwn3t+H7wc6cNtVC5jEsErsewdZ
l0NyJwKUrpm0iUy+KfJAmCBYtCAlVCCtGFybSHQSok+lKadzPuxM2Cexc12Gj+pvxzJIhMR5FzYp
NiQze61dXmpTN15qMqAQMuPN6VoYr3iqmRFdP9fj/LHcDUeGCgoVwuDFUbZlh1ofviqM9s0tcVQd
6bbvao8zkSIcIcTjmQc2PVvPDlPZWCCeP9Wnnx9pGqosVMIjBlfyzsZkJp5jNx8YyYzjhh6zRmmu
u/MZAnT9i1JygYMsbmKdtHfOs3Ekb2Yv2/2jxjl3WacABHAzA6uBRhe4ru1qNdegxwQsqGYuVazS
N6aUM8PEtwamnV6XCeDM8ydO8qfbLkirWVy+2l/pDQTe7+vu939D8oH5WchVsvnh9lbI53HAsjCa
suLuTlmMtLcPC7heAPm1F68BGw2iS8wjXhZRVFa8Owt9gBckt8ygxLJ1EeuIvSWSoOA+ophw8qvd
uaq4qTe7K39ArBadsZVgWdQyyzkkpWotEc6h5vBT8/anYeGjb+2t6bD+q/l2O9e8tPnrZyY7or6s
Ft0g9qkJ9H/Q2sntGrgBGRoHvTYUD02ZifEGqUlYtx/9VAqbj8pq2yuYdj1lCNdoXMqW2IvnuXv3
X9f9VkI7Sn+A7A8Rtqk82w7YlGMwmf66/bsbEhQVLiua3k62xhrnmyFXx0BJg0MWGgHn+ng4pOnR
8NU3zb8iZWDhQkvt2pKr+cW5YHt4TXvihjXI5ddK0J7bKhK8v4zqSn/IzFbr031plv8IiaMK1tAO
pdWWG45NkHetK/zV9BQkvK5eXC3m7Zs1O+NtzjmhB5/0lcQ4jsevuPBG3/oGLHWcUAUDPJkMjIeW
Hf5x+hQ5ddK9mnZ05n5y2xUQDV0yRxqHYh5lsJqYquz30cKfhn6Wy886h5SEiURBabDgZGUP6Ff1
6nWE/kfowyrlaI/BGg6xN6QGSv/8ljpQxgnoOrXsXMYeazHVAWycVzk0axqrfs9O7G72vFBpsWqg
l+SeLUktLLa+whrxyeii0Tf5Qmpse0wbbZTwZlMtwJ4ugwx12RdtTHEXfmW9UdKFIxNpWSSM/x9u
uyPZrQc1VNUVSWvuVdEXxFYfqnhpE8yegQxKrl/0V9muL0AoW6UOQOB9O1Aq5/NPmNM25yEKyTKh
kibcSVh3bLwH58LFDBCAarL3g5BuCrqhQQt3v5da7bZq7nXJnijZF474qlhQXL+eKrymsK6ZwlHP
N0ZZbKhEcbObeQwVN06SyhBa09y5txPqK0XBmKSEHhuH244MfyGudY4vcMEGzI0Rvk2sL4ab1uJn
C6iNhoOSnDRD/IYK/urccBAD2nTC/i/5FMDNg+m7/OqMasoWsiwDXlJX1hStJmm3T8GN0gz2oDNT
EUsUCub6desisAYp+RtaRCwGHw7vwBRSLYPGLZd5jRtF6yZPFAQ8O0MtVLaValLaysi3i39VaacH
AaNJWhcS439PQGqmf9lUCgGzTdxtlbjwxevqbk7rxB157Ut86QrOYsC1BpgnT9FilPPq5EA6MhpR
glxuCO7ia5JQcfIvXOhtyUeZfgNoYl4tvbvPYCSX6Rf5MB5YGTfdoQK4h5OLe5IZLeoavnK01wOa
pthODD4ynq1Vl/N90p/DHbdlTMbgPoBtl0sg1A0gFNnZctbGWUL11KVy1Fjc2A29mJJjWv2mMYqF
Pzh2HYG7AE6uKn2JP48KGQym1Q9N3CNgYWok1tYVlxKwlh2hpRoXMxcorTGascLihF4WqyaqdTbP
JJZD9GH5BAjwwwJPZuz8dMvlrWdM74JdFzeCijB0BcadoG7z7LlOnXZz1NDZXNO6hVP2DSPdmr0y
lCG3qUJ+jVBu00xF5RXjwMreS7tEMvC3XaimrD68mcT9FHrVEy1vODoz+ymcRsBPBNy/lVpRU5kI
gy45dKUyXivt+/Ef0VElk1uWPgdINc2MuAH+698AR0ED0IOixMZQ16Bbhz4fp4MOWoL4KOSTvAQG
PJt7PDSQdzyJUkrWnmEoPfF/+PD5NsAhVzCaE4ToaDyCCnq9sJGcj884nhbDi0mA9UblfRhtHu64
04H3uM6nmmTnAmm5JjnlDEb7xAGpBXOO6uWZ2LfP2dGRfLj15XOupPs/u4UipHtQqwbswVG2H7We
Xpf6cM5/o7ncDyj53dCbcLmVWatn72I0sUT3ugIJV/AvySZJRnizi/47GUy914rszTTf6al+lFP9
CyMT9YlQWLgzO1du33ez8Qvilmovr0JsJgV7bhiVGqALqoL7+0HugJ04qaXtgMHwIEBiLHY6RzEi
5eZQey/DMs154CLXCo62Yq/08purpJ+z2tg5NDEYvspout9cpu4N+lwCSOzthtgLUm3BarbT80rF
2csxrxQiM9GktpBGR6wFqqZhUoC0A1zRE2m9raKDyVj8vfXrXGdQVcepKhxRbLaXaNBcDAELHs7i
fHNwkXEB7CB3jJ3mnailZuGmJlu5KKxN6fIfOZiaBJulDg55Ab+T+rEQnqMNTsmcdU02qhchDxw1
Z5OT/2Bz30XDcqkNFRy2GkqIOn3LF4zCB/UgBDCiQm2v3dcnD94eMrzcnoGwyKv7Mve9QHtzh900
dW3dLjg65Yc3PSOw39qghT1+wSOiRu1iL5+QnAZeZBSmhLZoQdHO6P64xXHXfKxWFvd8TkjCQT10
iIc4u/emgm5dHRWnTnJKg0+kPcYbtdXRfwaG45E+NfjKls/vK2Zd9b6zh4CjLQzE7cABeXTOy61v
5zIbnxanafAJQkgu8NtSK0ZzbindkdosJzYRMNDe3v363YWdY3WI9rvF38H1gc7HY89clOYamgYF
BQa+/RbhF2yXjs1PC9FInz4TTWVzFwNrwb3FqKExQ/L5nFlbkJ2wLEjQorPpse7Hhd7TGjgT+uzq
EX50/O3g3XQNwWZSEAAEOD/C8T0ZDW5e3PonKTLWJYE+iVlwnAYGmG5EBPa1ZjkIeF4g/M/uP0VQ
y0iTdxGGwXO/dK2h6ia2PjSa/rnjRD3yw/TkbxvZ6Wg1TEuYqEo1sI8/2d10oJyh2G90ZygM2w2/
f95JNGl2qEDkN4pE6Yps9JmhfgMzhJgV3IbEa3pMRni1YqR6rd2M9/A9Sih0EGqtGe03z2xC5plR
t62Xx6X5F0L2JDMQzFnHNLb6VKQMzpl7jpEh0wjoTnPXQIIrV6OGmO9taMZ4H3pLNcLpSsLFL1A5
W7XP4f9Aq0wNh2Ao/2i3qL4iPabcBPTorJBa4ixdgDgg0GPW0ToPNPBu2XpUthzAaNonllibjoC8
4nercxkGyr7jrxc1psFiNioAHPXXMfHbbn0MZsE3vkhJLNkhs+Js3YuWElF+W41oXwq4XEdHP2cc
CzoHBUZCDfZ4MWQTI9lyxdcV4DrY3eww3m/A73ZhI/Hrj2DWkZ0Fhr+liw0Sq6jNYnP+k3iWSme3
hCOclSDm+moDyxGWIFunHCxOngmX/esFsXwQ6n0aopSXD+llJv0EDyHABxAwkMhjnRuz8cR791//
QIYULWRY52oxUIRaQuEzFCeRdtU+++c6B0a4OuQUbYhIDaG0jpu6CJRGlfxhNe/E2LP2ESOQnkxP
gSOF0A4d/12KbSFn5nZ3OCIJsijqZR1cy67ZSBs4lSZTz00UD9rntMoQruX5GwXRy135FB86Ba8e
QCF2BOCnF8NKjf5ZHBDMoXrtYUtivJBGK/pEOwgEgsXjDDvdHJk8NpPYw1V/fkM8wqVwK0UhLfQA
b+BxpdUcea0Aa+gnON0ZVD5SNvOiSWB1c8PA7SPJH023g2mFCNK+K0/xp+lXF0Kjau5nnEMc53kz
2t5qf06eHoPTE52hWpuUZWUzNWZma6bj3FYLhUok3tX1iOy40Bwpv4RwYQK4/z+ZQ6QqoYZOG62t
qztM6q33MS2je8IkYOXse5ArgIrULguEVmtavM/b2C+1/SREZQ6zQVpnujhWTY3UCFOc7frOtaDX
+mmYz4SGXEVVUc63PzDVAj+5BaLpRXFAqOCsbWV6e2ayLC0UbO4C/r1h2o3U+xMt2bGHmMib9m09
FQoBn1Q2/MM8a8gYrCyB5xfSFwa7xT/uyxkx8vz+GkqploZ0y59RqDg5ZFILXofXWGVRakftdvtj
6ySGAZ3cALP3geZJV0DhYdemZYBjUT6xSx0b5J+zl3gs45V9LSje6fwAnEdQlAzlRjzt/lDW2iz9
13on5GEZNScIGH7CI/mSnPcWN2iBXxIOPqCS9vAOB6GAjVynxugMIi1Mmkn4wSaKeU8LcafIgLs6
0U/KmoZynWTi8VZ8neK0Mqq5l5b/FODPj2Yx1uBeIUrcO20W5GhpNjO7XRDrxTfsMe8aqkP7zTyp
jM7/OyOLFH+tnHJKfhPSUeq4M7+RuvVHt4/qbVZZi1zYNRWkwTgO/QtPDgRN94RUsscvpsMCeEfV
8koWpGqLMIsIoLRmgESmZ4wiGtB7ptjq10ysObb/fdqC4WYV28NiAs7iV0I3zQS7Za/ZpDAo+v1c
OrFzlFrSLW3q4GvF3u1gMaPp6H0a5g8FTAJF8YHH+KOGO/igXr3dsM9p7zst9caLuyLyKtyiMWsW
WhkQ4h9c2ZPs4gQOiVfHlG7ult7lYZeNJipPicUgdXTMBFnbVdPf6M1+jzo/OtjXkL35Gmu/BcCZ
Nu5CEEzxQV2Wt/gNgKwhTlzwurbZqLC2JslSkCvSEHm+CYY+g6j5LtJtvFacD8nIpmBTNZOFn/o5
fuePxzfGqB6ZqnbjOEeAvf/jfj6cCMPFSIDcCeiQ+CcQtEuqkDtmzeNgt+xttYlycSHlvPCReXik
/6zph5F23MtImwBk/pQMUqJ7H7GFs4BOhOHK0To7ebPapFAM1rc4O6z47qCKg/QM2rB8f6BjogMg
K6bTI/7cZa6rIQJM+46kVoYuWCyUQOfdlUYmd6Fq1HR47wuz6PKLWdEdUkh12JZhnorzETDWRUIn
htLO81KOpm6mIaaYPXoQsZfnUJnBOuCCfgKrdtUgfwBJvqNoIgb4ZZOqWjj29YAhOl0o01QVH8Q1
Rcg95myXBfyZxMuHufHu9OqTmXmcXBIPPkHfSV//whhs74NwycsYMIYr6UaV0VZSKf3ps43/9gl9
Lqm0qVvoDQCkWLALHzs0/3d2/Fek6NBscIn1dXtjVzR6ifCg6ltFyC9Fpe9OzXekppyQ27wT1Anb
zb73q4DAXCDGcdAngXoyGMvx7blC2QhgiF5Q1drP6hH/W5KzZ4XvukrHaGl2+mvvwkb3rvDfmN5C
vBmmPYEBUwMNauK/zd96fIpiQ9w5DUJMl27IaOgRqUSBERG36qJjuK/eLqR5w/nyS3sqdyhW+4fp
EBJvewkv49rNUwn2Y0CYoQppQHReZKBa3105OrcdpjwbKWe3XB3tEQQNV6VLAnUt/FG4aCLwrMCO
PWNGfTbDWpdWFj6SMaA+9IRyuVX8W4MwdlH3TF0tAg2EBM70TU2MWlHkOVyA+9Tv8U2cjaboHCHL
ZqvPvYAsdDdX3mXmWLw2+G1xv81h1s2mNpQ3dazzGYJ+cjLQ5TfpCmAw0a+JY//DSpn+Lc/rKIlc
6ymb5t9PqRkt/9BPT67GPsUFPJ4f8dyuwWfZbXUXpUE2Wn1VCOx/usMVsgoqHs77pP7SBy7dlCr0
rU8pLpCmYde8tNXX5H0cR76NYqx/oSj/2YxGWoF+2LClIOvEGO7fW91kDsZg+ERDxz0nPnkTwxYo
shSEcAABtIdcZh4I7yYK1dW5JVSUcOOzbMLnkqTiqEtrcNdjUi7WFUehRuo1ySr6uMHwCYRB99hh
IcE4SPul3BR/fewFAfZ0hnwbW6Ygwuk5TLEst/Iov3EgJrrnYPY3+FSZxJ6vZurlTfOUkFHqRo4D
xEDnIEEohfD7ZItpFE6g8YQ0h4c1qd6kz/NM9tbnZywBrXgeVtZfGZgjWeqfKQYoWVgO5QKqv9jr
26rKt37lYy22adDTenzVgmOn2SwYKANG50dw9FnqFGcgbST3TclpONMzqWFZhEWuKU32cqe+3QeQ
Hgg7C8/NY0mI70NubYeglZ0HLbAwzA700y3YsUV1exYZkEKXgrelNWiksm02ipw4KuTT4Wq5EFc8
mqMp6ThwVaTSXF/P7RQIi/AHeP7fzfOVHw/h0T4dXSZj/tcRy/yB8EGgSSSrpS4hpum7J+itBbGL
CoP/57Zbs/B3C758bZTqZCNPTffg6UJRKlb1jbUpwwOf0Lcp+guCWTxURrRUHRYtM80y4Zn6l2/t
P2OLmBmltRmcrZfSNpXvhM7G4TstHyOZZt90tO1sQAXXAPp++/YI/m2DhX9E0nynPPfxDwDaUnSe
u2wGip/iip8PbihX5fFXENHoBGJMOvU9pf7niieCpO8XnVRLmoepKELg1MGduUEEWuhJM+kQElaH
ByiMp8Vq2a5Z74Y2FFf5P4SAw489E07Z3TUGppoPfIOqnWY5HNgbegy5MRqOVGQzKfQYbiINe7KE
en1cBSq8kzySAAufRVGchmsQkR2WWF7E5ZU+xfJ5c7FRLD+mxgWw0JHkD9QfTXO4S7/dbgnKrVJ6
zXwNEkh4NHM0NbT/e8YjYP+Pv/aORwFphT/w+uThDs215oGaVemnpgY/Kpxu67MbOfaBdb8M+hC8
ecGFg4mB9y2NnqPlLx59AtRWCcUODaivE9q5P5Y6Wmz98xI9GMSTHwK6SWIvIrGSehpaaIoxRS4y
0FI+F+JjSr1oREK8mchUR221aC8ZCSSO71ZRy0u4z0T9epg78T8+ZXtDN+GViJJmHTzvmyazl+Ej
qPr/h3vm/jiATOozuP/bEEgXaBY9nmC8++beoUG+4yDpTj1L2Rptd/rKgBW+IGGxsazrIKd3GCoj
je+EadYZj7lwlamxD5JsChUgzgj+OVbGDEbqTYHfLaVidtKK60wp+Obq0vvCWX0DSy566l11j9qY
rvGPEXvOvAnsaUmLt9mm5332EL0wUAdkH64YfJGU7Fx4Rlr6WyQY9OgDjdFTD4l25bak0QQiFo9r
UDQmL3v+o1K8GAl5VqD1rk+wrPLqLIEada8uwcts3XjBgIV9VZjMMgRkrJyEBM+mL4ALfE7/BPz4
LMZ8IJdLEgOGinIjPxI6g+kPTUBMqpSbSNUEbpWUzfEDkmYIO6mm+E4lvG9QyvMZxT9ciFrM6Od9
rvQh2TyFQ58hbqoW/vwUwjilcYwaahlAxBRCDqhZ1kztfJFjSpsoTSLESGW4hs9UXq1cNR3Fhp/e
5vWNJ6xq7m8GVqE4v+tDTLcdCQ4C/Vd7MID8Pb7CktUrOGnw6Gun1kK8vD1o0dOJR44bmOgomah2
j/CrLrRX449xUk7kYh8pfZm8Qh6hGCx9vlxhX6vPLMPvouuMAgCnxfI2wzrjfutHxkuhoPr7k0Yk
WG79ejJCb0Jna+7XKEuNmRCmCzFieSj2+siQcvaFh2HbNqeoKNjGinBbc2DkAUUj93ANgDaaNNJa
KxRKo5onmAz8vRJxbxn1ghfhYAOmnzZ3b3eTKdqZlQNkazUhEnyI/aGoBLKGexDTiGyzeZsxU65t
fOTfzC3pSaXfl9gGuHpTVDEdG3R/fmKKvv+a/y5irh5dZBMigZg5mfixCoCBEqOnVpTxSRBDkpDz
Z/oMeofNIDC88hus+DIMOwchVSes8126OQSJkiFEX3y+rSE5fxnfa2kl4QkQ2I7Nx6MdXIHTVXC7
yFePDzcJRO+KbQBt78OMMFppAKMeOjJuESporMHnok0PiMcsUAkv6mGeamYkIjEY4V2YOKyKJbaL
zLUBz1ouvrIZfh/cJMru+RciqqRHVn5uo53b1pwlocKQmGgbO1nbAUSSPuESlthfIXVqOGQaap46
+5q9o3y8/Hxc5W6g6xnX4P5IWk+2TZxBmGsDIkbG8XGrnuNapIlQP5bp8Snr0wN5DRNEQZb/eOSX
ysukzL4Q+kdevRH+kxOY13VXvYzzzI2gVX/2xpBGEERIsN9JkXs8A3e17bRe7y6bU/PZ2Kr/FeW8
/FXLvA3ywgtJeSnuXnFHLligxaFvY4Z6L02abFCCkTtqS4HM7zOHyZCGftqM6+GaExGLPw5Uav+W
2l2z3EgvEcdCphZXJpIQVJ4BZW7mhy2fYTc5SbsxA9bsxk6Tzomgv796rk7HvaMU4D/5J3Y77CKC
T3bXDwQhwzRUwFt9eh92c+EjW7FYiHOrpberWObHOhYeXWcbqb4R04aMc4OL3odBIyIgpw4UGgHG
5Tu4e10FxqcS57dj5sFbipdo84orkIoQhprQ74wKXbyhoZe99SRaRsa3QnLnkZ2f7HessaXO0RPD
x2kPBCOcYY948F7XKeu6VGmjRzrNtm2Wa56WpAxYQgNkanzG29o8YAgZZr7tONz9UafkQil8YZRN
/sJLfL95kRvk4DS+5GYEHdHRNSrf8WnlVIjhOvpsEDgXo0KbLrTHOM2GBDfkBdqK0LmbvF5bk+mN
rOQv9qtjGi/Y/hh2V4kjSmioOP8gnzfsd2In32aoY9aTKEASYGgw3UK1mGQYv0cSN0HXF9D5sqRI
c0UKmjuRk5h5rIFHiDKezsyvyxgInErxIYXCeJ7kKPghhU6ZYNuAKBfAi7Y2bPUVzEwIWAYzNnvg
EqgRAgT28dOtE7sSX9pbeCJOuVY6dGlIypCef/NCzNpqlo0ql/JR/gW/c8RvLwoWvvoj3fxUIbCm
+Z1MyxpB0EQaIMoaKu64G8WW2pEUCrcC15ajhwmlLJjLtalMH6CZ5a4FCjOdGe/c0WEbtg7DB5V3
QEkLqp7dXu1VmYRS4/zTFnlNpIWaTHQsMLD0CN79u0qJGjwH+YrHdnXT22OyMNOdwegd0qUX/LCL
AWCcL1bWkrL7ucr7RuLvL5DzJLUgnrWSkwNmVxg7uppPNIPdvBsuToJ/W/n4aRvRNH5lfVRs+BRb
8tm6ruy1cy67YV4sOJLaEVgiuXLW1ZsYZIXakdYq4rcTWgGO9ov31af5UTRqGY+s4zWEM5GGIxbG
1wrBea9rJE2pj5KR5O/3Rht39QQSZrlGt/HPunFD9ulvnexmQR0teJlDzs/adrWxz+38aUqm8rIE
kpd7mx3Y226wUVrbRW+jKSO1FbkdQ0w83VcDNu+c0bqA7u3RBBsorzaOtgP3h7uQc4ufc5XcL2dz
UDx8E41mhf4Vh8sHcCGoI5/9zbjbUoX9OtkvbiXlxzdC6H2XN+vqucIcU2oB6nI3ikKVLkZwyxAT
bXEP7w22y4/R4Y9Eox37itWwMifD8H1fXqnX2arYYBBqn+iyM1JuEgf1lEN1pM2oc2GLL4QjjvwK
laMnc63TcpVh6ORwUZSsqJIRj+a3DTce/77We4ie+ig6IxpsKz6qtZcn++YEdmbLbDkIoHlsVnD/
/u82VuxttzkWr5Ce6xVGYSJd4/poH1FM0IL4tCw2sGEiM9ncsiCGwqZVL507etQiXwDYKws/s5KF
vvQzvXjdGqFG23IhnqCPo7dywSsARl99cB2tbkohcfo3tRse4//YWMmVU/8BTEAFejUYI3Oe2G0Y
yhLsQ6Rley/4FBlRbDvNTv2pnaApm6b7EpJ4iMsUUpveDVU2tzBvTPeHOHjcZFmIdq5oDp4i3HcA
TYTNyPO0AQACZ+H7j4rfvC/iD2Ylqbere9iL6yA4/eOqQEKx5aT7P+2vkxQDwmtBi1vXXc3g5LhG
ThMHka+R1QjITFThLAgk/qEQrLSt7BDZZ6iPtPusNYdk2P2ScnZRvvQi94+dFaLekI1DmmR9UN/P
nWBdmlyFtzsPWr14qLeejCTLrg/y5/hCygo1DLYsXGr1MyJ5/H9XBzDjdJISBpeMpwwwSYs6PFIw
fYGga2TadCdaane2KeUF8eShJHW9WrbDs3AdON/rQRHhWtUlnFIcSpMKtLP1Pxu5l145hwwDTV7M
oo+be6pLYe0BgtWrZ5YuGbQqYFhIqilk3Y94tvWZta6b15MuI222SILz/ugO89LDmYUrbrgU8oaD
8uFCV+knJvmCP4a/FNLQncYJpp6Ezv3+jkIWTleJ9wZS5HbyZcBcebFTln02DM5qnty0zX06x6zE
McQbENCKXqkW6nklhqXaIF2fJdjc2n/CTNDKNrkFkA4IP+KKua+kx8o9jitG1GXa71M/HxsZgj7X
8DMo/iJvt8KDgbpmG8X64XXgyeTJXtUgFKVVtDCqvfdBd4/JBh1xlw7dPlix9S6jDlDsmqGqytoD
BhpvZscvSE8kjUhl8axRaf9Ameozx1+vYr36plHbcRmbo45eGyEqAKsU4u31E5fOOkgmyCN4jxfP
Hc8JuFVkYtTd8o6J+LTE7FhRqp2FHj0sWpJAb9G2JlUsBj2D5vstlbm8H4p6gaOrOc4pQa/y0fW7
6dYJNfJd5kOzFMc/uCzK/ovsYzKoriP4RNMXGmEhhG0ZHdwPZi8oy81j5582lGb76735GGxmTJ5V
1wy7bZzGrJ3oIqhX4DzphKYv05IkziuiIXEKQsRz9Gco9aB6Nnw+3pG+s93NDP1kY+iVMsemdybk
rSC0hGyDjBFPMxrLs1DeoUJBxfuCDafxAlSnb+x2yTpUyLEes4nG1zp+u0YEBsnEzHKHfargMyh0
R1rmKgbwMEHGyB3AhjbENiOElgtkOD9XlvjIRa8igrGEPuf+M+9ZccsekhzqExqFRMQnYSao7BHL
1z/oP5IV6M+nxDWWT13Znyw36fXeShFUvXNS0+J2cypdczaLJTKnugnipg44EH6w7j4kH8x0mLUv
TG9O1tqT2OyrCN1dgyRU00Q0GfKx3kfes6Q3mtJ3kryIALGz3m3cZnX1EfnMAIHWhRLXCjpIicIr
tVEXIJn+Lay+94czT/pI5Dfz+rzL0rxiZIw34AxcuA9FwSAfI/I1UuEshF80kJuF32bW/ntSNZug
UhNYyOYjeIkDmfPq8bBtvkT3/Hb7ynQq9N1rMQwVjZ+yBnVNI046amkAxHw8+hDT8m9x0Vom4ePR
jeSDu6IxCYZKKQq6ayvi1fxXaN5qIXz2HwoTEFWLuEQi/kuqWnnVyUL6wo6bsnQZEqkoEUzQVwAq
97v+jchLXidcMs79KYgUExrsuyL9JZ2FqA7Jb5EhGGcLl3NymC62K41kDs6sgCi0bnQF8/0r/z1z
Fo1n5+dxYQS3CGMd4ZcavUYGgutPCoowzD+/oHqyP24PbAGNo9S/eebvccH03Wk++xQNjRPx1vXr
ecxhT60WYCPwn1j5tPnM/3hBuRo2nNoV8njMI1uGMWDYwMm8Rdclziz8iu2ZSStc/q6rMl9VaswN
OpUGc2q5dSGq50FbxaREXvOOA2/x6NI/INOqFWA5mhNwVECNEyMz3aPKhVry+yLiZQUltgvk8d5U
7gDLGRhLt1uCwB4WMduASFq2/DcJceRjLy2buRpUnnpFqvDN5GdYq4dJvIimMC7REoIjf7/d82sM
A1VfHnJadWdDyavcoiMKJtbvQIZSoZmmdqhN/OF6wUdS7OikvXxQlOpPWmfXz1gJya+Mbqbky1bE
0Va2WscLtVeUeYJ5onFK5ifR3JsTEInzUwaxGaprrri1ugktFQx4xfGWOd23HXVxgUxJryNwlaeH
/IFt3Lpozurfy5Kn88Txkb9/lCSILObwjqMemShM+bTLpi3SLDfq7veO5Q+Ear/5t2ihIiT+MTOB
JV6mvgzglNJmmMbltn13mF9DsGUFQsJyZj+a6syj1nFxkGIC8A4MWuQUcqwHXgrkaH2mlQXCMj2l
ttYakOha5nVzBNgvzjaK6vEhfppm5xRV2HAdeP8TTb7fZImwsPc3E2KUy+RRYzNwaFpbE9cDDz4x
J9bTb5QGKSufZRdRL8wIM9rZVW2pN2ZxCa4E3wu9r5ym3XOhal23h6q629PGxHQJ2a9IGyhiQUlz
3HW5gmUov7cQPKa0g/+LORgJF1irrKbTuygxpGJ3PSBMqSP2l7jS/OZiji/hGj3XDJS0OPS6dwG6
U3jETv2qabNVxTX5gv5+PDcaNSJdrGQXX3LrQtfbVmPqyDYOCzgVolLv84HPB+TeT6AFrnb8BUz0
eJ9li+qvSSJiSK/exDU5QiDITGXTHfLsxnCFWqlRyO5ZiI6VNdDxgGvKRH5wdorGz71//Bd7kpEh
JL7qOcHF85IluHXheyxI3ZFEA6d8pf5VUdabS0q3oNyCxavJQP+cNMBF4h9rZA6o38+bxL/H+p3r
T4h2KvmrgNGl6g70PIkDMrI1VdjfYIdFadp7zAhT5Waroa/CQ2m4XFu6a9tqV6sWu4D0M12TQVSB
tYnZGvcMcds3Fc4KsDbkKD4gnrWE6oymZjjHGew3fUh0vt1nb1HVrxGHozqjzbntdzZr6GvxEWBi
oZ3PlFx3mDEehv42I/C8LUPeyV3BVUqF/20GBqDBlwHz8jLEbGv1y74gprLFJqJnAVmmnKyE9qol
+chcila8B5BzHse4aas9MD1PL00CkAHsfkdXGX0Yjwql7+LbvBr728n/aGkmf+0dAf8+wHXUB8bf
Lcgo4q72SMxySfl+TY0sIfFHkocvtBUe996cNyeTiRAD5Q2IjMeZBNGDEjIEjymfA69dA4rEEAuw
Y4odMusHNCrtSHn+FvuFVzf1aWczQ/lB1xNlsJGFfk+NHssegutklumYoHgGWtfNPEFg1j4HRpAT
+d7D2+uOaLQmpYXVCQdlvoLFY6YV/bCW+VkkyDlV6iAD2L0jU6FFi6tQcVtOQT51VCJW1xTRiQRK
mXkY9uVI4eap5fUK46IwuWTn4BZWkQb5HYEFIrc2fk49R4RVkK7vAKHTRuCC5jEBDUuH28bnAZCa
iKbDY1FbjgS0280i1qRXTVNYpVILKB4cQcj1pbK8P+T08NmFn44Mv46MfVCuG2JmS6qBG1Kf6oVT
LLTLhelC+1a6I1SqYLzIzFqG25x+nHSaUAC5UBTjZrVYuMcRyJjp/Z9Me9FeZj1kXCAp5b3j7qNk
3kSXqRFFikq+vKCozvOci1rE1pSRAbvH1ZKZfqIROY3u2itgyuiQ+8kixlW1ySQ1Sfsv903wyZBY
z3T0KWLsnUu2WIEPoedAVq3XUCz64SnGYF6hO2vs1Vla4blOUQjlOk2O+Zhx3t1hlaOpnOhOGsLk
sohTHssMbWyrDjvaIYoArWo1DlZogbs0Fb9MmiN3MjCH24AjYr2T0O5Cmv4q8eUnnk9s7Ga0L1Y8
dRmY6MIL1YdiRPsVjMknEhFeQtiJ35gUo1TP/K869GlAVo2YRMrPtTlDXBgrR18PwM014VuKAiZU
YDMzYyrZgnt2dS37uFIjBcPf2RoyhcRate6TxOZI0o0ww0EFSNX0rYSYJSS7Ib+VNDHlX+14O54a
bPulrnAcuaheqWXC3onYRlgniaaicap+HR+SUBPXr2LhjivNYwO/3/9NXR9Qu8LqBd6JhtcyJru9
XA9pQ1hSfqNwBEajAYdAkUqc0IgG21cd7yjs6iKNJKhF6TV8tBPdjFEwNgGCgHnkok1qBE48FvwJ
vTR6MgtNmJd5W+qy9avNrURhtgYRJkbRo6CHUBjWl3XuIPdEconxVNtbU8bm+HEjtZkLDDI75STL
f4Bjb04s5D5ZCmlw8r4rxpXhbQYRT9sS5WDiSsoa59FQpap82bUFJCRgaUJhzmKJY7j8KUGQ/vIL
9mMHsLkp2rj5zaVplda2N2XSz1Co0dpxFKKxz5rYj6nHijVJ9JGqtG6kaMuovPTLG5CPhKMrtc3Z
QxuyDMt5fppuu4+ivVT3UbTyBMognf8uhpVY74jTq40nk3wB2VVceHjLi+eYYr3Kfx0PHM8BY46v
BYAHavkX/I4m4/RZ8tsGsK6Sox/7PTEVSRcdc4WzF1wRljbj3KnGwDNW8+EhD1oWoNmGvlWvsllh
FMTcfw30l/Z/RpFt3kJZb9mnumR0dz2l2Cj+VgRaLFojVdifa99gMkOkaSqPIq9kfpzpSNHl9yEb
/BSktRJ5kXBBi7zq7BugpaZh6IcQip5LioEhDejbzZYtHxyob9lSgrtzIGWekn6gp2aH9uMa+8ZJ
sJhJ9dL+0QhOQdK81pXEGQFARDR9ZYQHuz2D3squFEKiDOI18agQVmeClwEICSLQhHr5IRIiw+fF
+C6ieombdba517NfzZg3Sl9pPLU9gsKnU4StVczpFqPfCyyRUoOhgF8IE98eMCNm04jITItzrn7+
/vHp7psKRbkz3Pe6UQkVv1yBZikyWx3StK7wpnYaiJC6SJcdxu20flvaX+5L/o92wVrp67/GmXqY
xNB00Ip797LB5qIOX2WGF/NwVFeB5Xk7nrB+q8jDltAcI1Ok/2JQx68X0r1u7wdF4RNe98TdmfuR
/MbtYz0Y3e04zsmveFHJquRWtExzqMijssrwQ837GF1hzL328JxJ3VBR8JhSkQ+3aW5epySqcrFe
/xQdgTvYsi+Eog7hzCg0Z03oUXEAl87c5mbpYZ/gJgx8z1AoxG0vnK3FtL1qMxriK3ZXEuThCpEd
x3OerCiaLFZ0KIu/5k7NY6q+zcuHwuqHbp+f01kE4sCKS1aDx8aprESg97qWUdGa1/wSmTc7b3yL
co6DNQjw07yMNYnTjSu0yAubzltFdWc+jTfYQAllh/Dfg/320dqt4EpH93XtWDnsh84xkMaJXCTl
ViUDReLpH5OH7Gfft+O6WrDOkvr+7aHXxHVezsD5dyaTTROMSx44lp6ubcy2tR13/4dkCGI74jM3
eFbK1xui/XQ2s+mcue+jRHFYXMk8s1kJ3CBqkKxR3FBNfgEJs2u0WbLnh6u88mI0fJUfc+kLzrkZ
v0iEwzFxYBmlGX+/VaLmxeg1Nv2mZSiWM+vxEJhCCH4VjzunrrWToY/pFO/5HeIm4pU9ZApf1LUj
tI1uOTxc9BPNViqf+p50sZOI4Ir5Y/Ytpn+Vu1EQnvFZzaTuepnSKmfgYJ8N5BL694K3y0i8Ik8H
wqkAkHJNOisSBmXXqDDb2ak6FsaBgHCt78jkEkZcw5vUBiOBaSQ0UPUwcjc1YPUsHfm5/aosNFWA
US1/OjodyUkQnMJhNs4+eP3Ao8fGAK7lu5H2mr+nEFLQsoSIZZ8nVqTnmQkoN2R8mGBOCeCdsBhL
N714IIMzbU9jtgFG5DleO4BetV5EKZWo4sCSJg4G1DdcZwc8fNkZzWVDWvZQFU3tNmdb5t3Uk5He
Qflq/LIVBJ3VEjddd8yBlKJB4gC/EkD97fgVzXlrrKRiTI4u9uwbcs/o/9LeQsLignnz/zz1V4R6
BDfkJTHAsw1In4VZ+RIOZ3pbTm6ceWDhNWgKIAYU/7VPTurTK4QhD8jdKMGVB19CQPQwDErXht4P
LIoQlmvwj7wByBkSmssXADPQqe9/2bC408bTS1e2cXxh9WQjvImy2Mn6THbV4DVP7Py1o8pEvzy4
nSyawwensgmwOQQJEFMP0+aLvx/a+adlRWFIjhCkrEV2DA7gIeq0v+SxdUqEQMYF6wUcIXB33spO
RURmUNZst+5dSce4hWvkFg/4cizOF0QEcxMvILB3EjeSZiqGXrGH0PF4OKQeUCnYvJQg7uMlfiWT
ftnrl6/0vLRjhJmGpmOXxPUgq+NVZj3wMXnh3vEXaWGHaNbqiFEKJHst89XkjGVaqaNJaNqsZVDN
oAL7YJ+R0Pm5RC/VY5mE3hMiijljBftE3ZgIjb/6RDei4NQBQvcOAtfekYbng/fT5/mZMz0SiS8+
CpbWeeX/CJDp1Tn1apgbSEQyZHlu8FkAm5UgmI7UdWRUix9F0C3cxLMXkvzyInd+BkcvPP7n0Zro
VmZb/RBMx71i5G1czcfw+6wLVFjr8atkJtbRh9QjUgvd/nLYyHd44htAJpz5CFVRu6TTQJrLXXQX
kVA6JTHfGEIEeqnCHlmhaEheDHtZxiADYWiyntR8+V6nZPj9lJ7s1ze3bsXOofMoAM5iDpUhcNcH
oeT939+tGXCXii71eiUrLpUjKUx02qyX/eCyvrJ2m6/OrrL905ozuJUb4bOkPTlnlNUOwTlck3Z6
mVC3NxM0RzCaRnTpGBNfeGNTddva5gkcDoZkhFA31BMeRb57eZXAAp2xjssbDZEaY4chQ5v4M01X
MVD/M0uOaeix1kuyj25BfSxWZS1WWcCClVDSdwqkmzQeBhAh1ollxksqkyF6k81MfXzdqjDOcBuI
1gQpwJHbCWdWdZo1EZHA0piztuweOuo6t8Qsg3vZAaha5dgB/jq8FG7AZK6KnlrVXNfVsrCy33bo
R8AbLF9/+IKewaSSKnEZsnfTdF2w0k9Vcz5Gbr/98buTnN11ReiqgciKOUZrixQV8oB37JuIR8X8
YtAplcjf7G5RxUsUHMDSCriL4gYvWJX4GswhnoG/lTKQ7fRbrw0Y3qlFzQztUEbgbaDY9Y8pL/ak
frdbrQKoPXxgaMLSdOmMWwNEE2jnqJzRBd9eiXnvNSStp/g8mehx/o+qDabnj0sXGhjsMs4MaN+z
MHqnl4oMx3b1GO05ebW4e3x2uTfsUh3ngDvEdTMjKkPpFZavBeTA1uoIyQDlMUEZSJaLrmblO47M
g7pqiaXdBVP13hZpAmqOY2RC8EgnqG/V/UBCS80NcFte1RIFM016Rfk7jJ/KM5WX7ATSSoMDGdhy
DPtpnm+8k8qikV/lmIuha0pwR7sgQqXJc5W+ehf5fjwuRIOKXJqz1brZ+dos7eJDMrJ5Q94fBiwM
+W4QiHBmTatpkv9ADj0c1BtvnQnrDAFhnOugQfyHHW1auVt39KW993CpzhaAUcIaUbFNi8O4SS5w
nRWbvaFHBBgjAICWblIXC4sD4NmL5Jr+eyG2nbxrclAqJWvQmEyczJUY2EdeI5zSUEu8aCBawccU
wS4yoBUPXhQZ/ud+fkyxQfWOq7O3QwH65k9ey/1+tF+sjHBnR9aLPG293/YmjB62sAR3lYIyAq7R
rHyjkFr6OQ0qSv0088URT97NOAvivybacpqzB/Z5fKFx5HpESCtOmtqeBpXjOGhrZ9iIaNvCv8iX
76ObetgkUSAmAlphIMN4YD6oeFhzjD9WW1g94gptMsJK611rDicXtZulhUCG1wWYk4cqWdnl2Ggr
NLMkLAbCZAKkRxdq1woJgvqMcE4XjhJm8Wkza3JslnBivhD86GlRhamnxKZRIRkCy+/3uHl5rbo2
2T8Fh6gP7Zz3Y04MZPLXJJZNYkhj2VmhN3FPyHTGLsW8bAq7O0RZX6FgAs5hpJCi9hN4oq66kSpb
mM7biv7aChS/lx4BxgmQ0uLQAQvarSRZWB28Th8+K8fHRm+Eq+SM+P7wQBle+nCW4uCzhbPHIu8U
tP/SHZBd2ub7cHSk+wlNPddwi2FsRppAacxf1+DFmDI2ZTAEdaegjQ+9zELRwXwlpHDSoZ60spXD
mjAjCSagK5yjQHi9vHtMf4AaNtroyCrKLgFUvMMjvMzM1ML7JmtlVuIqDVGvIGcbpLSHb4jawC2b
5lQGjDAPv8IpNk3gLyK2EyOz5f1wsTEaoFEcSfMMtqnBDLjzzClD4/yjX0iacJJCLRQqA9fIcbxt
n5uTg2ZvmBiD3DNNoZvw0KAnVZ1CtVRNFq5g6OMzgU23nKmMXndLGTNT3AgBCqOUSolA7kUUiFrn
1uPVTuaPBy9lC8iWey8qNGcqGX+6mD0Bc9oA75Ddjwq+vVD9N12C2zqFG4HviG78Ec3RTfuW7nGE
8+8TljXR3LyfTztBcfarE31kbPZ7HHujgcV+MhqAbp2uUlUz3aQuwbkEg9W0kipUc/cEncxHhb7i
I24x3uzpDZegUr4Ihb4mAV7Ng2C5Wqb6vsPCjTA1mfGCB4MbJDueTh9oT0DGLTnvqI02X03UUfRj
0K82nLz/iERWogYXdcCylAKmq2kj8LiX2L5zAhvZ8/oHRMYTpWKTz52Y0OgwkBgdseQm732KrZ18
FJXj/NMfY24xsLddOpgdf3fsCS/wSsCwtgOSQK9V7pAY9YzfegoORNyCv7e6rQzagEfx9FpjZRgF
9MqwO4fQFtymX2lqi6hyqBphG10nTUmiABf6O8B1MWaMg4ABrHqKLGUMLSuwkx5aHOANSIawNxB1
zvBzPEhQFLtDctmP/ueZlPWIJcDiX1aCGpb211XhHYtPhoDBLRxUs28qmt1x6ZKP6B7e1wyjfr70
No7G4wKcSNesU+hj163o2D2WaH8TsquiBHEQHmzg9M05X61O+0PuoYMn9SMhn4fM3ncInFu/mW9l
TMe9ZAi4ADVxsVrzsemvbBtLkV+Ls4zLGISRY0vOTksqln7qyBa4SpfdhUGA8s2VS7PrpFvVVDFV
Dxjq5aauJlonr86X9Rs/h2kZgaj8aKMg3MhMZvOJ7+zrj4XypyxY4yT4WSntuRyA4iwtk1QdQd93
U3tMQcIerK6oIfWukUxdaLd42pW1o+cLVn9XWBl9tlOpH96yicTRL5XxNSvDd7aPXWjBxZTj99gY
iNYGcwwM9oHJLeZ/E851lhLQih8Bfhxp54+FIOCuGE5wnF1M1fiUAU3zAfLiF39nnNJxPOqNUOiG
ukyiCtOBjgGCelXBHJK2wmp+h2TRm7i+MnG17rl04kbyLdfKGZReKX69qMiXbh345bgdHJRx+D2f
ZY8ywrBpQzEFjZ+ks/5uQp93KIGHZHCwWcdSN4FsBHN500Qdw0DTnxRox9fSKQ3zHKvsi7d/mJiX
o+Kiq00DjF2gTHUGgrfZlEr+RuFC1kkFVJu2AOdZZPRCXV4OuRIGwvj88SA1agge72uL2O0CpNec
dz75PGwvUu7/W7ooy8rAVDUxNIW7YFnHzQcQLkjWcMMr8RTvPdR23ghKr3gAEHpwu2iNzbhPmeKf
nL6AqtK2xMITgA4GAgFGs6zCFqiX2M1c5fIYKCngAvVFsioo/6ppBQF5vDBGKQwDnYVOT+qwQQZi
3ZHjn65H8F4vU8FAcqWOq/QWOUAOac0TGIb3VJip89GAnmTkP7i3iNgtAinbES9fdDmFiKHk1acQ
+CeTXAABaXXGABqeFmUhsW09W9FWS/sENlWlDXhaxwyq0Dw7tX2s+7qVndgwRrZtUy4q6IXQCVIe
EwokIjZXj+ay4gN/ZbJ9v28CYe4F9lrgFnN0CdTzLti/FCuCKfghAQlk6O/nxpvii7+XCh9U7qiQ
nM1j/HyeOCjQgzSpcoTPQWpX0e1eHAEy53G4drCIMWpM6a4EJumzkhvQY7ohcDOcdxZ+rK/8UVLt
Y659KXHMXMRNGnGblGlJcXVRqbsXppx7cJQgn2H+qKefZMVExqP20Cw+8mq/jp/nkwX/WcMj81GN
KcSGTnwl4tyQnn4XmXqL2kAWQk2HTHSQcRBUqzyNeA87JJJ8zIUCWCN148UTUnaB3y60VVeOLxzK
rqaL2gWE4nYVTqJQob6vWUap+jIlp+cJ9xhK8tOcOsDqlugyDsBvoftAdvm/2/0Fykb1Lsn9vLjL
IEZbE3BpAwo12Ugm0aEb68UOwDV+oARw/H9rKt09biFuChrh63tpu5ZEZYCaXMYLtOjSK+nUbnPd
SHvQ6GWAe5vR+DNmhzs3a/daW4DVcP0EVvK43KxtEgiWZLxSc93IO36bgmeRPD7Nr0QAoik8Cgzf
TK0oOm9P2+3HGvCxw37bm+LfnUBHY7cR+DcBXEm+8aitOmmC/SxFWv4owLkTaIFTFaW1t9qTb9JB
jEcWuW0FJctMgHhQvNoZlM7YWFkICOuCcyIy1eBoq1/z0sWpzfeYFYY0efvoe2AZ8mVRJOczpR+M
rTwdGK6bc+yTl0hl0uiXIj0G3szNJ28DHMLKpO8pWgchgficfyJrpIydULJBJVmAXwdxSAZfbvNW
LSYCmK32lwBvlUR9q1vcL0d6VNjiYqu2XZsgHC6HFFTSbjzReQFd4PwJMMQxoDjfAb/uolbVbt+y
rx06AemmCkbBVRKIreMS2nieyXx0h+hBa0JC9ZjAYrSlClCatNe/0VWV2wYYPlyt2yd9h1b2HO2q
xWaEqmJxTNXcG1FD3sqjate5p8vLTFWD+fJ8avP91a9SuUBqIbbr5QMuKCOpBfT+G4b0wYjS8SnY
EgEHxz9Ulr61hjxKRxpv1scWD4sykHnI78N7zU88J2vlv7MiSs3sTZfL+NefvnUXa0T3vbFXK9Lp
eIIESRwtRSMDpfj4W5AUcAx+oNS5FS4+4nIlJoCY2stP3YGFg1I+UZAaUmAU/FajAiUMpIvuMc1b
cZ4ZocupNlAjvy4Qclzz8sSsW7V+gLLd1PbNzRvCbnP79OYGYCUIlGiFY3GiZg2McH/Qq4hd7jjp
UiGN5PxGNf6NV6T+ILz9hXWdY7qp76L89ANwxJ9s5FQv/Av16eaerQV0/Fi/DnWe0TeUF/wkCIZE
Do5bAJMYgzf7nhM89ivaMMSRvNKJUMhjdal6pyVC3KgMSsP/OP1uyPp+jBBztzMNxylG6/xdu9rb
RGnqhduK2Ob83k/VtihoXD9OX24KJpVuX9oW4ARAYh5HyG42V851CE/fP/z0erg9YiBCDGQfTLQy
uGLQdeUfapwIeL+coVODQ5GJ5hp9eUDbg1qVGajvU/af5FeHw1ZVorh/6EKfTwIVO+8o7ocPlbIQ
cc07RRnjzmIHVBbtkK4YWrHIMhVQTW0TLewPz5ysG6zL0yNhbi/BwL9CIflFk5jMNPUaz/EvtQ+j
3XWP5q46Q1F53SKQBUoupL2nLdM4t+vZ4Ru72yCZqgZoXMTDrQxFvppQ+XK9Q+9sp6Y4ok7zxDH+
SuKUducrnATaoo+4pRoxbCCHMLkOnIooiN7pDYspPqb+QweMv7HVYiVpXpIl7z+TT0ZbgR9067fR
4DbXgT88h2fhU3tfDN/aOCUz4xYBMnXJW7HHCM1hN8nWB7deQj9EGAv7KpHm9dzz6iwHc1jz0KpX
3UEjU/eTOLalKGtM/UP/nwU/U5r9UqUXpkHrP9D9IPufrgZwkVzL9zGyKH41XuAVxqr1eLv5lfUe
tNjTH0aVVGAKKCaJ/cnqolWhfi9H/HNQjgxngv8M/ffF6+dMQsn00TGfVpO8Tshmw/Y7kYNzrW3e
2LNqfBRi/X6ZaC8kkcCecT9pk2985RZQp7nBp9KZw7DlwSIvac/HuWFCHVntRHJtPnOFFmnWSRWH
HcOYXDM6SZJpbSStt5hZzuU+mdKYuc5XrUXFi2zOGRU0+VC+UP6Bt+LgOa0gdvj51jYxx26aJI09
XcJxeki2+BdDgu1IUcvfEZsLkp9FGIwQ56aCK3cXqRz2nFcEBuw8T2rCpqsbNxzLh0rgzcmL2Xtg
0ux2KZm45//Nd7JFRKcM4pqvdAXoxYhxXUAJTRDlUwiAB1ONip0akT1yTPh9YGv+Opko2x+IakZ4
M2fB7zfH+uxs0ymLkuiCxPVLYeaz1rtZy5rUdax/VpFTKqXEQp/adUflUoqjvYTSvx6ZGLhL5FU8
kiaFZEKnym40uEeuaU2Rb1WjmmjSAQuDg9fuCywjVXLZ8pAfR93r3t/QiB8nLuTY8iVGuJXJRQPB
iQv3lqXEjHQZxM9lpvgP7zHGYef1HWaPquIgzdC0IREL4THpGQZc+Zm77eLgUZYQL4sOcxARA5v+
Y/CpI7dYBf5I+EKuYQjHngdoIsKUU8e2J7D2ln/jkOZCbps6RSabAE4hOcYu4gs8nl6modQ32Gn1
wCmg8WVmXYPPhanBwnB6sI88L67QFgXV0GNdLdYQYX4OtJEzfmho778ALM4N6FE3j+YTqAKKC5oJ
4MSVi5NwrVxyFoA8zERYf2B6jFvfV6KmNoQmsDkATR5BAfcMnuXBNyHyfx019URwL+93eA8uBaez
g0R+XZZm//GqBaZ1+cucBiLuwKnhvi+x0dmgsBJpWnH73Qk9FfyGObtb4zmPfIoysOzrbg4i2Uvi
F585YUKbyz7AWcIgwtHzyk9DMld6mxPNu4uvYrkdrrVPsLY5kOqXLhU6ghuQ7L+pFLEOkrbYJKVF
lWsw1Zu9bTsVOYho02mQ0xULk4q0+A2nTB1rhx5ZCctGSBdn73/YgH4UnpEve1YGpQCA1XKs89d3
luKsY376In4QBYvhmmhwGH4CTaSltdHu0hW0KU1IxhUV9BJXmz8uJzNL9Vyqdy5wf4+nK04mYIMq
KsLrNgj40GqGY4K8mZyZV+74bCdGl8CYefRYHqJD4c7MAkKcaB4UYQWgr1k1SC56+qF5ydANRFeX
3EJ5cpqS9aD1BAi0k9gORqtXNPSpqCsBqOf9nHmFNVey9bl/n4VZc1C/AvBta67vTLAonzuoRHFt
P/9ZBIU0RQywrcc69HNTL72WdpyyIYWGxe669fm1W9SN5Eae4GYLrVXHc7H/MUOhou//dOY5AgFd
4H9N3snuDGe51VQEe1NabTq7YJpo0CSsBLU1Ccie4ebD8j6hcgihuGVxCpgCDIuQ5MP3SdYg4UeE
roE9C4Y+N7xCipxNAkQuWuiIprGwUDNJFzazd6fyn2Uj5dSFLCZebupirPEeEqNU9vB0niIW54s+
7zV0MGeDmujs9bVZHMBvyiIlHGSDDxcsaGPCtOmeeKuYqgqKhyAY0JP7JEXtL+1T5FA/VlBaD2nv
vH+/IP4mzwatf0I1rIDb5SvBQ/RLW4i+AUBLbgzjXzDOVuD3OJQLu/V4pdsNEuBg2eIVbwabSKaY
kxe2zN1mrXtZQ7J+h99sGgmW2Lzqhi9tH3ofD13+sw8ZZvQejv7/nEyrLng+Gb92Zp8EmlhJuW8d
SgBWJ/VDrHHNaDl1g6bjpucN5s494pGZRz6SUciJk19Ekqc8RVvuWX0E4cdRF67gxDQPlJvtQjqE
VOYMQCsOXkOQcTsl5KLBEG9Pay0YEP+fufjeYFMhYWYgE9+gVyzkdFOvrmzUUwefbu7O0wZOjWKF
NaKZoRV69cYpO9juD+SSvhLDolhTsts1Bo1kOpgVfAJUBnX6Sowd5NqfrOpErYHHip8tfOnFBkg/
fxuFkjeu/4fVd6NtsgJKJLVIPoDBW1adcMD4jZjm1djfZOxvXtr77uAbSjp1Id4irFgmW2GCbbe7
Jc9xHGaTgZFAeoPeMQZGU4GRomsW2LNmVi5LvZMGbHuoMtH52LE9fQX/nVTKbjwqCOSoR4CIk4EA
FciiE5nkZv2YdnwHzc/tvphzDfXpHoRMkFnS3XHVTc1LH8hWp4jSAZcgoMDGEJRHIBUUwD2v5PDj
cQJ9W3VJai3DyIaOIcLhzGNFTbPhu3quG88o41wAnVGlhWzrXsYTtlpmbgvvbLDn592o+6Rx8QhI
x4sUuGkGdrh4CTTshTwS938PHyt/6CJB7gRLw6FF8KhvAIZowNNCEgBh5DJJ0khs8WmJAmnxY9tv
7ZOYb5HQVbmtd/nBGWbW4FfQ5ZfjQMobRmUbHacxPxbc1QbMQdhY0nhFmOg/MpAsaBuUbL3aapVd
T3YJ9OCCcwDcXlfBshuzKUyG4vKKa4fSAdnm/kSrrJj2mxvMbtD1QYMJaoY6GbpLFNlKlolzhn7B
UU2QoHlYUI0Q/mJNfpqVRu/QBbwRU9+9KvsU73NFYuLKp9Yn7BQpH48Mw4oo5jHn1P6EEZBAlR51
BfzbDvoRHxaxRq4OuydoIBBJ8K+/2BnNghi9N1mPpD+hAcWgqMaYtue08DDhfMeCWQuVGYxR/XCh
1Gz803+vzzCwQMiLf9OvqvKt4WHgKlkCzehLCEGXUKyfu3MY/0NzWAsD0/nKjiLpBBYM+f38gbgk
GjfrKYE3blIj0yWf4ytYtPDTm0GdlEYbqPDva0N2nvd604KVT3NnbXWnoKaEe+dwZs9kOk2eO1SP
/FJJsbaIcz7yJRaESfecxPna7ChF/3lMlKDQbZL9sQIxthmfVX+M95cxwSDzFLDmEyILYmku4c0W
Ko5G844JuuGWD5xc8mXeGyTKNU543Qwcp2QhdPqOreWo1VYbIoSxU94gyLWXbTPwyFTqOcHioVZr
xkGT2RJYi4+CBc/1MJfjju30OD5qQqispuvPdNKgZz4wpXyYr+v5dKEDQPaB13IebV6RQFNju+Tg
/V2V6pxSq4riG84SuCuAAe35zkTgS5nk3OwWpSJzOZhGyzW7lnZGp+iowecCNKEYDLSuRxDpu0dS
WWb4WT9VMU2JVZ6jN5+tO+qIvc6jEWG22h80NQqmuD9IlO+vYkm/f+NF177VAyFUw9Fr1J37tlWO
x3ZQybvPwpG/2oQ0NeUciTh2XAujceVlSXRUyq3LYLBFeSFZItO8/3vxeTf0LfhTxRBwFdseEG9Q
gzLRHFWzajyz3yl46H78zmQg1pLz83LTgMthjjqKyrvuoe2KcIjDa0SfGOp4+geIAiRBbdUSXJoE
UHtGps3URGKccTdfx4d8+2AkOT1ol3pkJH+R+fvhVlmyJHlomaiDpofPPf+S5hGEFqek9xq2x+cI
eWTFJoHjNNzqreDHOflBqEj/ggl1DMfjObatMcTeV+acMdg0P0q/77/H7EJYvxpskCl2tKGTMf1C
l/IKTFy3oEoODY9uEUcZS7QXCaholLTMJbJTmxb/CYUsRm/2UV1m/DzlyyPMBcmkvugr60tSvkMM
N7mNTZPiAfd7VMFI2IPoa7qeuEUp7KKu9Mp7iQwr+EM1lhfd1OlQ3UTIjSdqQOFUtKhQnYeqkj8/
isGFXaGOTglpKz1n8n37mGdTHMIGaUopHWHpZifDGEPvasR7MHn3G+t+F3iUF+aSuIhZK0abjIzn
GTINSAz+fVqlTVaqv85dmmQbyC15mNUmlUddqHRpiP0jJ4BUMzLEvhzNautRwCbRxwN3l9NT3ZMH
N0tRm2kaOrba5OZVATZy4mUYpyOV3uYL8i4MD/tn1zjrISoUpd4Ti3vSh/2bwfrfcnKlv1ZVwnO1
XEaZZ/CCrngfRPMrXGRZLINJXuyC1pYu+ODIMTXvqFIKQfgUdOC3xd8RRfZpFwRh+aSD/IfJufNK
tEPAr9uRe3d+BXH/WZBzK7g2HOdysFO4Fj3sB9jvmnbaA/QQIhjDmRMAm0rljqU2pST4d2A/f34f
DkZ1Puc6k0emVQiJbLD8B1AcwLoQMmmbFXOvfctqsFBa0eWESW0kXcCwzdd4yw7V1xwP1OrNP5uM
QpBd7Tpqzu0LnwwHZ24KsExtxjokOR33OaXdfJzIvUnTw+et8ycmM0TiNXCrpHw9Y9z1j2oHCCvf
aWpnuceST/4z2tGzb9uLX2yFezsrvtaMlk97/63eZAXBFbywspcnjLvbvSPcVX5ZR80L284AuSt0
lg8f+1mBSZO12xyLYha02YiSa6+QSjjGdxgCZdgabWEiF0KWqQU2RkPxDbxnHjOGIJvHQpLedbzj
eAZjFAj1L4ApARXSpZweout1eNls449xZKO7KlGLnJLv94nssp0hetTBjnS86omq6i8mG6cwoUcg
0p1PWSD7iv5ca7X3GKnONAzev3jj2xeRJkBn89VFtNkagIOH7L4MqBmCgSyE4/iFkKOtOtypUBMT
srVTR6oX1KHR566hWcup4BXyvJZyKk/gj3xTVNlLcBZCaxQapihGAUBD1P5YUye+tpaKR4uQjaIk
GeoW/A+VO8GZ3PN4+xSRvn58dAi4tZkObxnMo8HNnSXuo6UeIxuniNfUUCc9w6TrtTuz8mNfWalB
In2IweObSYRtwF6Zh+SP0H9rnYEsS3+5ipccBLjXQT7wCTjT6sIPcY5vqBCvxw/8LUNDY6iS1Cm3
7raEVXJ4lTQmqV6L88Ef5tcD0qE7aXJHbGNM21cgMB+Wt0t8KT2T9/+oZjjJp/Vz73zVyBXK9SKM
GdtjggkqSGP9OXNgnPLtQaZOgx9qvicAV4sEsciq5Iy0tm3li0enV6P0Q1UyZtPNx7NUC8RHvqVo
VnO/UOo9oyaw2p76KIUS2gXuFxEfzKX2oFezfYcXA4McTn7+EPcK+N3oJDPBR6ke3CbPnkCmgy1N
46BlQ0pxp5bI5eCsaKyQ3DNu1aTS9/MgUN1oNXyvYHre4Q61pEyl3c0rwpmlD/gz+oYRpNVEBZ0h
x2ACtGhdMjdLGBYPVAXSHoDIt+2SVTJa7vA9OWXOguu6i0Kj3bqG/jlcBrkbqrw+RtNdUNbmr4Uh
aUcP82IgRPvHyJkjEUMfJMNg+1CPwQ18vYJOOvWbZ/vgVAe2g2Fg1Jbgb9wYLe4WksNa9nxVdKSr
BocjssYLajpc0W8qOguNsU8XdmzuDVozwfIN8Os1C12UWetNcnQxJcEFni6kUvGFYdGsVwShRYdu
0ZYpVHLYX2D+mw78f8W47bxrLIou9x+hjmUjldUp1+ZXoqWX+6b/wLwLqATw2QTzw6f/ImFrgll8
V3J0k1sxAPawLso0nhLTn4e5hmOrFlPBqIcGV8OdaXEt+9etVf1H61zyEJEWdWCdN9609LjfKTTO
Zw1pRS9s6ygDaj0SHID0RxSTw78gJHtGvpJgFfK8FBynyyowXtlM62q9D8v/72qZ/5FwE82Sft8N
NcFNiQWRA/OF9JqKvP+RtvxPsd4/rN4++KCRa76MvR2RKo6UXYo+Z3Wajgqo7H9SiB8U0Ch8pWTZ
NSdK5unI6g9pPVwYKNF9d9zsla6EMBdB3nM8YMI6EM2tkjHGqCWIy9gZXvZ5ac4Nic0yp6xq3kQY
ukKgqb10bLZ2VmlYH1w4gJDA3k8EvSjjWkkjdtODIur0J6wzBpSJas3G37llVuoRFmVM3XFcC5+m
v+70TN+UnadPnrnSyrFLtmgn3HW1wGCZMYcQof5ZOWIkGGnZCJr0rIq6b54wrLVOTryyrNecRMtG
IvZxuPbSPHpkh0wj1IFGOsyoaxaMmLz8K5TmSBuCsqOQLVKCjgim6k/mr3TQXUzuf4ZqPR9dzAZb
RBWIPrSkg8npdBDIL4L6kms4sZRYYdEupPBTSMFbb43oBA/wUXZXbNGsFPlHiA9q+NDwrELnlABw
17rYxxLDtySV7HDHfammvPu2Mg/L1PyN7KmTOQVMB74T4EartcDsF5rzbavUuFMBLPEC8z7sL0dC
E5+6WNvn/ksE4KHfqjn49F6qW2EwkZmxZFuX0jg4bojNYoSNvTN21uVWR2nFrcTU3i9ii+uP0nw8
JNiJgQOAoIWu0RZtY22O28rPFCFpREiMpWZRebGxrk7V713L6zQmFTaOxr25uCK+BTuaacdsZomL
8J4O4sygkfRew+tNiyIlqj2b0ZCRyIObG4m89KKdjS/l4TfKjBPpq3T8w11CeojRw7/vmXcunhvP
culh5Cl8pDANOl2nUyf6vAklDZ2TcEiDBQ60DH/4oJCLNmncUG4GhpF80TDdyDehxzP5OAp2ZvIX
Gr1hauNzDciYuniKRAHtugk6YtU8xFBI2365yvsAmE47c9eX6+gCHgDcnsSlT3BwiQaCFCdnru0n
Q0u6oIw38W9koJ9F2bXLV1dC+mZmJRbUVHHWHldUhzBTOdM1WEJZlh/knVEx7vu+M8L0vajgnwCD
Yuq+8p3MlInj0C8XuGRJ9mlM/02rYbHXTBD0+Hus12wHXb+c3ZWwo4js8YJ8itG+1Th3tyS2nFo6
nZ6cIbHCCbgwMKx3rCoEhj6MtiFgOkYiT3mP4vZsLvoIFz0/0sj5W3BDg5Zls5e9HbgZosvZBQ7p
eNETtQTF1fiXBUN6L21CDotaEthd3eGMlBD1Yt0328l5/BajI8sQmtv03UaoOYbnIE94GGPyi07H
XBK6YslejGzURz6/O9UyUS7a9uM20usQtG16IZ0lkR3XwIMdcRjFXslpuVhXcartzM2eJcDL/d9v
QAgg1wA1fzn++hCU6fk2fUnsDJtVdHxi7OXbU7uZv0IwsTFlmupV/OY7qXRr2dHGX3gu5gTlY8Kc
qJgakLJEw+hrDo+rgpGDCPhZIgj5wfTM2x1UrusT0YP5kNbuY17wmGwxMQLUNTrDCcpwRPxCopEG
kCYAMnllvf0QdWN2yq/a/qubUokH3H3b1ZSPFrzu1NHiAcCOHbItQQgIRvm8fLkfKhMuGkF8yIox
8mlMbGNSP0Shfe+jYj6u0/lbkLjxajciIqa/VxLBJYujDAkafq6FHqdMpmEVY8TtTltCKMpWl3BE
B3x2DuLJMxmwkbQd9v2aqDDkzwSEe1aIgtkL5891OWgDKiUWrOJG0oqV41cDCvDBdxsFRPQ6U/Yt
Og3PPl4GJdRIfl6Cmn8mDRXUs5EMfW9oTq8SBNvd1wtG4c4zRwN9YlxDi0pWrib14PrRpBo6GOOo
lNd3C5eOuZlwJ/kp8uvWeUC6Ln3ZlbQBm3moCFTXgPGI9/4ULwP3Rpkk6bwO7k089RsILxhv0Y8W
15kqm7mfDItAvL+vfI7BTQvxzKmDz3VT8+1OwBACXNn7u0LNaOkQISOhZnOLWsk03+ULefpPZahV
WY3OlKEXI406g+YUgDoSM8zBF7P6ycLgC0RUmC54MQVpG58ze+mukDn5T2uAX/+aAqaVRs4wJ41L
eKWLTuLice8IBMhGIWX8qZ36Ig3AQof7Df02DmXKjmSTT2NilWpCj9K89j0Yrxtf5xgQIGJyCFVu
sV+nlodCFj30lpXSjlb5qYzcVVtet4zv+2cDXXSKGil0cXR2aEUDIogfSSoxQCGyqGou7GxmycCG
YZ2qVIBNLO9IeS58mVMIgNuroUx8Z9Mtu5RUzcUTT9RXiC5mvpX54IChKYmkbHkXICw+qvsW5w1O
IhWJ5TNj/qy58DFNnSc/c5RCQB9GXAuy7VKrs4Qs2dJwj6oRL5bQy4WjXjTZK73JxEdzXTCCTHxS
i5hPVYOV8c1AjEl23mai0cL11S1Wbz3947c0Cnb4N/0ULSCMAMlRkZ/eYyUqGsvb9vZbtq6JVfsf
MDHsUlkf7MijWhSGhVaaTfdQFb5gsBdl9uytTS7Muv2IuBkL23fXvMKXdno10XXYUxWi7/8dsf+g
zVlnN6UiDJkT/C5iaNIK9GhLE+avAOpkn2w5yY+u+ior66KTzeAL+OtIsRAuMPiiRMVu2kr+pi3Z
jfb3R0OoTB/8sZuNgm3Tiyt5EejKDlx+gNCR328guYFLV4ahJvSgvbQVR84y2s6hcrSUiS+1tpux
WDQNVhj8TaaHbN7gFEFM6g4ALTOYaW3avk736xG7hqdbZsk3eiLp2jFjJThekQKRvX4WtqX/mkuj
sYXV5fnL09O+nzik8GdIT13IYllmWDjpN0wmIo9zBsKBb4blSdcyUWcZ39O7gau6bN1cC06DiVE5
/+i+mXRR2E1zfSH9kuDhVUppjgpVC8X0Ze/gtDuqaaBTKrHA9obJBF/jnFdIuzZOY9Y3rkAs+Vhe
Lba8+M+nZ0l+lmNmGfQYpk4xNLNoAcUW3wj0Lgf86mjskNyJpLkEVsVBAGt7TsCdd4jSFQBoU23A
hkvzSl6YM/tf0bzRmWZ/0WDUWxHsNZKouWkWZHCSBbS+nP2NWtecVrjEHtdWYbVXtH51rdkEmhxu
nwmoJwazUwq7Nz/gQmJ/1U2WoqDeRScgd8CtkNWTnegfj2rHFOBqe+YbPyNh93dpsiRrWbRzH/R/
gyPwuhbfB3COB/fwZ64oE0nMFGHbXInXMdxhDld7x+SoFv+nucIOK3NfRRPmzjJOccpAx2HYjOcn
ozUglyaR3xV84sSFsLWvPTUKNIsK9gl7oV+WAqt8fPMXmreYjZrBTwaXdbLQAJOhhLQdsFSnhPBX
D/dsWx4KhlyVOtGY+QnhUBs1v4TmROvTrPBL2H7m0bVN9s0guS9evkiWO1Cocc0tYxIH8PyVsP+g
ysfpRT5xJf69X16njj86PznvYCzHA5Cbqevq8XymQ8UOI+YF9cbnzFWJiyYiI/Z+TO3UdrhrBdAc
5U3tzlu3XwD8SvbnWPY+3YZHedHx2D01qv3PBhAih02Rh086Jt+5/b1eeeBFEzhKcfNyWA5481Y+
oPQhqn/37Tw1nGHtHatk/ppqJAr8vQfxqnROqbK45DgPMaSbjf8O7ZeZwushKUaQiM07bBG2CIZH
j5Zx75SBYtVvgbSrZsXxzvVyLT2UOcZYqDyh0vLNsrNdMsYJU4QrNf2Eh6lXgA/afQKkGYEMTa5m
ZUBWZZAYI3U81w2DoWT8d5xhoZ5Hlgmm2D0bGBTEgHk1xg7SNmtLAnfEKjnlbpXCpzbTs0AE5/Ps
+aXEagpTAlogNFaaRFSUH+K/RDMmWpNVGST/GNQOnafWmc5ijVMj9GcaD6TU8oTvw3CnH9YpUh4y
isByo0s/hYLSf2/n+memxYKyT0zJyapWVJoiIjcWqGNKO5G7NmHwVB0z39HnA0dxqMON3lr0cSW1
CbrlSdBD2yJP06xiCgKF7Xl6UI5HPmAVULzvg9f+cCMW0Yuj0XoLTUHXqOUWgyBJG5BXYmIuiuvC
oiVTL6K1Lylhjnuys5CBWfVOV5iz0LEtvh6yVv9l1NWAoylxusGP/Jahasr/wXIXaxI9YM1AnWFY
KzAha5REyPjXx6kGe2C3BTuIOd5xXqXPukvfw10DkqNnxkHbPRq/n3aUOn72fiOFi5e3ygXV+t5h
N3XzUitlN80azPBQnAbfglnvADCJe9e6XfEUmx2MXQA7UJnHch+T0J/nHrwibh0U1dkunQpBxitD
wJt5gXoSMHjSBCKcK9EF5fPHsMiyFK+FL9ILr/aglSWgMHVv7RkSwcX9miWdUK7FtZhxosTD2Frs
X0mnZFGwR1lGo4BNszX4/tetfqq6GWnhUdewRORrxKDU3u6NN/97e+qBhrJzVkfXFml1TUjuawm3
aM/U+GMhAuvP2UbVefZnySd4bnw4aAh+jWzXco2s/oPnDkULFtSTBmNBv7uNCXKLX5UXI7Y1Du/Z
fh59kdGD+FxjKlWOT9UAJMbAI9Sv2luXaXOU2tCfqeMSgXzfvY6Wa1FpGFea0TcxD5aNv5FyboB0
gXI/z54ivD1FnAurnU1mbIZ+uNlAhLtbCufncHCCZFb7WFPHEbJRI1oJIc8wvH1ZxVSQmymUcNUu
GTLDklci05NhHu9ydfSd6adakD9uvCjyFOoY7WQ8YFxESG6BOTajqaoVi0NlZX9qDvUGJvJh/2Ke
e8jOCjnTyEVKUFvzjKUyWJD2F5YLDNNpARTQZFle7Bwlyt8dgDfPnBXkY790YZmBUrHzablYMiCx
orsKO0toe4ZrBRttjtugzwxJ2UtXyMODUjt68RFL/Ff5/LtiZWFBDmAVMKwKEvyIdJqtI9iDIrzN
scR4qERI1GCEPn9yYHQ4okFFuHYJVxqUfh5Tz+8SwekRoXy1nlanT4YFN9y0g7KpdHfu+31VTZVR
VWhoiWz27o22+x3BDpbw/ARvC23c5DySd6TdwljLSogHZ06UbJ84qXpE9RVf2QlFIKns9vI8id7W
+QaHxo03b9R5EQBecF0Nu0YPl4FJR4umZmGAGYMXZB90WN0joPLUfCdwLxNgeJPR4TATTupcdgAE
98T0OpbBQvXH0ldDwk50V8FRkNXtTTsemeY8tPH/u/YrocBDEqXgrSWZinqjbhhUb7RqZRmLu8Np
R04lDk4z+O/sK+xwrhm5g6Ovy5iW6OQ4f4B9NVqY4Oke960KpJ1F87MaL+/6vnbCDi2m4r1xZoiH
A3TBp6qy2buVPV2My16OrJ1thJp/U028wvvi2L0q+BkR9+moJJsJSYOZC1xEFC/PeHW/j2TmAo72
YP+b7na4PfysV6lcR4AleKXw7qXDYMamsbCFfPPtwzbZPeWiIQ5BC+Zv7iVeIeMGmjm7zQcx9A+/
5zBBs4bt6CUQjeSeZV3Lwg6+K5+KVT328HoBUJEwjkHrkDC5LdcDO+fI6RlBGqHqL/aCLDzjxpxK
Vu12I3SP72Nh9h0lPzrGfmZLm8j4INJFYXsgiB7vNksA8lE5ZP/XfUKly/sI/opp36B/FMGI0Jhv
yz/6/GATOcSnrzet18RtyPj8giBpZm600Hvz06oAre0OugA12FrXphS5OJtn8jlFyF5GaC1RCEG6
1dBAoH+0lFbZRZ/aOLqQCX5E9WOFyEFDVpHI2Kj8rz2/d9w5dWGhihuCf9YRZs1lCrQV4Ea0Edle
YmBBE5lwxq3VKepTp5zQmm8dfC5/ZJb3DmVNZk/ZLB7zWtIAKepoYTm3HXMIUvNPNNq0Y8ENCRVN
Mry641KVWk4UROf+cRzaE0pg9GbD1mgILjC7K+IOnIYVErubfNRnP2b50l06qPVBkTIbgD+0Wk2K
077oQ/SmdW4jyKMHgurCVi28AnUfi1A3ir4jTe76+3CEajGUhsFGAVdW2n003tgfar4mKUz/xuJp
nVVDmy/Rqem8n1j59fTzx1jcCrGVs3vYjs5tgYi0FbuHIek6pVWIGCwXgMJA7tapbTXnUQFIN3bx
pClP5UtKKfDDQ1v9Dr3NnwyNXrQqtct3osvG5vZd6LmvdFwgHnd8o3eaw7QGTkUtp4+1ghyFe95j
Di6ZJi6FsXFCQneUt6fNYY+S3y0UgRbfc1m8a5Xsuc9YqBu5nJfAeugDKzjjA8zvD17gERs5cXLh
LBSu1s4fNvimY+F8NSWmgxzPzEWS+gQfPw4ex8amukjs2LhmtULCnz6lj+iexRWz9vn8szz5hzhf
PVhqI1CFWCC46otYqDs/WUvX/iINYzMpo/K4OOW5sspnXQNl6RMlmtPM+p2SwOHAkLq7LspeOmF2
mHr3P9cF3iah4oneuLB/a+7xgGK2psOvTF/PqFKBZvohctODsIfGSi3I/nTo2DShfvwxxx5eIoxV
C9BJVlt4ErK+qByxkWUAjkpcwsXq9+mIVGxVmYskFW8EuWlhpndo8k5ie5aS/ofMRqoWpJk+hv+U
g/P8m0rhqSJAwGOmLz32/kVfsucQI92S7CJQWwFWp1TtIGCtAcd7THNGfoBp+xOLh/OTzoCv++8M
8twNdSmcBL4oytwsRI/Ddr0YZ3GCo1yXrUFK99lV2MXAppNA65b/pslpHJJ2rSnZjOYDq/mdhaj/
rAzkXy2hzftCjn2XVD48O+RTOHjurQhWUW9dtKz3aqZPag6rgIJtGKsR0h/HnVg5/rW32yn13TmU
22TTsRmI3ParazUkiDmM0Zb3x3RBdl/Ddv5T4RnQoAxg1k9CCswC3R/rvT4ueJ4A1lSaAh0qJFIF
61XL+wS11vRCZ4QgEnRtCApGum+gkMExxozPmwHhiaUMUJ0GiH+mHydjKS4ARLNnA3aDd4v0n44X
PZocoDpPHKAEcWLnslOoOt8HFEOJteulJ0XiT3OQBB8zMibWJKwFzTVdD1fH+dBssFKpH6O5juAp
rn5U6OwB9hSnKagWYmRw5gckgDh/hWomolIGlMGU+ta12AhWlENltIp/huZsrzdshWpFVTTa9s3A
IjbdHEGMlSrTOau1XpiKkTIC1N+cbDLbobxMbt/9ijh0BhgWH8xOvTPilGksXZglhIuZlhiHXDuq
I0zg7eknKQx1D6rgX6RdbBYu8yu9zpNkSISXemmD+JR9iYZ3wCC2wnRReyrFdxRQpBHyUKouEEdB
MeUpjIc973r0uxOJgXc71qtbAFFOoFwuv0garr/9po+/ixR8zuZmyKGezzwGe8bQHbDoRWBOYCI9
2APR9slUL/szwsUdEeUlCv4rAXdcApmjRBBOMHjOy018qKBoua56B8fSC+JRdCa6Eohj17oob0JN
yySor/nQpgXvxiciIejISLO5GcCC8GRYErF9uAmVkFFjoGbF23/Up9dimXIEC77rTOaqDApz4+Is
cz4u2HmHp4u9OT/QywiHLar6uPI4zCtHqocGnFlTyDqYq1XF5xpboXVv4exMpO+XWHd/Ys2wBTcJ
5xRwi3G4LnipizvNBNJk+6OLHRtEOdsXt6D22IkBg5NM2Q9Aw4jz/fJtvcKCEPjeS+d785Uc/3RZ
Bz9CT3iQACd8FXCpqkd+LAhcJ9J6eyXJq26BxWSO6CmEfmFgL0/XxLXflrg1lE26Ep/1ZUBkcXD+
MRMUJCf23wMqNW+R2sZr+OZpTPHycTJ5DjaVdFShwwOYwXUpSzSTSxeg5pBdo9Y0DizRmKwXK6t9
2v4f0E2FP8OXdxbjMNge5jrxxE7xlBehu3x1YuqBi7vgQETOqcImQQaLFHvuF4zwGAK4k3xy+psx
V9AlCTONAWpd1HrWx3cVCSzJ48Fd7efl69sbqXDzwgQmVWGUBPbRZJZUMp5UZbo2k1h9/9mY+CHQ
UzcJOspyLsOWmQG4HflFIKbVUmLV8Z+U+Xw1KSAfBxpgupkCjfnONZNhBrspNvzo1PveQ/FEekAO
Jyf/Xo71P/X4bUr/FVESTIoftvGCMRJCXAaWEdK1qZAONUcQQTqcvRZMiQVWRaS5o4RRpOiYXSpc
5FAwwvrubxiAbIty4Se8eFXvKl8xZ9/MNzGMSuZk5Lm7NoHb0v9kCG9Ks/QwOeM5Br5ui1RJI1Vd
mGM9hZBbP2zIjRayxkqHmOZizVGiHg4fcEwcR/iRROWbL1BKFADycm2MaiNYXdGXaMkr5Pz7vPqY
W81QdhJtqNtjdTsdR2L88uKk2qKvehkkq2iMcv/1vO8BAXMtXS5wjaoFv64EOFZJQ9hYoOabCAat
LhLYoMoTytFkwEno/F7qKSmSLg3cd99kk/VDPQTExmrbPaJEV8CPwpPWopkiIiiv9JuRPjbluFva
6HSgLcoV3aEGHQP66fBPOTOtLTjpZQZHFLBjuNo1ku5lYmfItXYslmDLYtphxW6l/4Cfasr+VHtt
+BvvqWCemREX5uI26NPnB96CmtNoJuSqwLd3X1X5ua9rQAoF+usbWs+AJJm67hJNqfCJCPHoiCtX
LGK/d7xZLvYGj4iV+FiEfx+k0vaJE8N/m7QeC5yHtT7b07E0ik9VLszw4bEwZEQ8dR+JTf0zltMs
6PfPVsM/CJtVngejgRn9ii38FiWRoVJQsJEYS9rycQn17VY+WqsUDAtck/kBvG3A2N07bgZ7e6Au
s1XBNoxpRtRhxriPeuPwxnNsETJgQYTQywPMu6TV3A07UcvaGJ0qMrt9Byz9uxfusrnZg0cDPZXL
zd1kyifPfdrnL2OdeYH/n+K0SE+qu2ShnXCqf2mTRM3xcg8OP+OuS0lNta96qq4yf0bbzttM9jM7
tMjTyDe26XV+08EHWfpytOKn4+XDm89c4wc08EP1gchNHku1oUlyMta/LS8gs6hEZj59Bu2ioXbF
rbpa7BeAz5rQjIVRlAPPbhzeJRwjIt6/DnBRv1wU38qQ0ER1g6IvaFHyMUK8wclWnlonSnPwy9ag
sHZf3l2bN8rFUNiycOInoxCaLp/8RnlxP/4rrKsZJrMzDJLV91b8EaKcT2IEXaoLqvG36oY0dAEx
zy7SYFnLrw+mdj7ac7dwcsVfFAG1EfzF07Tdu2topWUKaC8ocQTeEsKsaRigX48x4g5AK2sZQgcA
7rNCnZPqu+EphzYC8jqCtr+BefQ5uK5eagkfAme6Mxu3Prni4FVxcJGEEHw0QNB7b++j+Ud9Q9ln
2eCjj9YfXk0O/JIMNhbbx/LZkKaQ1Twz8fNPaIqz2tRjDfPi1/5koXuO+e/+Spw1l9xPBzwkGDH+
NQfVmfgJZb6vy0RYWYwQiMPVphLAfhluJnTDNYm6Rw9YHu28qTz7ZueVO6zkXoWu4cUoApmDURgs
sLRSeCRZDsRfbdudUa0WziO0agX+98dZvWcCcVcTMokp5Y8fFXS1lmT16jvqWaoAzH25qx6D0ip0
1ouNWF7PEKisIbmkAdaBJAljkFTN14/JWnV0hkNV1zN47zfI+h9KMFMSZ+e+zet0lEqWhxBP/ftu
pnArC02WOzHahDrKwJ1y4mPzOfqUNfmcR93IPRsu/WPDcHDLolsU9B/2AK2yWI02DUOVqCFxItd9
xLd9J4Uf+8Nm8uzTlrOVtb4oQAlpXhXrx3EfZ7yzd7lrl4hKrgS34lTCTp8IjfL6kfhwbrvD0EkB
f5703VhvID3sFmd+NdmKGzfKDZ+DC4UBy32TgTfVlVhuWUr9vtqh96doZIRIdUNENnfWpFY+qrmH
FQvtxroNCyTFoIXRlhoiEKhgJSHbDhbOXdmzGSYAJPU9TrHJrK0SVsmdnwDNYzyiDlNH/veDFfbT
ABuLwgf/13Cltzd/6n/d4guL/dPVrJG6wtp2xrZh+EBJnqKKsLRRZzgfjl16Q1sUgvvTpoKEFv31
COtQcO2EydODZFfBHNkiHFmFOop6BU3v3lAuZ+UYIFVZc54H2eG7EqyhUIo+/x6EZrBB/GOrnriv
u6av/G00uQODoP04HEfu2D/a3T2/hryAz54Mv4qdV1Y/iMxjAAp0a5HTYjaLUHo9nsAPnEIHNH8w
Hiym34h2UbB3sBplMMXmc0Hqe8/8HJ7CY/04DgSP5FyxYxXuI+470IvgCyDR3S3ipr1RywRW23bM
61mUtfNYP/Y9OrYnkfD9fzRhgXPNdV+ApXH7S5/6m/RDoqTrFNlrf6PtGzliijnG+3BWTT7Al32L
dm4Ss3yj9J4cfgiDP8ZCYQDjOTCPXdBVS/lJ2hsL+rXYKANVqrnJK3PCrb0vAfJZRUTWzzQzf1O7
VbOaeddahsdGQPJYdoV2n4upDU9JcX2zzm1+hSKdN0IF3No821V2V2h+/Who6oVYzYOtMDArG1Nz
5BrQwmYxv2TP7nrQu6SVx/eoVyfrspLdPAyydLn3yT4iMTWqnrVszdgKW1vZ7zgy0+im0KSaqEpZ
2n3YB5KsOsgdrtGZrHf+uJXl6/+S++l9gHGQyyzC8JpjpF4pDs7Nd87wAwdzLHu6ThhxkP17HxzY
fJKfrWfG1f+FEzuJolc+6MRTP9zQNeiaLsmuNshzdiQtY+3XkFplmgNm70m/uo0V3bJ4Yqhz05mQ
nGkps3MZpC5tZL2uLdfpvgX+TDod9BLgkgP6S6C0GxQlTZKcSiPL6L5k3KIhHCQT99aWxMkZr1Aq
k/srmOhugO2rzyAnnLhiyS49LW1fmggHDXwXwQzph6bgfxg3zWcbKAlCwS6TCOUFJG+GuO8jyATV
d73xqrZZSIFuvWnGuhWUe1QmMhFAffQzZTOt9icWFJkPZ6WBdmbpHJgHdRUnmyzykXbx3tM041kN
5H82LKRj8dOrdJtDXjVCvmByKPwFQxV659HBjQTauVWOQKFf9kvE8gT+dB0IMOsv69EigfOm9kAo
H45ICzr5IqmlFMsyc3GXBMXlDOF7F6SE3OD4DJ4bwA9SY9FT/yP0sweE0piyqhSosJu/bVXyMqAq
g/FtCk1FURuvF/N9vnXLREnQH6pA2uLMEKYo2Wgy+4owU329F2UaFyPuLpQ8pMAV/GHYp3HzNi3A
fepccI6XyEHp3hL1UVTu+b/f1R9VYbGoY839JRR5XHRMD7B/wt1e/0Bixxy+vpt5yr043ZeKkEAL
9b3eEFGPKN8zSXDPYkGgwOidG0AkXUAcDim2eoDuphj8MX4Pp4EtJHZgOwoDD+xPcaUEMN1eiYju
xYakibtxtoT0uMWcf6+aC0t0s3CNq8Ba5QIi1yUQynLwtarpNZJaomZ+TxKpw8l4BSzkoBqoFbQH
+poTstEr95wGyarpifTA2p1CbZAMTepEmEp7C7y+1VPgURJzvTtaz4uaf4EKqzITnnPc5byzp6ql
6OWrYjiWs/1xN1aGY1uAW318XUzb2KK2ns05uz7ojGp3Pm77x7fb25db+t+zlChfkzJ4TI4FmoAy
pIVzgw0Hb2nJkZ8z6BGfG4YikjfVz4MUOeOJgH7ce5xv9WGz5w89Y6daZhtK/rRt4Qxco+N5qlCk
udoEFYqDzjK4f7HxbsY/YeCJIO6y5l59LpAoVBR71+pE701po6j8ruWJAxgBQ9DuXqPToNjCuELe
xOj5MRa7SCeK3R/FLpv61j2ltBBoqecuPWnykJxxqPqjWOb3KZ1HGU+hwKzsNzEmoGgQoo4323re
ConHmJFpS0XVxoMA6Km678gFOdVcaHmbhUcAyFFkTGwh+5uq/7+fd0tt2xLllFuy4bZAPXAXFwAW
tflL8Ur7fg6rQB/CMGSQVy7f9kz7ktrvkW1gG5+0dfFt3SgJhx+ibQ8pv8SVdaEk3WrEgRxSFrJp
ApLTh3X7bLM1O49pXJ12C+kILTI3mmWXdgJv2+bC6igS5Evmzerg2FQrUm9J74MM/lt98Cjx+PU1
d8sz78eFxJ7ox2Vg2i8GrPSn8DhcnNtLER2A0JIljHs2dUI8ikRZ6Pyhf7iTIYH+I04UVfz8XOrx
7oS45uyB3rQx1l2MHrC6E4iat1mG9bL0jTGqNeDbApxR40Ap2/exe7RsNL19jrFnK/DI3hq8zOnw
x9H8twnSrVedDWWCxOnRKTjnatctpTyGutFzghqut4okUIs+mB1xMc23v9KfVGQN18+d3cU99gD7
KsbFwMVcpVnG2Igojq+OQVaYauVXHjQBPNLGetKSQZwu438NZsbtlo4NKTzNBZ/GluxhNYmiUBVF
AJ+vQkBKkSwqKfNee6OMLNwY/5XwSZGyk3pLXKQStSSUKWPAxOAUjrQvQeF6cYHJq5sSMTU5f4HV
3vSHQLs6rXqBtbfdyUiqBWwFXPj6aRqyyShj8vZsPsQK6E2PpeQ+ihWeno5zuFICncykrAdWe6Cp
2x62q3totGx8fzqI1SK2OA6Efa3O+t37Cz6G6m+3jTjQfpZI4x4+ydIJ8RuPfX2Ox+wUl6Dp3imz
AQVYmCxWFHhTuE6aYpDOXSfFYJ+YN4zZFLMvL60luAK14dV4LQ2NrVmEOSnnUzA9Nw2SQIQDljrR
4tOSwoGE3XuDffY9I0Ud+jxanfbRbA5lDZ9JMY/Kib3HL1on5BWti5JYNH681FySRBlqtskbFqzt
E0lkK+3xKhowKgdJGZdNLUh5lq84BTkQ+r8pXf/8KO2gTLVVGc2G+Z6q7KN23dePjwoB+rok25wJ
Ceq7z3yJd3ZnsuDfkrwuJSF3qvsB3U2t/anvwmxigXi+zP28qEE7yk5eklouMjtKlcndxQTkAGlv
I/GmrjYB6ZhDreJR+P/78Ko5kLfLnmGUPNI0L8iwpMIsMqkSHPHrZ379xGEkAY0DWaUbP+rpBvAr
kQf92Nlcc9uowAbjy/UfXZFIxB6PlJVPsTF0kyiNzg44ZJFS/7OSZMRJ0VYc6+QODLAw+9alLVAm
Hc3ILAv98R6W+1ZZUSQOc/HZEmHTE/Nr8QNtQF0/DjzSYfw5h3C+MEcPg5bdYCV37o+SavRMlNU4
e2P3QYcz+J/47Sy8BS34rsafviBby0CngRwWc4htl23Y1kA9sOPdm1kRHDyi1nl44Xeut/ltSDcE
YcdCWsRsuK6YsjqkiKixowlMxWL9K7XfW4PkmAV9DB9sN+0BioKskosDzIt/fzgLb5tbdUgw52qv
IcNkg7MgMTFrJn5TNgUJPq7IMjJ1b79vn5oHwIvNhta0rJgZYh7XZoBn0DlYnAmPMQ1FlR1bFXcd
YULYuvyEEj0JnuGooIDuLdlmNR9vaiHfkW3oBT+q1DBUSZIbTPwUp7W8RtAn3E68ZbrXrE6a/zJc
3CtH6cuwCzHslyUb2GFfDVcoUmBj1YyrVWR89l4WQG9+vmUsvWS2Xboh5Ec66bLibTB/j0jPDNE9
8ippIiMyo6Ay4HyLCUf2mQh1s0Hr1ROoDtAk832XmMqwXYPVWiu6wieAU1fj1YUWdsPOHnIfhYyB
PnCGT32/ylzTwTDrSMSbfxF7YuV1OCT8P80tN03adS/eoZIDaIvi2jsCymezcz0UnvQilRWqw7kv
nTHkzQAIUmX2qz5fDofn9ZHfdjJLUug5w7SB1M2ETh6ZpiT3wJc6Xe1dNGXLmPkdvhqOyU+rlKl+
As7Vo0gAtwbo2yoc8PJ7ndTs+EYhYw4lo+cipiIGvIaBrMzFWyoN8+TXrq7ib5rpyPkcmizVNuTe
XJDiOqw/DsEArfQOyzAKdlT7Lg6s+trfVXZjh6EIFUciaOcSQSnJEWNUEMmpxiGY4OVVzhNBBPXK
3DRjNiq5kTeqFUP0JMVaJCXAWKrJFTur9o3hNWzayugjB2YO0ZZk3zIN+l4RrjHQ9S7+opLPmc+q
yjuv3Prjq5QGtHhVrctROqTqEmoZGMVtHvfS4bTXQoPE86aQmR0ejtPqqj5j6v4tLpRdxmBFKNC8
n0WJnfasSsUoI0HwFvxI4H8o97JYgzs3VycvrBZRUmfgUwrU2b1GM+GYwJVjPvejIbinxplOo3p1
2xTgN+TAXF/0dmwxlQfDCXz2F3Jp539wJ31w/TkMW5d+q8fFyHH6TK7PUAwhEVojJ3S28RpWIwaW
eroo7HFyCz5TxpQg0c+8m5AAhyZgaqofqvY+RSuvqJbM9WKVE+DEfEXb4LWK03jOO163orcaK9Qj
JN8z5UyP799kY3Gd7cndm9sFMtb+0MXCpfIiuUgLah/b6mTDfl0oyUK/C/mbHyzdvwcdOrcMFZ/1
QI5XwbyNJAc++tVzrJ6p0Vajix9vzJcr/7LLdwIplH/uoHryXrXGfTUaNWK2BE5w1iPvg3WYOXG3
YQWBvWvOJbH6XqiW20swy4/EZZUxrNZEo217SL83nvDo47ji9Ws8MX20eiJeU0YsmsENrXVBTYgs
+/jPKlbq/pr+LNAoOuPl+7JGNaYFqmuQQ3n6tjWFBNj3SrktOMFH/xWhBCKg/KA1Cnuv/RHruCAV
5Q8ekrhKDf18bl5SnZDMZN3ywGJ+cnxrJ6AJocfhwHo9VJhSWeTx88SIFCcgWY9/mXWys26EhWPR
JglOcuHWVY2Hv6REVtCmcledvPNLTHD4egfZwoodjYU/qJsebVL+OxLt2xo9Z0XZjmjXiyHTlTz8
M8U8R1chRHaSCT9Xomn8HE0QgVoDPvF3ykpJOhn+UeFob+q55ZVaWrpbRPvtEiuCdoqn1DZ9QQ8I
7vwUYRSu+BVGIXBNnK/nYrs5O/GOyBhrLMtG1KFoFlgkcHqO/SWUdp0XfI4oY+EwBLwuIHKldykz
kUkVt8/Un7/mfX5Yf7GlAG6x0MQgEblw4cLJAQdTsgZ9GIyFd2y5C7SXYagXPEv5f2b9szS/9D7G
ahil+vaw25KpoBlkmTmJLZNL9dhw2noHLp9iE259eZeczgo7oGVk9SoMf8uhAaOkENkUUw1T2EwV
AZKkmK6l2cxts4Bf9pTCqitX8ELxTGwkuc8uQmjHoAYBbh+WGmZCq4m7e87Iam3OrANFIpTffvre
y7a69J5wR9fBqJL6CR/CrEf/GVF34XIgNN3MZhWgC7agFxp3VjWBwsKX8+3toJwux5K2BPzqB5zx
XiCkF4sjjDVXBFlJh38DAdN9kZiE8yvHpWeBoac+7cvgbgoWYf+e6njzv6F62wKd154T3H/Q+4HB
vkCNqt33NJYcfiLqdMcJdGwV0cD1jLdslGKBNaFKv+TL1uzSBXyYqXEPuuckTeKjoQkjblwNgZ2t
ZKzKSLQX3NeyH0THYdwoKKIFQ/bIVQd1foyYnqf3l2cMqV4tKWozojrsHczgLosnQaNG5R1G9PlH
rruwIrYTpvx9ckVYG7T4harUU6ZGN++sAW03K8Ki7m19i7tRYq+45fVvuxF+Y6c0aksQ0u4T1GcX
Ele130bonfaCPaecAcU/ahly1j9qG3ediTlJxodTUDnmPcTgyoZf/7BJ4Nt7PyFnE0yHMa6w8LmZ
tUzNL94n4/H8tfOri9bFNyoJG2vFxp5lTAYks/JUaYAoxPGVLdUJXnWpozqHnyZqFmJ6A/1bP6eM
YwOiD/LFYkmXsS2Slocbfq9itp92IF0n/WF/c6JYrglx5mqiB8FCU7OezhUzIkSxCtdaHeka9DNU
36i8/0/b3csRqoii77Yl0gF9fNo0+ygQxyWiwdYLhehT6X/EThWeM4vWOtGNKHHikWCJULtxiMB4
Ux7sWj5egP0AQM1MszWhaWYMK0GpjcxfiZgFSC5bvG47Kt7soeNgLJcP/SmcN5ruVm/cOL/P1hXJ
t9oXeOkcqD9W/6+vnE1BTMR9g+j/pNdLx0LxIlQiluyqUar9TvlgWNPgkuhOJDGEON0SB0JCBkE9
9zMZuvGS7i7AOtD1Phl5MmckAbodkB+g4Ypv9j7FRiOayK/2OLqn0zt2ICMBqqpnFDJdvXfVCkwp
b6Cc8KNNXnTrScWRcMcLaxtwDlD2Bc9s5zQNy6QDimRmZBhs3g3ljAaTAAIT6+VMklaaXYXbuf4c
m1ZA23UA9BicASQs/3/6e6F7BXerbNdgl99tjW7m8ZnG6mqxOgPdCRg6YHt/kIkdm4mSrK8wYt1g
vRzfWawRWlUURb0FqQ/2gVeXLqmPnqY7Ono+IXCooinTtVjsXpmHbEMld3e0C9dHOd6d3FOLzHbO
fOVrSGaX41hMFtd7cNC5BBTciPdYiuXkASBviaqN2cffwhb+YaZ+Ovk3g3EmYrF9ZMnfhc4tykI1
jcOIDeZyU0NWc0GFss2tmxvgdw8iKSs1fVoGbJnKC0NelRVudm6ofuPI52ibuVFDb7e3TaMM6vua
i9nbu0FSA+YzWp7aBJxCKgFEQtw9za/zGr/El1tX61/ZXk07QXfweFKhHI5NKZ+xQDMLMFqGA+It
gOqP0of3I8Iur3hIgeMV+KwzfRTvM7q0t+MGGUQcMw2MY4n5NX1SvrFbblhHKPdBA89yEyR+dTQ3
f59L2w08scPWhC2Ocsotq1QiP4wfs212+D0i4ta68ykcyyIBwv6IyjVljemQHFMoTHY27RTbF7Q+
WQ43vyrbSlLnV4bdn6aRNW+DAdZmI0fUaGHblZ5wGOoPFgPBofM8hrfto5vMLaKADnPs/NQqcpei
O/ikokO6anSNhQ81KhymAOs3bABAz3UOsnfJrUfB9GRT4eavkjSi9zxIXt6swnkOxZl+zIaOkMMN
XT1GhIJlZa8Dyxieu6Lp0/Xt3LxV0uCOVdmSjzw+K96ZYu+hiVI1Sn8gQUcWCOvu/9TnI4g57GIT
h09o91Vjhs90sXhSeIly3KCy+hKnerEIFDc4lZfuO2A9QhBwM3VMS5p4euAxExtOfpTm+6kPYETU
IV624GtpefBXDYjLt3/0Slqrx3Hi4sMFjbYDv8KR9QlKgHq7EUnp5yJ8RhynbTZNfLLzsdOry+JS
N4eSKuEw6reBYPG5oIKQbKmxWw3SFqEKWpOrgDr0LAKn7VAT7tOmcwT7r6lEXNaOavXN4Eih1/XM
gwpCxTMjiu8+ZFVW4IrwdyYFJPB2cvK5bNTc4jk2i+Y71jYpLsfWtYoGA70AAxCLgk5PTugXOwyp
ID2guHNRuYKIj8ifYChjsRwfrW2ijIPvru+0/XLrT8QDRddVC2pVtQGR/m/pI6GEFoidW8/J/vzq
j+exbXLQtLN58+AIPzo4AU8ZCt8NIRTJWHIScF7+wJfFs3l4lrnbOOpsnaHs11BpcYbTTkFGkKe6
wEySkdoQhcksLtmIRwdSHaX7U03tZUZK+90v8/a3OMCgQYa8nxQLDMVLVLQPJdm1a2OPF7B47DT8
Hs9Ns6irR/fgZSOE7WseZ6KCW2Z/tE1ZflrNvjpZqTf6TMUb0jDEMVDnAUpC5OOY+g+VAseNt/N+
RUzBV7Ott7leU/VcZlbQdr/mTnzNVYAwxHw7/zsO5TLx7vkmYIKpTs7EKU1ZQpLd6bllplFS6uLO
9o+7bU/3d7v9xtHo0nkvjewsKnE01L/WNQJpPjVG+VawdFCeq1HRnbBOqkqr8P6vqZg7wKrUOryx
n2DnxySCy4QJbSciueeRA9NdBDUU4+zfRy/BrkfJZG6QcybWWw7MSAkNpsZKf+NldYAnnRXPOpQB
HZ0QZyTJKrm+QfkkNyR81F9hCYNqwHcjpSNxUZBcTy4xqBXDz5jPE8chP+gCsjijUXygVuMdTnSm
MWGLJWZIeT6zzPCDf3GW2KpS6l4m5iM+W24+BZH/ogxi8zJ41Pz4RmM6eC/26qWgCUI84iL8PGps
rb+AE/OTOzIwVH+rSNsH5cT9XZ1kPfYOkkm6M++Lc9/OvxaFrjPtIXf6nkV7AKfOQU/5wFtn+ikP
t70Mv/i/AXlaKqihH6LALDBSCwQCmjZ30pqf8DPEEYJGUWVSCeze8Q3w86jrhZsR2j1YXfNMMIxT
gok1gJsx4kA9hwdJB48RrqpIrnEpVuLlLuphL4ZA5yAlej8I5ZYUUDWLDhG1/7SJR8ltqRl/bBwo
wwDtTsgfAkgls7az1uKLY/9UQCJeXhNlf2pE1mb/ZgDxFcpSNKWgBMV8AwptLE8A7bdYOE04QfMv
c73MyViZpAWz+yJR8I0p7JMju/gc5N1mGxa631Exxrzp6NeNz2U3x7m1mGxke2z66KG63zaHMiUd
M73zOFnck9mupFUDi9qQXDmQdM9Qet0wdE1WfIBeayruyUpEzC77EgBLzu3RZnRoTJYH12Muu9FR
KBNAioo7fm27CBNwZw7Cw/QI4yL/jsNWaW61d/Lm1a6IaCpGvObOrrIdmJp2tP1Q/oKznh+u7m//
wePDMlyYWljFUGyLeaj6OwjzFuujOJB92BnRcDegfIEm3bXDPBcRkjqwVgV3TnuDTVcaoWjwL39F
he3hlgs4G7/FGM74A+xp5TGl+4UxBFkGhR8kL9rHig3eu3/AHw+j2Pel5hy7lG7W/WwsxEIYapR8
hk7he1WRsnAFztVrpAA1wSL9zjKqk6ZkjAQrL64pRs1XYjbJ14DtSIY3IOZN7mqAT9oafspbVtYV
IihbIXdbwVcEWIL0GQP6aFyUH0i0bkpjQG1B1XejIebgAEGTSV+Xz8agUq1FwZlOMj1aBkKrNLQZ
9cSr8v02+pt3QK00eShFzLshQxnl5asnn81oPUE2U/p37/QRwIQIt6/vlYN0pXWL3SNPqZzhgS1X
t7u0VCDErLTxdjyK3NHo5lcOaheM44BsOm/7FaBqB8Xvy7xiunCXXGPFgO9engdnAXBOeDk5WGgj
ZEK40JdvDJy56f1Mjw/oCgw4bIoHX4OQ121hj7ASxbZ1QbnsPuKVRUnAomyu+QO227O97SopwOXG
egEARtdeL0XHoyBPlVtBJ8l4yxEMQSN2g9a9wJ9fUHkiNcEwWbJVndFaoMqSX4xyLEUWfIFvSFFB
+y34fz/v+14PL0XuyOFdIWmCfmSGG9EROAWec42d54Yw+D+4Yyab/I7Nq2MKqJfkBWn5uOAioXA3
TXv53JmEZmMHktYQ7HUzgbZ1xE7D4jo7783vX6Hfa36Zr1kdowtas535cgkm2RRVC+tjk/MeejPl
kBp8DAB57q4zsKa+NDAHnzMGpMYfmBviSfQaR5K0VVdMqEaz8Vk+T1R3+8bmqJ1q3SQSmNXea9VR
YWX5HV18E6wkMg1He+XV0jHcEcrw9s9Fom0MZ99iDUp10xKCaOh2A/Sg8ALZpK3q0eso2lHaCbLa
i+FD8MRoEEeac5nwObGQWe0TqfRleFRZV0q9YoV0F09c9iy4ZKVMzuMDPebGUYJsWS4wG0toLE18
cAL0i2PoeTe4Du1rmtKK/KSmbenf70FWlWNJdad0eJhWSqhi0xi/jnMcGpZeN4VGNLMu7Yd7aSY6
fdXu0iRqLnuFiCFh3s3JNL6Rn+Pn6gkp4h1dVLBsjoL8wsRjtV7WgdPGc+ekYfISYux3czoOkMga
8Xs6K3e/oMbToqsz8QMNtPy6wJVm0PVeSvVXB+Lrg1E+pgOazktTozcnFK4MfL6ZvCD/R/OUx9UO
X4vgFciYnLN36IYPkAnFAOPnFW2pJYiRtBlAXv3tr58GO7BhPNj5fZcQID0f3zoauRuECjodKS9+
WNQFOpycT4/hPqsl+XRVNDWe0v9BNQXvgu5V121C1gYBYELf/ju+WuDjQkt/8vMdlYroStSsQrQm
pxtCkczwqokZjSKWLRGnm4JIUSToiQvo5Bz4YPAgfiQF8dWKs26bXTFXGXmYyXvHY/T67jq+6Mib
kIvLw2jkZMyEH97kWwhSk6dx45fBGHunexRhm3jcuWnAUdPV7U3Ri09CYp3L7PPVwyvJp1anMnKA
4BiQR2ZqXlYtQorGqbQdah2hzZzq1R/0+gq+oMIJUgWS9IXp/cITybyq0qfN9sFOB5iBahIsl7cl
H8rSV4NWaRBJSXoWr8dRDmlmtSpCHZU1ZQ9gdzijiOTTw8nACeVANFRZ/0Gs1weIv1+/YJNoqMhH
F9WV1kgAh/bDGr3dl7rIRT9v8w4jyF1ERmb3Ddqh+3RbyY17T17uTYolGq05P5ApAVAOul0WLVWL
5zV9Knj1eQBC3tQ+zBkYSTuL95fRkh+KA4heE7roOtHzRxheMKFGl3v7hORJcPJ2Me5TKUkXnbVB
SrYldGxeBnvyRACdxRjZo5hGvLYRaVhIp1P7+A+P4zHtGvLP8qKhcRt9ZjxcQ1208eM8qVGAk7uV
O4OpPw8AfAfQsdnzv1wxOq445s5QzrQdWw5t6364hqADCzOfFSmiECCAajgqUNoLh7fTzhM7oPsj
QyLsRdHBeKQEpVRzGW3eWeAfMeEzpMS6/zHjR1Rm0QkAf0qJFYvuMyy3qgd4tK1x68QwN3yFN1Gj
OhT+axjouKf5RK5KDIz0Eti+K3P+XUPv8SKIqOAf7AvzALkkreQX41K7RX0nLMtyRpBqF/rOPiDq
9sutRuAkbI9Qr38rcVKm2sgUIYHeG0gEIjpzFbdhkRRg7o3RFj6QQl5+LmRZcHNmS1YTMl2Yk4jh
CS1vyeXb/9XNgqQFOLoKKTL+uRjaUtLC9wrvCl56W/yR8YmBqFIXXPZ9ZQXaXfEUysUEXYAG6vCM
wJg4yLpR4YCPXKVGolBgKd7DXmi6TxY5Id+ru3uOSWyVP2V04fHoksrYOT6xdB+BGzo6F+nmfk34
GlWJdEp74bsdm6W/CU7a+10UCgPxDGGKHwk1X422vcfXycwlj8fHfeb9oDEdaozQfO5/mVydJv+q
KIV+FG2BAidl5k0bsC2B9vio44g6A/WgQpPLFgfSin8sF+YPQIbrMv4SKflMRBrav0il+Fcvkz3q
ZtzG6kItWEttg2K1C7a1EN0gcgrgHwDtiR8vYN7jAarjhV58mZMrgPhw5rZGqQ1GksFft1QJI5+S
Kbz8OMOIDFZiWFuExwT9gMtdECxu9aiVr0r2hpgs/bfZuLncEwqeCXDJSSGyiXUuyn7FgLHbV5Vu
08SXC54cQPG66EqOyn+YRshE/zrgvIwvZDuXqVadMeWTymW9EVewyYhtpdQqtmthw8iJ7XS7bew2
gagl/0CH0XnAW2YErTGsUVNNOJe9hekpu35soilOJN/NSq+UWKIqxLZ/Ifkq7ELyRHowq/lxYZJo
Qx5h5kJ2JuzOlXE4VD4D4waQcNeIaz5TGf0nGPL/Ba0rN/GKylhpKD/BWsU+yL34sDU7yTgoY12p
iU2Y/49q8le9wew2fl8QD+l7DeN6G54XS546H2if1CRn0aUcCA6gGY6vJc70T9YpSu15Z0f0H6Nt
i8zj2+vC6FkdMBqSjDMGL9tSSXzH8lUfO6xYP8UzmSV+G2s+EL3jR6NkrD62P6GnwqoMuNWTQJv8
ll4JfE1Vhs/oVywWRgCsRahI5hdhb2IbHT69DMhy8aUksYbDiiZl6irP4k4+potwSmCg9iJAPfPQ
BhlR8cRG9J1CNMc7+Ep0DG3qZTUgatK0Eu1DbKwiR9Uj5DEhcGj3CvhOpRzBEmIX2R5Oj7iJH9iV
aBzyFdKOEQGcXhcrfCQJ5Dv33QB0V2M+jyKipuQfaCppxEUx7ekM+0Pts4TKTtnw8vipcMh9UIUK
rl5O8VjvOIBHDYex83C9guqncEpgIaJ/Rw49/MiEwFnwkL0rvRBydhJZ/k/wmucSL0bYVj4jFz59
9ov0Lg99BqAr7QUKto7CEIEl6XyaGfoW/rF/R+2oDyv70zkl0RBEXoLNTFofKqD9Ww8EBHR2SB70
vB076PU0dPLRNvchLlgXsueP2wp212dy4br24S01f+wNeHVTticMamWvT8jIXaIalmBC5DX27lHV
i/u8LlsUFWVDaOZ5FxKhc1jmDEa4acTH145dMsLg+glYpptWt00HGzwvYhQFLvKVi3ulssn9Nx2S
pDb4cGNCrBvYRVNN+iad5R2I/dxTKMpqIEkMfdkDPAayjNmPlPXmPpEJvzj5kwWh8CakgOnrfVXq
VpLGCXCc4UhzJ+F2syb56qJhO1FGBvHNlRw/phdhQn23TkjQr4lQeNDMxB8sZ8yfZ7HLULboM4bb
YY2X3smmolmiQpAnmH/l98JMfvE+Mj9kdr0t0hVZ4mTaLPNVzPtxdOyPR/krHTvdHolRtwjpaS3O
I4wf4E0D0YPkm9yLVd12mltKvUdRihZVLJDZ03mTmEMQHo+Q9eDw4PC/umD5umg3H0Kq6TGGJG6j
HgbXxSBPq8uNxQnk8uPUGRhgo/4SwTMYzbDPhtIQlzKX5NYWs4bxmf/fYCsbap9o0ce7I/oh5xRx
YhtNylVLWHpQ6aspkbDXpUuulA82PZJ6A4QaiOVWAQBRQAXVfUnJBSP4xlQgoePy7iCr9nru8y+7
H59EtTbp5b+wEr+6AcSf2yVY7HlVnNga+eRS7fvY0DpO913F7/gNtXUaeSBnAucJva0CpVlQX/Iq
Yt7yNx+z2Ff97mhFdCHyYyabTfeWX+EyqoWBI0ApVGgKthwhz8+idC4OU2o9vYNNRlh2ybdAty97
LHjUVSNZECV8rl/+c8pEJXb6kwDVpV/S/1W1oTIY7SWj5Bc7p/NWBOkjzuf4nqL4r0OunVM09r3q
6aGRvn+TiICPNfQLPoxsTMOpEhgL0AjGNQ/7yzAmMm38B+UhNiMwGbenuw2Hr77p2rgAQ6mdQLgV
3f6PsLvxTseq1PkY1UlfsiCwEdgvjZgwt8LeR/qaq32Tz2nIoX/mw9fQYk6hJ8qK6GOUKSjb69WM
LyMhgwkHclbOg6LAE+ghKHLK3yTXC7h6tXfQSgC6B+sqQ63FBMusKkqD7ybgSUthioDe722XvFIN
emGW+xbl/YFtxpvgvDcHN4elbK53JseqjxQbAmcOJNPVwGmhJbo9tfru4/gl2Bl+BmDbj807s6eT
Y0MLjG8YIkWI0BeK2RPfvXVq1OuNZqVO5yLtWNj0quymJfZm+wWmInCAs4rwpylLjjZ60OvWwxxQ
R58ntWxSVc+voOc++huZ4oPrVCz48/ct8n/lNiveuGqc4H29gn4sCkGS/2Im4knsl7fjMu97doaE
mnfGJ8Mp0magOtIUvEkTvkv+wk81UbL0EE3iAb2nO+QFzZkeu9hEPjFypZ313/cOBs8Q/RjFONOS
8AdH7vzRy+OhDFUmAR3K3dYN4/yRbmua/bZy8gDvbrZPhJh1VfKCR3ll94n9Y8/ttOB9t0QE5bGa
8rt1PiZR9xWR1wnkxVNxP8n0thN+aa4vQMSCgTlPSInVFrc5cgKe+JycdzYRjYkEuUKTEEjn4+c8
O4bJutQYBq/9L597yWSQF1l9noqUzJ25ZpTiiRXTXK1mq2m10MacpjLrLB6hUAuw1dFGI1ieB4vd
iv6v2yzx7eBxf39M8AfHILCqlTX/VFXkoc1gwxKWuReck0dTdv1RoN2DbflGn3DC9L8HDPwX/rmz
14/6NLI+BtS2tEZq+j32u6M+hz1CEhAG3iVIqI6f/VhIGEmZGCbwfLgBSUrtJ+e0vU8yBH15GJgl
lZ3NJUXorw2pdUbHPaZCBi5ixOI+PoyPvUEmBxX5NLkkmdUpH3GIOitq1HCV8kvnOiHWq+JNMZ6b
MwiEOisQTO8cR1/qjrkFyJxfkGv02I/HbO8QpZFXEDaXfMpIcFpDvfHs6YtvqyRjk5N+RwOINhI+
qu9UD/lZqsrdHw5hfWQqg3k/nbAZj6AAzYuR6EWjgk5QeQ9B2sgl6gvlA5ESndnG3iqnmc9S1x6h
o129Q+OgT5LDB0NtnQC4lrUFJzf6TWI6GbVWaJg7ZHfeZrnZJQepRpKOUtGcMKb8iTNIT+UF5foz
/L4odDKGGeR4uZzS3eYJdnsWUdf37l0rsZJfP3C6alnyKSN2Exp8N1Gr2cdMyYKWsuyOSlwgSFRm
2khvZFsNouq/WrRZtvk00F2BGfM+FVU9BP6BPR1tD+eMAvVrObC9ynToxK95hFLDeIl7gzkTaZNP
xZPPR44xbVqZ27zIlTRoe0GVU2bdW1F09Vw42hXfDfJrB426qY26wSgyqpG5MtrK2qK0+ui9ok4f
hER3Upqmt+TYNYSL+eFXUM/+kLRDJD1kDYdisGc3uYSao5PgGWp23/J+9uEjDEzP5lbfxqjSSxhH
w+mnO/u8exXuS432UXpf2N1sdxuGAp+s0BUib22h+Hg1u/UxterXYXSHKimZRHPcmpFLb3AcT7m8
TrX+avMQBrxsbTjiquS0lCVm6gpUVWC1AwtJ1+blu07PrHkK31Y6ynR5IQe25DhOI8g3ZqkaNt/Q
n0c+/Ox9OQ+D7cUA/K/v6TC0OOEDYEooG2w2KFE6xZAGMfpiHpoJqRe47VtSYyJjqObqE0884BdZ
3/t8nhdnsocXjEvPKCQk+S2vG8on9DZxQdkp3eXeZpmGZt9Vj8hqzGcRsREcG/dTLzMqfMjOEIuQ
6gYMygrgi9WQs/QqO17AeQ/2u1DKrC7h698dzXa3Nd6WXrEd+rxkMC0P9HVDpN07gbWU4DOvBLqG
gkKJPvNWM2l2ET1fGaDBP2gvPuiBWPWAGdKxWin8U33dIVQrNoTdXtzSYR9CDwbxFdyq3C4hL/DZ
lUGdmtS65ySIOTXIVwlKUrzBu6BgS9N596/PntSMSHvVgh6A8A+EjAq0ysI9hhsR4bsg9AwaOVVG
eJEMDlm4ZpnyJwyohH9W+cuWAmCXuiXKVTcMc+K2oTUaFsXDqmCs3eWtHwTlb0LNl5GfzwlVJe6q
MPc661VRfxByegi+/Q5uVzkvxpX4dD20bGTxJFsLCmZnEcABnFtBE5rq/MZ8dctTC8ynjPA/gH/O
A2+bMLmHJ/l+gSqzZKYS166JAL7XnXFGeeXZRa2urKKcAWV9sFOh4oow7TjJZzzZ3h02ymbEmTh1
Gqrj07axub2BVj3MXWvq1tpPbaKvFc8zm4KTzieeUGEyTX5RwZcV67As+EaHOSr+oOUv+dOpAZs0
BqoHsUz+kdFwMQl1RXfRNLYS2haFgW8Z40XIGE+hTeyxNJ1uMSNAi84xGSUOkcAfJvSHancJxwQV
5JKzl+iBpfVBFSxNrXKEhhlpp8xiCFPhhwOUkXANy13hpwfX5adzbxDfqLcNmHJ2YRqSu2xO2BzC
ctOO06F9nFkGf5Uper96Hj7dsgtO1+Nvp0R6YZTLUCj7qBd0XfmyJJIaguz8kIcE7WGwSjlpI5rh
dZsVV/igjMxZlcyfXo4/RnibErAR5n76mHNpRIBnCp/P2ABHlrLBNzMtWEdOPmZNw5BDOoT4Zodk
L/uH8JGz9y3hUwI8VjaW0WCeW7e17TJNk7ZM9/YdN59h/39HbkhQ0FXUeWJwAfYQJbyRCAKI5KIv
OOO4FhfnWHkmUe3i0RYBp7URyyd+v8X45EnD9/+Miv3C6gBTl/HzdecICILCsYX18yyz24xilh6A
u5nygr+jRGZxoIbuKkhu1M4vxGC3VAyTu1SebDP2TiwYxR1muXF+vfOaup6fGsoIQDZiIHz1kgtn
u9Q4czxd0FaF9rbgbri6nQR86ahdL/LozKOFcFKrhZLwBXz69bfMzim4HGK8kLHVchgB9ztTfUTh
i+aNBhFVIlfHc1YuyvCOfbJ9oB5MTUUp05Lj8rgIrSZgs2rnXy4qKU8tlQhvpP6FzsKsyzVtB14/
gTNxeUTbRGIEcUS0gA+QKFf2E2bRzC9QlknaTDs8N0ZAjBpbUKZjRnEsUaAT+u1/0TNlaN9Aq5U7
0MGHNQJ3Xb+eucI9XoSSG19cucMWiKaEhWOLa1KH+HGXKp7FKgmxxkH2JBf6ABRiPXoTe0KT4YJL
qL26uvWUKvCOxr67YyLXnfTU+ikEJhtOVKhYn4lP+SApgQRC6bBQ9SE2O6mNZ+YUeSYiCd+D/ExM
0pKjNzpsWon20TeN2f/MNNENG12BRnIDdfN1ZtmDZn6oa4bb39o32545ZJbJg9A24CsqcT5VtvAx
0mfbwNrWm8q5LGmqlQmty7L4rPlCW9dXI/cIVkoZ5JUSbvUkdKJj77wIaypA3+OD+twZaUwZphL4
Cd5MG8ELJS8ypd2S/V1Lmr/Qm19hNHuBALyqBJudym2VkslPj2Rml/Lc6meXwmf7QXMyTsTYJ8E6
Kw20N7ukpNe5qoJdsQ9OSjMha785BqBppJvo2itAo87ZmEMOg3vSxO8duPCkAv3W/mFL+LombhYY
g8VsWBNjmshs9qAGH+AiVlwqfjSxBBQucsa6XJDg2KcqawvnIQeZWAdy2YjA5YlkG8e29snBZLNS
/kOoEfncwmdNyr6g00zg27ZQHlmPaapYW4Z+cFvni+GJfkV3idoUhhbbhjyBcXGQbiOu2huovKX3
RRqVLFAYNzOy2e0rPjdCR37QTEvdJiKq95sdiwrJumAAZuNR976fJAR4KIB2000UlQnp5d0a/zSK
d9d+YElv0vHBaqTlQY791dVPvEPEEniSdN4zUMxF+8y1/CXPcJ/JehmBVnX3F15kQOeE0N3kS/PN
9xBLdQkAZoxXQi46g0gwn/u2ZXZV2Lxq1X+FAGGkAnrbxdcQT9Q8ZgIOcpGbBmX/lQqu4Cm51JoB
l/mD4/avcgVW9yKsoSv7MR0n9FZ22d20xsOsMaYlr9Hm+lMbbbliVaRluDlQmoQb5MmG0NIlgBmu
+eeuEw9hq6Vu5Gbzd9mqGAxco339uDzQw9YPbx7MUJjnyt4UjnXUjEp/0xWIM8LhPaDpIpWEMXJN
GGNkvbh/2ct49jlb/Zsk8QPpHQ+CTuRhOTrGJKi4KVlVjjRqEK+MCK5/ljUdmiYNWzcpODEfDBvr
hD+5MEW9afbZT1iib/teurF/8UGqc3ZnPaj/6gUDW2JWX/0Yp6DLmggTomXUV4GakhMLEULF/Ggx
Y5BK9BFMkM7N9bVupH6XdeTp/XbPhwERMyc17prXAfuppbHKGrzE69oUKmkjaoitYkb6QyPx+wVZ
8BXnJ8HfkzVO/x6Bjh0hwsQoThU1C7kmm4XxltqGdUaTEwH/wkef7HzX2ox5fuQCcHN5oruK12uZ
jWU3TYqDTUHik/Y6G0T4s5a1DhjGJ2idsPIGDdPQXSr+xfZcoWVzyVAJfdO88F2aU3p9kRypfjIT
4Xw+scW5+82Db+5OyQkzDop/SN/D1E4uj735k2IpZxtG3tI0KK390FWyPgKALhJeeqsQ1gYTj6zU
IYLjy22y2H/xKcv0ivYk5Ea0ANNNu3s9bvYEXfw74HtcZwtNvTF/DBcIGbShj7AyAd7SPGIOVpGk
OzWKaylEUwKkYvBODUGlV6L6w/qrsZ99Ercl46yEu1HG4zI/0Tkx6zXSoanQgqpy92fdrmEhpkke
SBmKhrIy+zFiUlUwl538CjTMsaZtk0U23MeDff7h3ysU4pMJRrEEAZiIRTeE17QdxjKwgdS957I4
MhotHco5wzBkt24cSZhYlj8IKkiIps11vOPqlJ1ZDIFo6OtzrGuuUXQk9A6Z+cqmI0YrF+0AJucw
Z5pE/XVrL1ldLQJxTSM3WOiiRMYuHSkJuSYJsaC5lRZsoWKvoEyO82hZUrTg9HBbN4tiK+lEzr44
+QTcbEkOUlh1BMEiQCGEeFRxfh33ikPsZEVc5F2wCA4+qrpL47JOgPQ0txKVj1NCN/3hrpsnG9SC
lp/qCZNQffXYxAFEsJpA7v4T1AVhVS1ITNHbtueFBRSUmyJCqLwuPDiaeQEllBbAXNmCj3fsLUbu
zmspdiMStjp9FNwK5YjbNjjlyIzb+ysIoeAyBtrXsJBSl5Rb/BZLBYy+eU3GlgW1IDmWdoexuw07
3jugYtDA0hgXo1yA3mXuWmSzBJ3Zwa4J/73l+Chn95CiPU5hPl51QGpaHy90QaWLvR+Jm4kcc611
+BECo8n9k1TSzTOgKadFttIT9q7DAM1aI8fII0ChqDwyh2NU9/9dga1c2/6i7A4mP9T/z+uQZDyr
Sf70X5c99D8nFf+R5rz4aALlxwDYS/cPMwCp9rHa1txRuzptbC8g5KouH0BZH7UqMFbbLwkEeYxD
PU1EVcTDQWCqbhvN+bU25ULl2/HNYXwDILYMhpF9TKe761uYxrPINfTixxVDL6wxZp+57cOhBk9g
unzkirm/42ZF6hPcCcicS0AdqdZKjjuy28RnqBJya58wNDARBAodsU+Y9JBjB5jjdYtn0g7MrrPR
1gLg/M4Gn6OVj52jCUqbB/MS0D1bfEk0wfP/HT4/Xz3DwVvBYKMQSAP1fQCdTViwmY/jA9oyxuRg
d8uFKh9GFf/hiBSeIdYO0rfAFDKNf3qTdqgh8oKZcLONC/fMMVds/eEhzVunbdrKhHHya3F+WnJR
/ZfA2F6aGCz3BRf95i51TQNzaCjuPA4SLWXzMarUs7gTr+x4Whf2fwVUMdvXy6G+JtKU1e7p6l0Y
0XapTID0EYGA2pqLuAyH6NhdeQ8wZnAcUJ+tK2O4uqnib3RkNltTfRLF03x4tR2sTYe9oWLtPZc+
bESMaLcFdl/8TgAtuGQXVMIawSLLLDUwwCCD7a5pCe80XpHFqEHPhyuKef/Qu+jz76FktX4tQC1v
m/3gqZ0CR4vzrPjd7Y3F6AHvr613h/JFg8EFku/MZW+4W7ZX7rlFmZmlJ8x6h9pFDL+XbC4PL7d0
au2afI/cc7w3TmFqLhObIO8ZFLxrVWLt2yKn0MliGfHH2s4OhCJ/ROodRRIX3mBkVChqIug9xYaZ
Mlsxt9QA5NLNzM+W22XaCiBg/5Xh7N0f4l4R/78XtZzPgnHd1jLaUHzP8bBOH2BxXizdUi/ufqZA
/BkyMOckr9iF+q73V1rpJEbC3J6jNLE9kliLC7DP8RGdtzQJUrf2RADNtCxWKppGh3h5r1U1W7xS
wQbfcHoEGFFXKWfeg89zYl9ZglYn/PJBQ4AbJYJEgB3qr4bq7TZnXeBh1kqxxbcCGmuPbSdd6NGP
RYBg8QjFleMebNqndy13HJfkVWKbJ5bNyrwyqHeK81D4n0RRzaZTv08NeKn/ROFLcigGFqv0gBcG
yB+/LrOuachKggiAUiUP42ArZQNd30u1WMqVc2s+GmBpkQb7etw7USnScWNGOk/mytsIvrK27hc9
AIqz5onjgGM/pTy4M+XPX5a36POYJGszDvdev3++KMBQ30s2t309ovO7z8m09Yx5gRyUmwjna6NZ
I4CIppzV+ueFCrXvrchqYSrprnbL5W7yRrn77vxFaUDBLM/S6u7MGifcscmqNWDhNukP7Fbnq7uF
Nk9sKbHA394z3vRV10RWpx6BWKsQu8LJcV/1psbXBLTYNveARE5HupTNF5mfc9FDoN4EHsEMOBGC
sPqkHbKJAgCnMywbm4J8d0uZblQC+HvnKtV2+x6FZSlHTKB+ECXwr2661myWmM5Fi1Ms8MCfsytl
DXDPcts8x0zN0L1m3m2MTjfKOPvwJnlH3DJdfNPMDuWOiw0pH1Wk4IAw5HGRyf1yHZ5IWpVkuTFK
qXhd2cnpA/E5b9rcMs0KCJRLmuZZBLp8oynP9voE19arh5P79FHmXv7AxJL2AyiMCiHfWnAQJlVy
koM2WA2ElyXFu/p40NuQD/RKF00rjuCgpJSYKwkGC1cMOcbeovFPxjK0GDbizQNzP6Ze6GqzDILZ
DXtRy7PUcmAgUTHTtvS+5OlgCYv9iuGTrtb9KdvuX05ZmixO1pW+JOWcjQjgid4aQWNtgso6Fkz0
7l0a1rtX4XA4UD9LaM8Ghx7qHN1U01hREOP6lHVTZLR1nfEZLcd3hYIFegf/aBMP76Uu3YWHGFfg
ZCGqwvPV5xtasAcuy7Nrr/DsUd6o/3Q55/2WBCYDvu2DJnK5YN3xbGzgZeJ6dIaBl4WKNqyzifeh
IQuRs2z9Nn3WYJ1Cg9vwrde8D46KnPW0RxWfI67fBhvkQwfCQucXol5nf8ZsEMld+yH4py0K3SeQ
EX6KVZFauLc5c4J2UQ7NsOF/qZxXBLTKeY+xxKFe03ap8X3ztH3u6JA3I2p1Uw4GjGVs2sp58791
OV/6Q0zBXOrH5Y9qsmNhhK7jkIzR92B6yUhNSEu/do3ffutPSyoYe/Kq6K37NM+gB696mPaWhFdq
jZwcp135N38HfC839bSBXvJvlk40CA24n4n6gw0+KZKDvV5Vzvi/kE1Yx3NMjerSZURz4sWDx6Ab
Q9L2PYCLT6HbAPPgme374IcriiFjz9zZYzNnSQYw0keyUWYnXJKxeb7Q2I2YpAVh7cbUnUIQ35lf
k0qEfFd8C1s0IyrEcCHJwe/I0NvTasrC0WI6daFClzi0BzyEz+Q0dOdL0xhGZbBD2rwrMQP4N5N3
j00BqOuXgnyynKSh18t75+D9kZETKtEi5kzqXaodtlc+zIulG/eL9h1JP3CKcprfixAFd9Sa8JCS
+FFfJbEl2O4HCZZWRK1+UoRZue0cuBOOhUJSyBaoS19BIzXJCrdE2QocP/6YUDs9s6m8dbcKv6bi
NrCluMI0tQDs+VIVLn7rirGjym07CwdHNxrWzXkwPnmOyVGnRGn9JOCC05pX4ZZEPIJiAaliwpyi
g2Tm5kTWhwZYS7Q41tdi7Lbqig40Pb15EAlr+f6XYG/YMuVelO+rXWjFGWrOYZ8C+CcXyliauqNa
z7VtyPoR8TtQUadvT1QeXLI7YwCfBHbuqyPxRtR+4xHzVjierBpAZdjpYnk169YTEq22gm+NyWp3
h9qpaiqwDrQbbNp0sWKhSDD4ckro7SPTDcI1BqGKAmdf7jrMeGnHZNYUx6R/GJhK/a1fq3y3g8/p
HFGk3W6XHV3jLtuOvVGf2EH+zJZ9vPbdRvg5Axm2MMgMW3ExEj+OPaynzIrF6yiGa1pGDaccc3S6
xOdWgZeCzD3iALD6Df0xsqan4fwwr+i5Jh7pdErt+d2QcWpbrmzquIUn383ko8nTslgw+WloNtit
tlBOZP3XYHlRDxL12962Kh1spExGHNQaZ8TP0rgo202jaL9YXPN+MMAmh/+YDaUfucCV5iV/LIvg
0ruVrnI4w4kYsbD3Vd3uG+EyYrdBodry9BJzP5V2cjstdK6tmg+ssM+SbNw1j7F/4ZzN7aWhwTSB
J7169xcEetM4Lx0uXrDeRn4XkYpOkxRRMT44KGmmAXzep7MCMxGPa9z6UqAwZCkxmA4meVJaaUNB
p7YdQpCofbPSZIdjnppQj+Q31GqBrftBSsVzX0juOGpyx15/OyZyT+n/Z3Y0BhjiUEzQ76bPDnPf
1W8MvyA/5AnCRJpeOaR105MEEa/K+YC9Id1gJUiTnW8FJQtomZjQGufs05mkl2BaGpk+0OJ644lm
8eoY9YidtRJt0YId83ktLXO/XxTXxuGuLn92TNOipBVjGCHUA4uv5mS6YGE5fnqK3wJIboV21cnX
DONo1upngDnvPAzYUzPD/NG8PrjrHumgfMijUDiAAUxQiG0voKjj1H5DTHP5j9/JNSCJ+M5qHaNw
UyzBIVFVNcKUq+MOE9gFoufpSZjQQMljZ/1w65VNApbY8zdPVx943cgXdNG8At4OzBx5xw+3vNHm
4oZtsoOPh9rNnJDQ0jgJEbYjDtjwT6WDuYTR3biGZalivM2oO9p3YJftRLyUBnvdssIPumN0Blwi
f3EIZ6uuLdxvCUgd8u2Zom7HXIYwnviM8LWHvRX27O+tlBBFvmD7WhN6glW+mC4c7LIaH4Ypfdh4
vqYYtMA22SiAxlwQvF242kXzMbxvrmlpPp7cZakyf8jEhIRcLw/IVy9VintnUuXGVH1dvSMIfyqO
/mxH0/H+mMEibOqFJ+OaSI0XCOUrsoYBp8bY5kKWhzT+NYC9+QBL+mqfQ03oKdz6WysbZLfToIrZ
Vyn9mpuHpPfAlYF7lJFcXa9YsCgULu/UHcyLAE6JzPFOkIGgiYQ4y3g12Tbg7UdbKMQewnaXEobn
VTk2GZow9UHFrPoNoYxkvL32Yk9SdTiutmkW0/YFbZlm/NLuY8zQBFYMIr9R8gzaeq+ZtNy7YrVf
mU1YmoBZAKq+2RfTtC92tHafDnC/Rg8IwUGoNIwKm9rvlQurRq/4+dEINlpQj2Fk0fZ/4IqNpT2n
rATW7v2LgOvsobJWtisMUQunqHjbE9M2RaWDwWTJH2fZKlEcYmtI4K0gPi2IPeYCHSbP+4ebVITK
SwETk5Zvv1DucA4xG9yko1ny3QY9H5qIJ+ZhJprjEz+qRdvBfCJCsmyXuhh7Cm2KmeWLbg1yK8Xh
nMlBl1zR9UEOpywU7ecy/I37kSjCpgBvL3SD+pFrSp3m4vbwjOb4KPGCluUEkTrFmJ4eDNdv/iZZ
LZtBsPz5E2FAX+G8Q1Rwi5qz5wXdLrsAjhIg5P81CjAhrXhisZqD9R1R7gQqiJiX6hFt9Cc8s4Kx
jcVwtotdYMxQCe+tzEl6Igq7DUCUUm36jMRsP9QUfSVAlMmHu0nuHLKBy1ZAvwpf7WVAbGXHr7Mg
WHvswZdi5/qsc7ROx44NsdhRcbWJwbQ/7ciPHuzA2EG2UBytjaTi6QmgSi0DJ+sXfDWaYn4NE1Rz
u/WtabVkvKVNrrM9tGaKfG6rqJ2M//WxtmAiqNSkV6RWBO3uf4xYJlaJnADYT4ByP2PzFkcSWOTl
0pv0pBqW8COI2kSJkYo0+OPmYjP/R2h7Iy2rNDf8knEGn3vNXRtcVzYfvERdCAiQ/VgYCtIKSagw
LXyCkrBkeZPyAJR0K0pNaJrxOuDbAEHwWOF3rKLc2I2wDS6g2DvjaXon64h0uGpAUUIDgeTMPPH5
0f/sKf4QGcHjJrd+SgjahY9nuRunRK9NXfzpA+yHh3VmDsql7i7F7Sy1f25As/y0u5DXTZ9GW0i9
MAsT47eNdsejXKJtpqsf5OifIgXbtRgV1NMPR6Ob1yAMnl9WtixKyEGVNIdgTsNSNZKyHWGoITbm
JPQeUfxPVw8Ag16Hz1naFG4WhOeP04DobvykhDYf9c94aQRLUl6ADN6Sj1qp+b3qAwhMhYy2AD3o
lU38yVGpPyCszjGzmUr3RQHoGeUi0d+HmNcgUwCMwrzpcGFRsA/nmT5acV+q0hHIe6Xv8t87p7XK
d2E1e37ywJJXzMbDW48+AhWLZfJKNiCyDH2DuHIBhIJVIvE5ugS9sltWjJwmyHe70pq1/8hSx5d+
aYLX/B9ufAfDN0dRE7xGgYZ/ufxlrn8ysw5t6+dIn/R/rinJLHSGuahEoerpR1RxjaGg6g11hzKq
VTUr/n2MkH+840AawebxqkZbfIdRFP02DdVV30aOISoji13A++lzYwMoqIjljOejYVm4ejKCoH7e
0HhC2gCTrP/4XngBqUHmEaUG5VX/otQDPfxIGx3szlWWKOptlHV6x+M7TQY+SZ5IEx5zcChEVSlg
WmtyHfxXhO6PNR2zW20QUvgE2wtHf5E/9jE9yES0tcPB0W+i31/opSv40qaFIi0rfknjzVfiDdJl
UzY5EXfjyb8MRstLTjY0rcY3md1k7cBiIH1U9jPM/IQeL8U3HoMChnDAT9+Scj8/Lhz7YPhIPpvi
7G0PS6bsyMep+GAbR/rp2QOhJMXww5LjPRfL/R3SNmMl+PfH+3EyAthk7r8CCK8bd+dSar5Q4NJZ
LkCp/VH6eneYdSOjWpnQ9AbwHoIdWIO8dSbW1Z8FACL4Jt3r3DR12AXvm0nILwDuWK7LErET9F1C
vD7CkghM/tVy+FE2l3Cg1RyC2MS2oFYMbaxr1KnqcKN4iAFFYorVz6AtAPAFJ29pF9ZA+nx+Rk4g
U8JWdJ1ZQQMczCCtsLA9AOboPal4Hk2Rue9aNes3Yb+wo3wbAbtAjHLG8ddOH2/83C/7Cb4P1nE3
Y8AkJFI5X0AVhhDnhkJvtPe0WT1wNjtDEWdpBfdk3MCa5ZWLbOzkxS1soq20tHkj/AoYAQLIrvVv
Qr28BasTILQnvlzydg3RDssSMqJNjmDiSwhSqMK4tO6X/ZjY3V1e2uBIti7gkRUjsEUXsrxYqvZn
Xj8jUR9JG1Mq3eABPu472rfuCaxJ42rDTXsihsFO9iCF5mQFErGtfKpzxvGhhPjMTwca5NCex1uL
jJ3iLumsbEM34FS2T3AwrTibKFpm1ajayOo99g9Tk6+tdYCEYdCpgWtEt9iR0AD8fTbT5cIRxY2J
GxKYDpGoZUvDDH54B9wahrWq1CPqVOq1P1xub7zL8+DBC9URl3YUlSnLrZAR+/x9Vux95bWLEf4F
MbT1GEanWfueDNe00VuAm6O9Wf/d+2rZ/erkXnS10BsJMmwydSt/s6KvhviWICUn9dNDe5uiSDM7
bIRawGPbUZaLKNzrmhhL9ycloEd3lo5fv4YLvvtK3aYj4wwyVaFe42D9z4pLWhPbHHajB2S/bbYO
kmhKxAwZ/wj+ipv0GV66d+R83btiqefwQwEuyPqrSKY2lNakrzOftS9xlHg4BCZPO5ydyq8hkdQZ
kXDvZtVh5LkvYTgFEfl2vRhg2ZCUQhXSNwspjkOGt0sq0zlMVirgFVnviueJuctEH1OPqjwr1k7Z
rVmSzmr+OLt2KSMj/kr7BF+l0StfZoMMyetW3q0A1w0X3kgmyJ6ccOKBdMoszhkHSj6+EsUtbCgE
ZeJsqYTmlgwWLzDbso8PnQyPGOB7NH1aLHFsvNkAnT1wCl1AG8yMucxRRrfos0A8f8Pt0vFwXMOt
k2WIJqta71fr+UXbdvqrNE7zt8L1p49CqGUVxT3qw4sv4BbPDs+mkuM7vfNKlYKRQxLHOBZywDlR
d8ImKg9mhTHd69wrLPn3Jwwz2C2nukVRFefKRjgICtFb8E8Xrnt7GxjPek8FN8AmE9O3g+WEojBx
5DnQxQmrMjvSmBqy+e9HFuQjgY0dIS4LjNxk7ZjaQKhwwT/8eAGa1D+SFCo1m6839dlgocVoHTTW
UZTaII5mgy++tUmoKGm0abo6fo+PJh7KHTb6eC4zgEw/lKEfsqcOyuM1Gid0BNp2B5dnTAIdvUQ2
/2/N4X5xkDyN/StkZ5gzSjkN6TfpDeaiiGqUo+3b7xXpdYi9vWiJHZ/SxWiqiGLx96kSqEn572oX
VLIMikBV7U4ZMZb5TtqxideyVYnkOhvlKGJhj7nrA5NU8foaOLjbMxsou0oELBOPU6uCThmcJPoW
U6jsnpeZsdXb11YebG3kNfhjP38W33R0u/0XcO919r4iEYNrqxlE1tKlOIwz+FlJoQ3RKdMK2Cgp
S9PDxGuNxPyyIzL/HiLfHgc5ysXaviStz9MoDeO053zQEMOOq3IhsgsSQDL0tOEWur7br1MUpy1B
eB1XnqDeHVwxn/73532XrnGUFF+YnvLDA4rUMlWhNaPA+c4D1U+z+Uuwvu2CoRBh6b668SVk+Dcd
hH+2vsSncL8Z59OBcrMV7JBNjrHQYqAteuButpZkhTM/qmwK8DpW0nT/SbkPB1pSu37mbjSlbHrW
4dWZP4UeVM0zV2M71WLrfcYK/EsJmtn6KAsfFPZrvcy6ZEHq7HGZjOZu/EssE0LSdits3ZngKo1q
81HUrhmaK456Ld371SbsveAk9eiCz2FrcV3xBwQWxgoFOJdR1MuRID6vYiCaXfoMAJ7rZgNoyC9S
z4olhtselJRsP1pLlkpB2/2OwMgmktFmYM5CsDWxZnteWLpGsNyKpXiw9eH699q5zrYBG7sFMM2M
V3UvDGLc2zbNgmQyNCYz6NVS9gpj4c6thEJ+xInX3tjKWKTOzmQJ+qFADcGPK9ZoEvTtOArMpGjm
4zxUJ8YTCdnB5yMVPQ5xijJWTRGYX6ByZGmg9WUa9qDlzFP0dY4URyBn2mwoKMs6gEMlkhhwH+Mp
CLq+43UBGTktWAVw5SrRM8rtzyK1EEJHoSCPriI13hvmToZa2J4SvBtxOAZhCEQmon8/IKNgyi0R
coETtsiaM+k8QodVMLULCJe2evMGmiLmfauVpPlZOZ3Cy3kGxOBvCgQKNhx62qekLfpy9s2uvwfF
SIxYdXkYK6ezFQH64SzPGwwYYG+GNuJDw3u1A0znHGNI7G4DSpeQAJiuQg/DjES0UszIwIvVYfnE
djj3F6CXK+2EHr/6Ke9/yiJeh/6hLd5szW45IMjW7W33MhCFBwqtm8X0XYz9Wd30qNKapB4NkBgS
C3mLnhNqf+Scswug1VA+6gPv3qH20UV1LsbLnyn2n0i9UyZCwhFZTY8NdyDrMigTUA3bBEV2iR75
pJDqQiTYxPi50Po7sOPmeh8bOHolhhpGI/JGrU7wG+y/i6/Y37zVgvxtfK1ekG2J6cHbczOdCgGl
H2esHkyF2HlgExh+dEpWY9r048dHre7mW3Zh6PvibckbRH4INTm8dHmTWRYeVBWDYfciNcIpeEuu
1+k4G63rhM5KGfYSP8SYBt9ynAesmDvcblRL5V5JzJB9TmxFJOyM8792bnSt+Rf6fgzFELrcktxg
xd/GJpt5HfKPyOxzqGWRCcOETnMhauG1txH935wHsZ67McQyjIN7Nvv0zUU6Dh/Wz0xR2gcQB6wu
krzksPhmEmDlvoBee05CwTvc8QeKXtHnxUzGMC4+8zUCvrgZgvPDmJBT7AcsWjj9HqVNC64z37AY
o8lBYaxydYmz6OFWXx98UwdTjOyGXPQV02BURJai4QdgU11E4aLtc7d/eL/SllSx5R18bMYnNvOO
iGg8wTlxVO5Rp+MuzPCXc0r4QF+WavWOSQKYvRbgpR9AqH+hsoR0ZiDuSoEHLMDzXe5jP9PVC0Bw
hBbL2It7PCA99GUJD5mlAYWovGtZussP8jvqQEN0kBmKB4G80Ow/RO1IZvndC0Z+IecD/d5Mpokg
p1qL3haWQQdE5IhfpMV20rx41s9ZEsbi5eVp6unayiqxbSHUt0KT2qgr+ZHCqQZ4BWTil15SqhoE
ajMjtaUto6lXBiAI+XaEWfeNcLQu32nO5592Y0//hdamU6/8+jY8sc30Hp47YrFiZzMHYl+btghW
y8Yf3gBZygcFfukMQeiDhUIGpJhNNR8RewJraGKQEUpjWC8ASAMuOe90Hu5lnHhiHq4f8tHYDTfM
hEcDNIesgQQNOxswdRkEdZxGukdJS3owpUcjSqGIihTTDAB/7i0j+pIp1BkRALJ7uoW8VG/VqnXY
UP/qmtBGYllabBoqv25fM3lchRm8pajuf8bRQjkmFLdN9VBfod5qK8sA1IYCXpdTP/8PT+ncc+v4
NexNVdR1Til2k0g6TeaemahsLsw0mfF/jN4idNK8fZ/EyNdPcrkOeENbYDiKQ4scYy/+GZScha3l
K2EVV7zUPzY2DRcxt9Iv+9dR1klf5RMGE+qzo5N84VWLQ5mu6lP5DvLUD8OoMRWdTUHI7bYcfPDX
l/Y+PvmfScgII2CFMNZQ4z8i6nBdCe18naS2XVWMUs2CIYmsKijeT3WHW6JkfIpVDEJQGDtKLe/R
WelfAUL8wW/fp9o2bWSgbMwpvKxKpNOhQ13pSjmU3vkcYvzkrMi547fCIUu7SIe5xgL8kMRPaf2B
328AwKmUY/r2Rri92pK9zJV1r67az+mB9tGs+WXM+zXDTQVQn0oIobCq5sPxk+KuGguV/J6X6qin
yDGjm+7Mvba7oFe95i6Dih1UfoAyw9cYVo63hU3iUbiLbThXmaLSCXR9Ye+LL9p01VfW2xK9TlEP
FB4v/BsN1oYnVV6jJMT6ztNrM4G1CjwORQvHKyd91JvAmNf0FRRntdm++f61ywEbhh8k+MrdqIcv
WR2LzMINM0MpqM2Dz9kzBW/u8D+8lmXqSCkCmm1uHahNJKufdX3pC3qKNpOmlPU2+SXBtN/toikr
yFPPxeEjPb1+/7k+2fqaA8zq7zbXChh8z5+0q700/cT8/Bu/PNHgcuBnrUZ8Imv/bdS69nXkGCkS
Uu42lmw6AeyYvoWSScE/Smunl4khus0YatUDPdgvVHBxrUy7Y0aDEHQRlHHws0qY174ltVykz0Mz
XS+AHTEUGJetL5pzES0UU2LZvt8Y/7EevgON/gssaaSSp2wW0WbuCvnrh3Ie2lVkpybbHy4cMlGW
EAZb8WGry59ZBqwy80xykCqVWNNfLOpa5ISxgA6zAeH4PrNxRplxhJvc0WCHNSJiFEYh7AxFTFxL
fQ6c6K8kjQNU44unsgxviv2kbxFvQ/83UBnodP6r84Lnx7uSnoZacQzI6lJxgqb+2eoYXg7orODO
iYWDRBNGQH88AONJzv6zEbjjOTRRxR0J46j5FY+PzvUtQGiqzfYSPw96ce4Uog/4flLhaQJHwx1L
WbO/q+0SkXJBNXtT1BwdXKlG/UNW5F9PxWctYafW/zIfaRFXpp4I2OQqvw04/zr4E711XpqFnyTe
hbREBB+YtjpInpZN3uo3eLw1PbUzMoOPRdx+ruNgX+OOLPTezAR10ipXPUv8xt9jUbMETeiJlsdW
0jJKJT0/dOg6iWyhAdE/KNd3MklCe468REZ9IFb/bZ7shY8j5vot/bSZQBDQovDuNRjmJIjDNU01
8TDJUOYFfcJEHAhE+5QkrP2YWFc8/mzQJc4qW763RbvuuCocQCkXuUITG5MWo/TkPp1rf5cjBezs
SphyvYyuPAcIEzTlxzbC0/X1FmOLzFGnB2dEPUVIE4i7I1BjlFWS7VTW2EaI3cHFmhpSyVCsG3Yh
jdRKpSfvEArVk6URoT2sPDXuSXlVUK8+1D/elUOp+n0VpBuZmU/CF1fF8lux1c4HmcNH0NUx8N/s
bKJ47u0lN2C9dP1SSTwgUWmuEewKV85jzbjUNc0vZA8lK+0bOhg8ngdOzxwb3iyWIFTNXJiWT1kS
RpcgEJf8d0EzHSbGG8lYdnIM9haS0Gar4MDBYBE319fVyuKNK4NExTyhvz4I8on2yVJT6LeXeMW8
sTn/RKRx8Nx5tUfOyYZAqW/3RR5Nv4mEgLpOZsv35O0sMDmpteqwDoshElJ14VcmMfxCupdLJz/a
m+t6ANCaTu6yJDpGLV6d/A2PeqBNz1V4frR0pUuG/d0EBsgNDSwRB2J1E5De2wX/W1/CDQUi0WIR
GBeUQk7zBlFNK+vbBBm0Q9vhpR9bC3oj49f9mci9mh5ZfIQmpBfj2UMtKKcDSdv0bDNV0ttl8gZQ
glsUNhhnxIfEwLk1RoBhZkeGyDpiEyItE/hCU2VgZN8IR6NUKUX9tRxyhRZh6Q+5gE5PpS22nLI8
kHucW+Jrnb6t53rw4earTZjIXIUkPiKAQai6Kg0lpHeEGVuqiJd+7CkTU/tiRS2iTsXvnZNL+meR
buiVKgOa+Z1V/yc8u+JV+WclqaDB0c/MJkYDNXYBHRmjvNfUVq3xkopTBRu3H+GEJY+cMjmHmxW1
D6cplCyhRATpMeJMRiS7xyTdVNzW/8DZ5/nuK4PzWu7jBdJZ6BVrPREYBta0h483JMXjqhFuE/gE
iGLTmHUHVsHYqHtRzrWVcvU1gX2ISXEowY5yedAYEcH8+Adyx7ZpOLLG7wZ3jnCrmOCyQidXLPfG
2eUg2IDC/3gLp/jDdFEuu5WLUrPft0cDz7SZ5QbFpXKBICp2uuPZOex+SxR9onsheh7IDZOdiu53
1Cl9UxFsOA+UVQvINvw03xJxg/HI+U2SL8YTUcdYBFF/FTilELLWE/dVKhKj0s/jgb2qOMMmCnSt
7ok2CnYnnU/h7tDVaIJy0fVsnHcA+jv1mckCtLS2demw/zjPDKV852CJin95ToLvEH5pYpM8tIS2
gecEoLSl9fQwyRQN981RYmk/taAww44+jD6JKCYQoArie3p1hw3yOaKmSFKN5+AWWdvFhQYBhPg3
KROdMDO2OYpBX4USqzyPMFzNY1G/P47aT6FGctohGH05Kw0unzLgfM03VQdq0e0gMp0g3dJFsFDE
aUxBSe5DZQ926h+B/Zdb+wFtiW6WfxC9MEOJYpVegVDxsZ45w6z3cj7oy6aUy8ygNw5M0uEL4Vha
9UfAAVsHy4D9BONLG5AcSklkFqDMsiOMcLtRsEDx2vqVRzFvKrdd5UsfE668mna2qCXxenl4n9zF
mQQMfetkWxrhrVb2smiIfOYuP08ggTgFsFQ7Btr1gVyt+ObdwteyyyZpDPCGVVBwPOsgQ20fH29d
zkTTYCJE1qH7tk4NWFIiVQ0PNCMk4nJOqNHsw8rLCSkoa/ycSb4FpFIP6oS80TC0wlElHbhf0nnA
mSmzEo9ulwrGIAekuzgYzrQBjKcvXFN5grftCaHyHO0oa2Qk5Bn6rlokz5MGg1ZGceJYe8iOhYtd
pS5xUwQ5UVRQr8J3OlPd4nnrr+OnzuyukeKWqTS2VKYIkeKEm5kBxKTQNJpKapDhYUHfKFNC9lBL
CEkU0fcFwSk33AgvkYlVClMilqT7LvNanheQNoDZIkrQJ8GLaA/VFCaXo5TmTXnXLuImBD4I15nn
RCBV2/0AwvQHgjoPprQ9zJ6c79B/ciB7m5FacF6sNHt+yIq7LwD/rdesQwiQfby2edap+6lUkzg/
MBmXFpx1WTi2JBX1FrO3cIRMDQr2uIkafaqg0JcyglcMtHgwOS/lr5U6UmgcX2VylUUHoIJBh/k8
0ih1A6X/6R350dMP9ZJpPp1Zkr4hasc7ntKZ7PgTcMQy8uWK2doMzUUPnMDEcDvfiBMq5+9QnuVX
Idn5wSpTruBsMS5d9XhTHTwdUQYADqvN1Fh35em4K5H1O2n0gHAE48G837dLFNaipS1+O+WQZRK7
exZiqU+8x2oKHtcytOUWzKNcBnoKEqT/EzYEvCVNaDCVDhKgm/V+yOxDbsZx46gHWAKQBl0q0MbC
DpGkn+aK8SIo6dcqFcNkQ2FmhbIcv8Nnc0W2xSA8MeCdWaBFao/eqtMvLue4ZdAoKOgNROikToo/
2CY4DbAgbRQeAaQALl3lOX6LwxhWGVfLBxkUjZZJ18pK3skJHQ1Ew+Q/casXFuA8xN3zHDo3jHKU
Js36PHSjwpfYRQg89T/4R/A8fk8qhqHTNRAvQ1oz5+YR5MExLadyvEV7SBnEqFUdp+4MVKFja5ij
IjoLvRKvMIEMDj1EI5sbgRPX++c7AiQ2hxxxyXawjZfcEqAS1R5RGAX3b1mfFeZj8caEU+PpSf+K
Jiwt/Pe+PConBiUFR8HuVlHgMrhGIrWtzcQRxhk9yoj42DIzeT+NrnHTTHhJXfpMQW+1KIQW4eKI
qzw7309ocXuHUmle9itYCFAeDxEBXMNwb4vsVOy32zFFnOW0nlVpxrBKdsToVjBUh/t3c/K/VblF
f9UUu9Bt+A0OdVogXNiO2afTD3//vHgoeY/J5kf5OsifxG80UYv0M+zH57NzmyV96hepJpp1Rius
Do5TQIvxgsc7+/ZofUAOxMezXx6gA/2QmAF3m9tWbWKnOm/TnVPRoWjC1HYu36elGor5ixM6J7T2
bXSLjlX7nN5vpA3Z79rvgvBrH9RgMN+IfjjkCZtd3DekJmZkmDe2C+n9XWjWXymrEkM2A5WcBZrt
mmx2gtEx3XiXXZbGVYHbUW3CdyPz8ylVgE2GGJzzfwISKcWoD1dT7xzLgS++/fM5MckowYq4doLo
z8B5h/YNkTaEggOgBVQpzUQXsdX9HJAlVGKM7kfkRP17zEgtkSHKP04kO5FunRQuO5LNeYq9Zhmp
3Xvgm5uEnRR/15cXiHqh+HUnvxjUt7mUSsNTaOGbAUYJrBsoc8J3gtAPuHNN+DFoVIdgNasu5mbM
BdryOW9PKZb6n2sF4q+X3DDeMCV20eP/ufa0K8tD8YXYuT0ZOd9Oca36HbjMsqF295SGti3m448x
lJlbyQUUSYpL5dUR5z/hS6VJeLgowz8J5vqEqWtxomH5d5vxlnQpfgmIOULddnGMFaMNxQFUYmVM
BUeCUmpxGCY8QOk4o0S5c9AJZslLr2MPCgbRVkRjdEVjjxMV4swjlOgevDEy0h2O26zqWEqpXex1
hTC1NVz396nHWnsoFcNmIaznAXV2hUDfpVJ/o+dhoijFoUaW3LI0QJRA6W436vfsRxT2boVlVrbg
aQpZ2EyF1yxSPgdVY5kg8sp4pp+7eHBpsbfkRn02RGwSyRqYM7tkqWsUbEnkVVxBYiRnoGyKx9Hu
uoED6VYQdA6l/tX7QxRyG4F1xKHFeHJCVPGWexFDUJBZc+hgU2hFZQGT30hXzjzxL6pfuiqD299m
nAQygHY5eQdXDScf1NbV2NmA/QDokeVhPULuKVdKm7SsGwmygGyE73f66d6vad1K0yhqKcoUcCr8
114Fs9UtcOJwcb125hd7S2Syd/Er8S+dAh0MvmWWF7XYN7g5xrkfh56HegoUvpOP2LEXwQl1dhcG
CXr7CEda/7YoNcLhRBm5qEG/ytPju/KVOSOoAbYeykGT3mioHGy8AnKpJvx1+GfBFKGnD0VPRQ4K
09c0IX2y1Hg2ZzpqgWtzgHRD7V4yl7MwSjVWfDhpIloK6cVB4A3U9qx45lrOTGsgTFjOdKRrkb90
tQXMWsMj6MJGyGuE53paYc19AURyqqtkdvEzmhmKUy9eHN+y9u9EzG76H6fQ83p5/5MDVqVCLPX5
LK2F1+joj1NglebAfv7kMPj6WrIedkqwaEBUsow5CJpkFLJGSymPPYno1Weftw8wHqoNqwjc3V6c
5TBBF78BkJMtDxYB9iDP67A5vf29LnNF+nu5Az7wTGWXp9r75zM2IAc0GRTLg48J45obD42JoPxC
fGkL7bRT8E0nm1BdbNoRBx9QBUxpMxj6IU6Uo/nhG+QBl66n+R+9562Brbaqx8cIxxsrL0B5wzgP
RoRpJ5EDEMcdwnHo43LPfE1ghtKgAJam2Tzy5W6OniZyFRrszMT/Lnuc5erZIVMqg4GcSrehiKQM
T4ThpGTXJ5yb7SULVc8FRWxUHlpD0yuuw1QHLZX+kWXvqjWFAMnf4gonu8C+OFU/ENnqeY+2phGi
fRKRDY+QwsHzUoq9F5afY+Wm8IkSca+ptBCrkdzwto7Po44xGjaMscc4PgM4+cQQTkCil4puu6dP
45CKaUJ+wPKgtHk/47bJHZPtORewTo1xF3SVWrG8q/dmk/vNgQBcv23LtZ98bnVGfcKgTrwqqaZB
AivKtt4jEo982x3GV7Hd2+cp6653E/Idctm3CIxbiBNgBWD9mrXJBOMXhSycRnDVkgG2gsCdTPdd
OEBVM4G3/5QTKgDeYeSzCTK4/lZ3eG43CZvyw1LFoOQutCMsJsqgsMq2MiTNqwsi56GWGbmUZpoe
EM7luoDtmUr6shHZ5m4ykbdcXdfwYkAFRXKaVDc/dXvUE9393vpjLTsq0zwKT8cNhVToC8KjC9Uj
X/Nu3AKxrrxnl4S8x3ui5c2dJAqNKjvcV1tt/hB0IjGt5uFoORzaTQ5amWNIXWMz2ymGmF8TFVaF
amHA4GpNDlDVCyhhlP78jIWzHG/NCyA/8HCBcqM8ES1OIQzQq3IH5e8oYFNqaC5FRZQRdZmRpjtk
lls2LmbyG46W5RuetypIH5UBOpAIV13ZP/a8b70gnQP5bd/N9eC1Y8BGJIDTBB5PlMj+Vnln9GOT
z7h7x6MXrPasdB7aQM0uDpJERo7dr0PRBS99IfKooeQ5LoMvGwspdPI4WcgbiRYx3WkjVKbLGkgF
7PlrBk9C1vZxB3e5BoPOz6yB9nATEkraeWBAdRE76EWZVnBVP8Uqod9RO9F940sIfZOO8/YaXHEr
frCbR7CSIjfDdBL59M614i8Mw8BoO2HCGmFWJRPuabtVbBziV7+KfqGJ2o+nahk9rIW81b8lKPLP
fyS4WBmBkPS1y+5DjXpAFrDmXUTPY0khHaOBhO7HcZAbw0VW05XdeJdfYLEdFJhBdvBbvNLqO1cn
CcJfqf4rtsoSsyreDARANhhTuPBDjbVevRP2LlaqhrFEaIXrev0dzV2tC5BXD5YMT1QHK86tf83Q
TZs41r5JzSPue0OKT613M2eWzr72twRoG2VBwsuJHX+cCmnAFZ4SC0hOOIQZ/rvBOfZIWtkiXeGx
Jsjh1+OdPzjQp7joqmfqJ1yXxkwc1AECKQBqDChDAlO0Llhs0XN5o6jDZIJTzpJ40PIpKtJmmlLO
p8/IF72pwJCh4NG1ApISRhxt1S95UqQ+xamBy0yrcDIMb0+aj5lJJ/cx31mchLTmMGAotGFuPifr
F5DJ1slFOne9HiMgpdcc3AnfD+7zrvO7qZnntSiqmWGNVYiS+N/P13ClHbPVp6xFCwUFFSfD+UIy
gEQIXf35UGhTP7YD0zuMyNg/1t0lYXZXykdoHDxKrqp+3pDSnWpQVIUCc7xAy0yslCnsQk0i9MQN
b5kYf53kRFPZG1pAG5zBI+DcVWDr5KbFqG/CnmOZjxeHGq988uJ2W1K4sPlJphFJqL6qdnCBLceF
xNMFFkoq1QnrLesrhyrvxlqD09ZC7x+smqCgWopWFkTdGIygBlEad1jYvKz//mNkUJTFjQc6VMBt
3mUX2pKQ5PO0pxH/y38dHV5WHloQfGdwm7ERXNYX1E0c2dong+2AbQWkBMTrt/0aABq8XpyqPZnP
2eV5VXJccUfNNVjbRhd6chBcetUbFG8wK1QV0lPnzRFsmvf7UCUptwR8byjsYeGijayOIGO4dm6v
/4Tya6SNiM1TQtPUpt6FEi7dFRcTRnvuOMu4zdf2GU1S2d+9OFs7KrmwZ70t9MIr5Usvi3H/dFYW
McSGnzGLCsynI8ulByYzjr5ULqwmjDOQYGOZ97p9dkn1kRqFbJx5MJ/jKD9RFbUZLvNjIUjF4PSK
2yYlaT+QTciES+VAO+naL9UEGnZ5HRKbwNWf9NGlzkBOtozKNL52TqnqRnhz3fWB+o4f79AKH0WY
qYwniJ8uEbpcxawPdJBiu1LoiERI21RXqpSHEdffrUrbDasHelMAFsXFlbXHnoOEhKpwCdQ6Db3p
9/VXsClHNXcwqMvwAC/yd0p8Gw5lNoxHfFSn5byXG9M7eRXtaLh72oj6PyqyPzKsohIJEUAsbWRM
VGKq+16P/jiGcNCKkmLTmDGX4vVo6bB8cZD0xWfHmBQB3lpEs3Sl/swkPCT46yMbzboGfNytxrHE
f0t70doYCb8X5gdaA+haQDUkK8RUkecCMBFu4tMuNeJB/dc01Tp1EwJmaD716gKKwpu3iyJ5TZON
rwnpPhASD8cPb32Kv7B7STeW30BozlYlKCfcvcRdCahaFnS36x/WYT+g4ouW3SeRf9C/sNLUmb8u
jFHhYNFLnjLgTw3lx1PY1xzexjGCF4fqBGd0mDJCyTVxRCj42MlJN5DmUKEOok5G9+0y7mVObgCF
xB8eFVt6n7xGWoqIsse2HnvhjaqQ3fSogRD7g0dqyrp/fS2lCdLdvrJKahBK/1S1z1bKJ7iVnD4r
VbqL4J4S1GaWKAnA0XGt9FD8VWK8sUoUzGu+G10/6i2uRzyzGCsruVH94sts4ya//niwDm8tUml7
KiSVhYykLuT9yljVprujtknvebB8WB0TVZCyap8a3WhzrDclzVCIQhgX7JIUBx7jsq7KSwvixPz2
/tg9KYc4KLEScNBdqfVljYLFL/F1XzYKPjFarkKK9HJKOCXda0UP/G/i/zQNzvSDDkfdP1dM0Gtx
55R8YLpPqo/UOdwgE0V8BZnyJNtxym2QocMqK4n+BDemjAbFz4XFBKC60fcUqxq1AziOoj+Y57uK
02L4pye5Jp3rmQ8kkCG7CPPISnHvVpyLumpQqdKG7XeE5n/H9vkl061a8vUGn51+klNmsNoVEsAz
y01cGWc8LKUlxopfMUK2UxEBBzlI4XhYJN2/udghYFeFj5qz3IkiHYDw7Q4/EFE9TuTc72wTiOwR
dB9LaVzEweKVQ9UvmsdmWHeRZpt/0Yumz1k7cq6J+ekkhMrBV3l9at/QHZ+Agytod1Zd13FvGnDn
p7sa4jgJt9RH6GwTpAi+PBuTz/AjDp5piSC17gZ5KF8ioh7Bu/ogsPhUpQHkqmEA5WMbMOwp40Hf
YXIG4X2kNL7qlZb20Wx4G0wnWrbJqX8iOhSoaonUQRdRZGm9Y4K3rd3zdljxsF+/UNjomA13XA1A
c/vEvX80FKqaxT83Y0gwVbfiCSd4r4nhxRLN5j4AgdCVSYNYDk6BK0ZRwU/ZNoz33+UkqQ+YOBwk
+0PSpYAxsQUUbCbev5gaHzglCCfQQe73szEuePkhrUeu2Fd5FL/+nk7PoVzTD5jekPXWlSZvfR1i
HmEUra17n71lsHw4euGilUw2mK4/O7IH+BrpdAc3Jyn7WcgVXMCKocaBCrY7/opbEANeXvPW2zCn
0Kx1YRwI8GM844VSl9ptpctM7mkxOkzwQ7Tkvhc6UBh4IJZyrYoBqIiC8hF1h6vcMGJLUQOxLjp5
++y1rE4S9xsOxTAEqW5mDlBtMmGc3zXgFECBJr2unEUs3Uw5j594ybd3HMDFVNuRY4ULclKm9L8j
oMjV/5U3diP3UH5BQaKLRVCOCb4RTDvK5YH2Aov8UBKJ/y2uBHv69cJ5V9kKv4MlMZRFeLLMk8+B
mpaWd4VVxzr3jkjIaaBxEO9aQm/95XrHRdhUGdXxtcre5nCWZfm0dSEtldcad3Rv3rggQk6WJSiP
riYyfyMrJUb+DOhesx9nGgo8EGn+HJ8QVDw+LIcUsZ4fpFRTV8J16DTwic3K40ZwwBQhHv3sy2u1
GZQI0ss709L7lgGLiQbqNy9OFtCGu1uUfjZOd/E/ITnBSz1/mGUgnmUb/gsSUdv9aRr/5muCUIaa
waexOf19WUjlDKCGqeuB/L+EYTEJ9+CKAZxQdc61ECtiNpYxKWBwqvjlwD5qPJ7kQW3A/Gn8EKdX
0S9sVgM4SEXN5AXfRU705I208Fj9xuHUpEknC2qiavX+zYG4v0Mqkz0Ie9UtHcO6uFGXA29WcPvs
D8kSOv4t0D15r3XmC+CMRf9MiPSIBnmkNUerudsldoqQIAdXjOakLaOjq9S7Ri9/IxGZCFuiWG6F
aQiBqmL0itmwPxrmJf5j9FdmJdTfXceLnmK3Q61n7Mn5oDHFhgKu/d0REK1RkAb7za0IXr3WW9a3
zB1P/sFkb95bRgfEtBztY/ohf205n8zsDnwkcxtY2j5QDzYB28zkgtALdIK2H5G8vlkHpVffGPks
eb8GlHjwqEnSBJK/8Zpm/vqItZPXsGiKZqFwPHAjB3OKur7kkbQZyHzxPFb9/7kMP7omVYr7ZnFg
6zhmU4RPg/8rnf8iB6N1Kkcmhx6tyGtpr3OEVwX1jMDJzDah5YJj+Ea0ek8wO1jh4JIMgNd8UFYF
KdZ1gA99Hj+KkTMjo25mHcwcSVBsWpEw7YLzhxJdoy65ZG9MjuHp/uLHm0vJo5ozeaMsYREZw0hC
CD/KZaDZu0l6mLblC/B1MoPkH4x7grIxAyCexFFF9D7OHl2eQ8BEk75NySJjAAE/dIbYLCwmy2iL
VADhVy9ukmykMydfnnzcn23xuAg3i8TB56r0cg5YwQfMdo/in9hM6vp9gd9lnHTDER4oNGEhFyih
iYRRNo6szybVr2cD3O1i6Hu1t9OvnO5bHR5L8gLdaOPKZqhf51cryd0TWk/zNmSnAZqKv3Jaldyj
71cDsDPzlL5mseXrsScYYKUZhG5aDyR8cDRhfsrZXplA+ghdra3Z5w2lQZ8O3/z6TAHa94w9B/3k
ePHGHtRnJNy1sc7XXeFhJ9PlQ70XYJoW9De13Fyu+nV0CRdlQyC8RxGvE9SbaKVvT3m5jMjHru0c
Dcrp6FH0qoE++nLvp4JsI5kJyN/RmJL2R4K+KDPsbicK5g+H9PCckYle6KxWtZbiqtSNL1T3QH9W
Z9ePDlqaN/DDyHahGrU760hUYsNI1rMnLGllBPGc8VL+IS9GlbHB4DhS5WsPpziCu0GPf4K+mN+l
fX8072olHU5elncpi49wn1Fwvb1sIOrKM1i74mCgFjgIUPK6Bzvh89VjYHXP7wa+mROc73Ys7Hie
jGeLUq6lkp6Yyp7Xhxm03KjWdF2UotjqLnTT8raOvfDDq/HAJY5ekmD0zRuIHk1WDR4jFLuzdr3T
y60Yg9VGONwpZjwyZrwZnfUOLf1pts8f3tukPaOfFSXLC75pSoVjlXQ/1H6irCkjrulWBReOyGqf
kPIg72mc8b/OeR2VSXR8XhCGLFR+PM5rBq1aJPslt8cgiJmsL4Oq05U90hMxwuSOrAzu4RyQB0xH
R07vLzuT50xxIFaW8l6i6qK2/xF92FNpQq40Id+Dq0kdrnbNwhoJ4sOAZmxWJSPXfnURr3EtEtvd
LqdjoJkn22oF1XfwU/yuejiT8PxC0thy4U2rzNG78pC5C3Z2GrEsUBjD9LiRC9Tk+d83OymxGo3z
y7CDc8mMitq+S1W26JlskWhcOwBfss0gz+irPyE1gFyE9mEb+bWMkxvvEqTy5rIpU8vwuBx+tMps
11YOVKS5H9Co8gtSAC8Iapu4tc/kU3xe+pYabgcVUN5MKGIZHOL6qiUVYjh1grsy9gIkA9Q5rW4N
Ype4B19GybBxKaGS1gNtaAKiQt1USpGtCAQMUYRhsXj3HMpqqavUuyqCdDjK2SfPNG7JOc0J66Zm
eEhReFcXoQvg74nDPDwcRurYwYwBk+dMffzfYVaPOiJ2ZB9hITNIcawqcU/qtSd1vzsTlwuG+Iwg
H9KK9RYP6NR5Rm9IALzR5hQGAK0AKAtFVfEvyCBSMd7t1xTcG2JZlLNL7A8UuluvHGVNT2J9V+fM
9NvdBH7XjudjLhWXJQdwMbzotwQ7VXu/yCT6qG9n7r5r+EqtVWrPbOnfgt073xCdFjIA35yyLTjj
sV4iM0eXzrlzo/9sNMUWKdU1otA2G8m9cwkeZTcNkDMEn7/YNouzsXgCKq0Kzd+XM5SxD2uZiPvb
ltFX5tLl/4mxVHXxKN/lVmfb6qYIbsxu5ZoMInZXGDd/XTkQTdmmXPbBr59aQEoTb2cELDPVRuQ0
ruXxciLvaF6x/HyqJ51uPRlD14UyUR0fqElQToq2KwTSfa/1Gq5/Uo1pAAlIQyZs/IFJLo7990Ry
u/W0meZmIjSmYSkOhM5VhVq2/rFAVx7CBnQM3HZlGYebLy+uvSoUNP35dVBqLGSR3ZWBTE1mWdCw
spWUpOBL4Cu79CngGHGn5qBA8ipuLzNr5r4DQWzKxbSmwNi0KQ4PJkOjNkSPnvpIHWzj9/9UVbl9
75QLa3SG4IxrStUSwnwNRglHHmbI47NUF7dop6h8D35yhkBGPvrJ+Npce5QbUKwssX3g9gnPL2lB
eXfzEx0TQD/nkf8z11UdfrI6A02srNFrX7INxyW1OLd7d0cJyCThTGBR91QHe1yH1zww56MRts0h
dh6gpAhXgG99q/qSYa3ixEvNEZm54hGEKZspd6vVPsqZKShroQEdSHxHcYObPuC1q+pVgro6GD9l
KTpIKq3aX+IJqhHqq8HIE5S/m0b/G5wQEcnehS4WQtxguBoYXQXjAWC7YlTAHRiIpy6zsNqT6Jgf
8RjXsIs6QsFxzDF9GBmEr//gW5KRc8e40rplPyX4Ryu0380MLA5FdEZi8sjyunVTDISGVuKnU3jP
o7OTm9QsThMT05Ubo6XzFp7H5LYLKx3vL7boNstCMjbId8L15LyApYmEXTEAVNPzN2YRfoNu8+yA
YDmaBQVWw6HGOa9VZxe98PtyQ1Bqjxc/h+Zm1a0h8N8y1pRcl9IMKWhgXenAnU5dVxID4WIXbBie
6TkDBEtA8nezeFT/LVFrPLrWWt+F0lTctWo9npc6vnKgKO/53WnUUxQnav+i7BKrRZzDttfJ5w9B
DXVd/Rqn0gWzx8Ah8YuWHBxgX3k9P7PZogEUJGdOMENlrsZfiORO1LNes6QZ6m3jB/FV6GEfsYE7
trE8zjkv9y9FqhljN/tNPYGlmeG8DE45K3CAZAl8g7a+jSN3qbAUJSOMmuRK9d5bskisreFHCL4b
kHLg/himf3otsUMQTelel/wJXFMqP+BGL54ZnRI5VBzjtANxCpvIDeQYRBwD9+W4GhtSzLuDABDb
y6ugFKGRKSLt1b97cp0/zrAZS/pqkEryZ3YvsnC58tyfW5/+tRvvBmnW40o4PV8nHh4jjG3Yxomb
v6VS3srLqsdV/b3xJsXD+vqQmgmRX9w9hjiEWj/WSBSCkWc25c7P846SAp6PK9FJSizBONxJ67ic
t2TUoOW6RP6B4leunXWVORgKz+hN0bk0akphQHgzRWrUmZXoalkhyOeBmnlIgVlUk3qdHZUlu23v
F3I7lDX+ojne8ssKQCdVXOVd2TJSiNccXgAb/CzWJ/xMJsuA8xemR73TGuqyxdc5z0KkSqng2PZG
ZvONyB161N/44L71tyRkeZVLHGnMcUPTBVSRgwHpcw1z/fntH+1ake04uqwfxUoM+nI8y6DSZ6I9
KbHl4xnCRXM8I2AxwBLvCAdkY54v+cyhRezGxalldtoECMJo7w7XG72R4a06D4OvopG/zCYi2QxF
7TS1IkgEwh2RgkctVm9jj0K3pxBVw+MRANdOunmJpk6kWXp3BKum/xDKMrePHoeFE0w+QJZS0otI
MtiPFppX2r8whGDF9fyue77j4NB5MQe8Z1rWP++V92UMBqeAdcq/V08kw1acBnn83aPnfJUqVUzy
HJWsDJN4Gb8MyR1nXoiQ9S6obWySNayYp7PXO3bAmlUCxeVKNe0kKQf+GGcUa7Q/YbVsj098cwU2
QRwOR9yK1lz+hoydHHUAIdedOGeHaUGle35JIlnWPiobJBmPpAq+48C7bn/CCWAb6ITcQEHqzGG2
+cm0qWwWEStZ5IwJThBueG5TlNoJxIcfstDWtBocwdBy+HqBh6v2hmFQpP+OCGHYXlSE2S/x4byD
u0gLibI691kWbeHl6w6VZmhhikBSOTTzoKjuH1XEBxqC+YJbkKJWY+dEhinhtGIzO2bNLWLo3+Jo
yzZUOSo+G5SD8yuOmz05ep1rv5GeWGYle3oNOacYrF+ZQL8QW/kLVqnTcunxNoTa+VnYviYLA7lN
SFw+r3z/nraRYshterw/TtlFY/a7CcNzX40AA56AX0of7Yhb3UHAe+SiWNettF6mEcs+P8A4KTnv
uvtOlbH9w7jm0nOtjWBQU9Q77QlT8hFF02D+4Q2o0OoR4TvdyIgaDd2TSW21RV+/fF3T5zSGBLYh
dZowi4KDd935381tCYhqw3tS1uxW2+kxR4F+bDxP7Z9+aPA6tKmUFq7SMVOVGqc8pg5VpKqI2vI8
UnJGNv6xTe9oitiqQwWtMAand8c6J7cPTBrnum4CIe0d9W43x7l2a7H2hFwtjZihh/ur59Mk3b5p
ELrtU93cS6KePcAtWZl7IDMSHGPPjvLHyIlbji+SqAHfltkRM6G+qomysHhTBD5o80ok8+EwrIIS
JjVRb2IiJxD7Wus+euiac1NUEekud3vJMGnhS/efBkxB66HQIkUO8XyyvgmQ7ORRDMhjWZrf9Eyt
46Fhcj/WnptcX2Ff+rU3mWBFIK8Hr0Da4PWkhPzBA+ZFrmb1mSXmPD563xUC8y9tGKBcfYoxn0QJ
7OOKVs1RbKJBciOAk5OcUnVSiL6ygXelBBC/q79hKOyKbqLP0TV59W8MM5qrrgom/bwBs7kQr3Mr
vCvq+Wm3wMfB8VbbtKw7N/EtiMJONJAhxKQERkQ/L0MmZZZYo/IjU2dWd4HQI3/KbVhF4OJRTW8C
ktZenpwf55ogmy3p1B9wTULm/SCQXQDVFuIl2cawQ6zlOvsnRNJMSXS2KFhjexjQsGkr2jCikZnj
igzMBweiHfCbFxbqPhdiZMixeI34ILm4zEHsP66Z4SqDslhCmvM2QgWzDI3geZFSCm8LOqoByygo
rQuJbn+d0daV7LiIFb/mQMkqNyXKcniaqLOLCxv5noDneur5cVFFPGXVio/br8tOA9um72GBu3Mn
Elql74kj5CvXysoGYqKkfwKBp6ynMjKXtEi2Kfbta0rPE7wW4LwRjgSC6R8s4fI7EXh37nBD1i5f
Y3ajQIntc6GdQBSaE2gmYQKvHwse4uPzdsgDy2Om1XCNHdBjD5Ab4idk5B338rzLnx0jVEbFTDBw
MZ0cxdR5unRcurTzmVAQSjVErfB5tnYBmJahl106/QYTJOiM3kjIUX8Z03ndH/aeWMGS9i+Q2b0m
28d909OS4GNJcq12IfWwgij8kP5V+31DLBZGbOFMahRmYbJ3Mp4b21QfD6iRKbfJ09+BOF74mNFl
wzooxjcTwjtofU80ulZUPw6Ju+Tn9HUulyL8OWQvbNGIDzAPFZLFIP5ruVY3sJLYkfEJ6tWjENPc
YJ3T5FRWvLegJ2+3fkKugirJrsBlXlaB0naQ/GGHsHWDBTN5FuGJJCM4J2/j6QbOk/1yw9Gm9YKU
shQFSbQ8P7ZISJYxSL+D9YFW9xzjlu563MdCjwtCqYFj/1G2mB59pap6ujkcW4cr1jhGx9CYTDJb
af1jGAnhlpCPdQMdiwjvrICuLiW00unb19gCXDTTjWJ1TKXPzxQJ/GO1QD1N2nq5y9IANSlDx70m
RNwekNWECSj4nMsqKNEmbUdN7tHJFRd/VEZssVfgJjfNTzqtEnorpQxpPOYoG0f/QTLUqd66tn95
EJoT+YmnqfC5sGl0joTszCx6xYSIbCWXGVuW24zrGOW+3tLfd3ZwwL+WjalJeou8n2jnBZ7Dnun1
quSv+Ie3YgHrpfX6Z2f8m894hC1eX3pozESv6j+fu1J4upkUvhVFuoAFgwkWStL+LDjKDCBottGk
5dsB7BpM55+GCGT7bJ/+asQBU+V4687r5pLYanyXMiB9m7wVXl0ZU0d+o1i+/OnTnGK2PwvLrpA8
vevAILLri9GVIpjA8NzIoUsZAtgt1ZaW/VG0pH1uixzlQjOJeFaCO+jMQLc1+9KfS1KkuusPCZfQ
ZBAs9zRrhZHNmfiwE+FSCCTELefVypmopJPfje0KhIUSM3ReqIobpzLegHVlTEZ8aIa9Ma/mVXuI
yn5tnDv70t77OoE51QBhnFGXdN4wYhwtUjsnIRAPShXMkLld+mQbNzLwjMVHCqxjMQkk+zv5excI
Xinp5SuUEEGXp7e6YL86bziM5n9iA5fIFY2dgfw3wDrs25C302+tOjURHqEmc+yHqH3hLkVQiVPQ
01BeVv8SzOE7eK00OL7T1IgP2ezlRw3+2gMys7yjaj5KQKMKshZIiEglmFAkUqDC48D+sdx0S8OT
0yunAQvH261k9dNbI+k9DOu/FsCt+B+SzzvGNBGlqlVa9sNXWZgIFpYkCLSxQv2cD9mKR/UL5E3j
k3QZuTwQR2E90pdWJdH8MnGWSqtfXdKA/C7cWK+Py4qfCqSRioupy2N6P+9H+//JNd+lYJZTUSnU
1BYOF6aRnTYJ0r2guq7Wo8EpuqElF/nswAtB5W7Nlp7E1jyIisZ1PNzIb56u1cRm8RkzvoLJKatY
US4B9V8Yys1ilE4QY18F6Qfh2XPTK9zBFpWzBebuR6C0tbrf0ASgOx8jULdQvNyn9wFfzHokb1/h
0uLkbRjzDtnuq+T++r09BkpSUQLL6gJmX/yE+gn3aRd+clh0MvSfW0XQ7Y/9h/kF8DXA0CBs9Ec0
aP2TcOlM91VMZF5HghyBcu8rffKUW+X9TE8qFYeu6uh4CIpZKRKLOvYey9acnNwHRxMlen3KQCXv
3vCkpc9fz5/fuPNVhXDydriQzaDQiy3GRwKaf7QwWoRZ2nUmjWgZcMMo4hNNu+gbNHKsLmb7u1Yj
1T+RAHereob4lbWxQOBx63XwMHnebgp2s2Fr6nCfOhkEiLncUA52nbGp5YiH1HIN0HEmfI0eIhWj
Mq4Y74bF1TGuXywDz1XXdZer9asBJSTP8fNlNeZqHqyp7QuSGGvw4IS5VFyzYBYfZBXzW8l/5AK7
QysG1nMkzHVAOswlLxwReZImAmLWc413jKh8xr3I6kCJLXC4R/cDvy8ysfmeWf7l7wIbqeEK5+aj
UulxuTSKwhG45yQnaq3ZpbRTZZw5LLGLktqGRYXS7Gu8aWIkwccPAKxYPA0SSwbMpVH/HUt99Bj0
vsEG/kwaB0Ts/1onJ3jdgcymKFQdNwQ+YVstIeS8vK83r31284Adn9my1L0Caq7xYmcq6061uer4
vXpCm5TZlkRF+xswaOsD1MUvmQLabXkqSxHomw4HiUhnLFgbZNEiZabQmH1RA6l9LEq6sgioA3+R
zWyjGdSkh+ijM761sC3daWWjiTeIvqxnslFjsa0Vduq9RQbQTHNbagWBzxKjIkVTeky5r5CE0Doj
oK4muQ93JOvfhHlrW12d7bv/PtgyTr5ILwK9IiJSpveZgs+urkuEfkA5uRFeDVQxn2Qr6oIl+izY
IL9Ldxkziek3ayGp1ynQH2/j2CdqN01gK0kbwsi3yNakxqxlgKwV/nT4EV0BHp3bQ3ZVxMNgMMCg
7hNfZHtScrynL/XLbezcsEuF5U5xhkKb1u+pxy05u245pBiI/jCHIAuFvWps2GWWqcb+vc+14/0H
/OiSKEjifQtEvXm9ac1aNlYyJW3f5L5Gwy2aFRh8JLFj5hplVuAQBHIbCKXXXqkex31l/G/F9YeK
5X1QOjYYixyu3EOmOABm87jJVOowbZB5JHhP1YXxptmVje42fV3UjWb+O2QBm0CWfznMYcQpuC6F
e7oTOslMFsfDWtcRwWdLn91KGE50s4hhUoDJuqq0pF30rxVtoYbBjOIsOcQf1/29ytmaqZ4EJLSc
4jvW7rVFVUyRzVnyCPvkfY5wfVpYd+c/PFaH2mo2jI5jQhs1DEEwEtlwMZHLH2EpvhEEXrHJ1fD3
VxKr/dvvTbiS51XniymfCsAn0udRKCKE9PSFfPVpZB+si+Vxa2Gg8dDe5/Vfs5kHTyHXQ2Vx3Ygv
ibeB0tmVj/+7sXW6U6Ufx6oepRTz/3TpzJguDAo0UONb6656M/AYgYuCvvUvOMEbLLd6Zx/joo5r
i7Nu6ahxZRLjcicrTTotxDzNMwM6I4E6JsgCH/KTsLB96faOpAGiKwCjPKuk1ekeHQBN9L6RgcMP
7yCvpREoz3b91a4J5zD6/nA3dtU+en8VusW6j5GsDsMo3t5FP9nDpDxRSXFp2DmBlD0h1iN5Za4L
ArNucTKt9LfqQumXClkvOnHw+0VFjmeB/1H/u4foe0EZcgSTwoabKbrAAGqxA9SHvLWXO46v/rpM
fe+TEUj141cZL/dQr1nuzw3Zdn+l1wKJfPpDtGB2l2skKbJ2OgsLZARJw8JntnKhxmffDZU/zZJP
X/WgA9ihRcfJtHw+Y8VwpooUbsVP1z+0AkJvE78TKA3Vz8Oc9SuzOBE8oogs5x366eNwR306Bg/D
pCIFtXlrYBPX04k0AQEab4+vWJWeu8vJ6Cr2fR+8NC1MiuwN3bE2oqvkH7i3nQyuBh9cq41TIPau
Qp/jfIIZ0VYcduzvTj5AQ7asF2KCJJAW5XJehOPnwynFTsSMOD0VvuvHdWPMXbKvBGz+TL017/sw
bWWNroJml8QXniXmj7zQDajYs+RUAmNvMJZPgMf21fZP8jkc25YfLWDG3GCHiAONIpl30Lrk6nHE
6ZaOWY+8XE4K2khEyHGoLLQyQzjl7GP7WWesYOeCETkewBsWu3+GT/opUOMuobL0+8ZP807/DRll
z0dKAlm+lEzzpQaXDMpxTfKyBTyfOLzlZ7a56DiSl4LKtzVlE1m0h82rqyQY9KIvu+N4ZG2qnXFS
HE1p21sYWFfOfkc08Q9YduxqTeTHfYMPEfJEGkdPw2FDoK7AkE5p1xn9eF+7Fvt7nYAVn5Uxr7/T
MrkarKpCprZmKZSbFo6sna04oJm7lbiT00bCIpJIAtMO0c9Ru+5MpmnKfUvRIRRoaV5alb6YXRNW
bD9DvYBu4yQoi31qQC10fFkJF1AjoW6bRE4p0eissdGHZbVIxV78hq0dOgBSR1SLCu3bkdrJ6wl4
qEUukwOInKvAp5848wczht7DvDNaDGJX5rI3lPPT2PmoCtjzarSKYgDq/b0ki7BM4HPPeUJR7zlc
EewtY0GhxTOaayIx4KQBsCyHj9kFNd3kHVayOu2CuGcOc+2CdsLVCDGXUBef49G4at8Wq90qVNPA
U44k1BwDhQmZLWyXFJV4X4uqA4+6+kr1iNDmpqyvFL2Lgvd4aullmUXJhgC6VhKADu1bXppBjbwX
7gQDLYU/A0U6oCfTc8YgYH7RAj95JExIENTWTVOY7Ezl8bKX366ADWFoOHLzkPBqi4lXt9f5xKTx
G3CsQK9vZ/Yi5ZBkVGZO4Qgb+jC7O1YlOrHcV0ieJ8brOpoYPDyy8B7+pwmgpAp38b5aLnU7NQmr
GvAs53uKP0xTlJO1IkrrbmwDwzhJ7GRWI/C5h+qgMDR6ZOsOt+NvpnvZeIy6Sxls/9KeS8+/XVJE
CtaGsdUONU7lalF5FWNViI3Gqfc38HzWXM/IDN90kq7xUMm7pZpDwW1fLZkrRjXfeyZfH7n8k/yc
VYz+sm8kAx4xxCEkDFqQElG6qFbDvgsc9sgg4rA9zuX2VbAbvRo1FjmQ3C21NTSLRm/9tOBqSJWG
lq4QPSX3/52ogIPHqMJsu3mMRgQ0VZZkleCzvsw50OZVk0bZbyFa3hQUMPt+K1Ggi5QSq0OazxyS
EahVrOV0pDYjFvpAFCCOnXX2s+4zjiLpvHd9wWKwrLXok/HQAeuZSse1utWi6Y3nIG0r4cM9KCvm
eSrTizWCOFqSIA3QbDOWAybdiQfjrqATLCoUr+LAAOGaNfYrNIDy7RpYhcJZAEyQWR66j98aphgE
3Iwtq9FbDgrOYN6n26V8KRH3UbFiOE3Exxuzj3s3n//GyMy1gQhhyq/cpex4QsH7qosEkoEoh2Lp
n6Tuw7V//A7JabTFcAiSlOhdsFVu2eFolcfEp459UHBwKEHqoLsTU0T6b6+Mx54daiE2TIClSZvB
dW98Dqjlob4N7T8naSWOJ1/XcdjJCumgWBAodDhqnTw6oCgWj5k2FobH13LUwWbD9ZRV2ARzN7HI
Yhggo0xfEpENIWzbnRVf94vbDwwWbgsko9XvEtTmqcwtFU4ewcyt+i7Uk3+yc811qG4IvXDsBOUP
cYOO9oEn+mn9xt5OMS96/kclYzA6J0S3t26BG9PiZdz9O8Wf91jKd6GEMO/XmDklp6+wW1Vet6VV
HvHO7HkaiZa4orq4ywd62Yd0r6scUlaBS0V2SfQ9jibh5SoxLYNpH12EEjV3HbT8EE5BoQIvV5ni
njjnboXi/kZlOP1iO0das1BeSxCNLeSy2qRgIIdsNYILvzVE7phi+55Y7Be9PPUIUFHoha4/RiYs
aEZWauaTJgXeC4oXjViqoAQ5ZiHKGmmM6VyU3RMBNpV09RbPTxc3Hkr8QM8EEeI77ahDWNF81PNu
TCnNzHyCBOwx6AiGKgsAMPktBVxxNfb7QMzGMW2sBaiN9x5+PEye4EzOXSm1VekhbUgHy6YbiUR9
+ovIvjTs0Pdqymr6oZFuPpDKCLCJLe16Ze/EquQSSjTB9wlEBLKvZ40GI7tDt8Lr9waI8wC1tayO
cXSXN4a5K/Jq/yQL8sF0c29nV8+tgKSxbo+YyPd7r6XeSnQr2V6VC/83jx+Qj4xiIf7jjg6YgrVG
rmK/C/Vzb3VArZkJJux+s3mSCnXxA4iNro1fpzWould833KkYrVbUCkYkhMFWH5NNpf4aDZL7B5l
bo2gF4ddq7gbcDWgs3xUmpvy5dmZd7HrCsaGH9ydOVZNTjOSlDFWP2BS3bDCKJlcHMUNuzanFgF2
lr2K0FqAUCYK8KQ4YjsUEPL+aS3+iFPXyNjlNww796iFzvOghIbHVrwpzkhswxEHH4c8X6mgclfo
mOReM7Pq+NOWJxMY9k9kiWA+WQ6D/VWlL2QiKk9E5qwhk4NM/kpYLJm78aex5gvwJQ2WCVVBJkAM
GL+lE/6ifAEa5ftf+lQ8klTByfyLb3pr/DDxOlzbeARgPfpY2Sjbp/p2x2ZcapR50Ghc5S+zzp9s
X/hEMhOea1ptGOFX5jaeRltVy86kTqxy14rUzx/Q0kFeDRlnQ79yWtrrddjcDJOK46hrxY4ucgXy
GtZiiKEUDRBECCYGJ7nZXnqtyXZL5EMuzhNuJY/hedztDTegWi+nK2gczI/3bO2YTYmJiLceTgG5
j7hf1EYT2w/50TS3ikRSohVZgLkz5y/VYWWwwFSgqg4kAutZs3Fb6gqpwFatRHX/tdTJsjGs2sOu
BWhrA2Uh2pnafORN5oBmvAwfQuKvlEXSnCRlM1IKaf8y261i1m0vN6ycH10p72VHwnrhgFSdAjZr
sbMSWyHMbEIYC4P3LzC3zBKO9d4UEiKgvWW4DXEdwkSpmHa47yYgMaJEpeTgbWpslEYUgzxlloCk
I+e88Rwqex+i16TDyBjq4yA0YRyTH0Qn83azsUfJTLwSCMoJ/m3ZysjC39oVr/uJ4AGpgoDiDjDL
h4MPlRaZ1lXFekh66IR49aDnaB15PE6G3hqqdq0zU+uGbq5mf+rWNRgzyi+nbGT1za+fc6shP6OM
bDGUYEGdUy+QEZYMqOgnG1W7+cDMuKBX4y+lhQY5744tT5MuHNApE14lIZZArt69qfIf8qduMyR3
XAp+BZnp/4sfOY+UzJ1UQrXAcSN5kqaedy8dCBGUZW+8ExnL2Pv6VVTtU2Am8d6nH0u8TJbt/hxa
XLsATKp6EwrqjrMSaECOO0M18EbRlPJOn/tUOgv/tSJEkn0kxaXIK1EfyW4vwAI1IA7QXoV7E0fF
D7AVP6/Wx0n9qwur47ociQkG3FZKhoKDOQZzlB+4PIpPbHEYXnq0W5mrsYc9J/5isMdG5oMkfJjC
+bNTg97TSIEd7y26kDBk8ygFSxlKSOcOOXtQbC5jK/RemZGWISWlPC3re+gZo0wv6D7sdIx1Wnf5
YOC5DQJpTNOWni+8d+Vei53fgbf2AUK1wGGNwyLMyMOwPAos8GKWpe5FK51y12m9dYUgbYzo3RVH
tfnvDfS+jlfLNMRoKcdWdyPqpWDU5/5Y/ynDA1N701THfSqYiWXzzBcJPujprxaQCv5By9mxPuH/
oLQeIP5fHjYcdJ6PwOfEvL9e260Dc3Yuz21Ng6LmhCZtOUikcnd9qpCcX3GTsaJ7TL/oJ3Q32lB0
eV+HaLyk6qrrRRgx8F36tf4sgl0rpIZd63GRjILffuydjq2P37rC6chcwqA8/zRaaDUKaRHf7T5d
7UdM11NYNSS+xZVDi80/9JX1ldP6bhHW4h7qAcSR/sO3etY9CDKalkQZVWwjCgj5X4LOctC7Etky
hKZbqRRt8mY9xzaj+/dYQzcHmogf+mi8XrQAvMj2kux340+2JoAzK/GSLjYnvKlhhn1jQHrw6jSO
+sgnWk58GaMnSqFW/4aAQdV3+xnEcyonmUHe9LNBIvr3dkPDwJOKNpSKuHENmbSL67DBk4FLNR0A
RnQrJW6Cq21mhr3k6MPdZClquahqQIgSItSqJXqP3js/t7HWdIyMRRcspOzxD/PZG0Kh513ThDjF
4RcVgJVCn+0Kqo+9e330VuoXrBkWlNc67j/yec0rkRGm1Io6u1y03rdB4YKT0rtbDzJwbcoJI840
bXFBdS9kKNNzH5du6I3uOnlIXhwEjtZMNJT1DmNP8Jjr2uJ25lyQ/lxMrFrXa/SFJZx3SkgmHHx1
6SuRakeNYYvvEqjQ+MzDKfEEwfsxVw5hmCrozCRsUEGqzxYv8+if0C/3FLH2WsHRuUubHwrGX8uu
48r/qLEdPNUuGcn34UbkDodyPzqHKHpO2mytKOADi/1zYGbHOLNF7mhSTOkXdz/8Ssh7fmCYl+vh
jB6Fn/l6nRPdMdBstR21x+Kun6+xOtqCexQMoYJed1t6ebec2KxOEZBpzs7TnoDCo+UKZ6mrT+O5
BipW9nic70U9V4q1BWW5fCGgbhKH/cblgE74Cf5ItXfxQy9SmmXMvZ/z6EuSi6FY037tA8InKQNV
Bl/c2mFaXWA35JAzDWHxjXtbKgBsKB1QPDqsRJmzAfbNH/YND6v9751dDS79dnMoAS+Mu58NIKZ2
gXkSCvYfTWbteH5F+lUBJ0y6vs5VJU5XlYEdvvG9zYbHN+jloz4326k0SAA+LEABdiLje+J2OtHh
qBjNp0I6mYDX4PkSDmimFDdqOL0h26uTicWxajufJbpKafBHszYwtq8wyWIGM0+4c3a1NN4iNg4k
VdOUtDZoBIfZQqnJg7mjKf059FIzeIQyZ/51uB93gsDWI/+Vl1wrcbQTD7DajwZklq6NU8rHA2Q4
zfymsgo6DarNSYaUjpl7WN1QV0v6f8Bb/HTuDBFK3+0lRlx4vQzhKq97zyugP/nSlQRxB7dnuVMT
RodOP4RQqfGaMD8Q0j7+gALmI+m4My/CtIvpI1+FDSZ5gubowaialdYBnE8TsOJ9d0FAqhxu5OMW
gwVovH1oNV9vG6LPMV7Rh0JdD39Q+3+EQ5Qsb/WLTyYZBCkSrgNCSQ7MN/7wJaw/PpyZkZEaNkZ6
Ezcf3y+InjGQYb4odfgBYFmSEVwADer5sRm6JYhLkVl8V4HN7WYrttFeg+Kl5qdaMMbIAPFTOfNt
TqtTWXQNyPOrR4iFM0iKDfeHcNCPxgIXM2GxocJcRexTiMcvhvnz9YZS+XmPY/0OIQajq9U4P6tm
Oj88wbdYIyxzXwin5g0FUsYolGNXbFIYPrO2bcfzkR7WHOpKIMIFPFQLep4f7os20OOXU52R6Axw
QotOSko1dIXiArDGpN5/7SEj75LsVnUBJJOJsebBcWWR8hFtESMsr6pi0DvF4QOlcT3dL1OtgSOK
qMYlM0ys02YOmLe74qjCNfdezzcskMYslZfmfHMj6Yo7wCni8j2LjrTuSiGxwJGnlYK8ppSPRNE7
iZV4v9fIhTqWqY40xRxUlXjiKr/f7VPLuMephjj6CW6U+9o/MYBvdMdTg+zSixhkoWoVVilvGBMF
ajsQpHcVkBPomxNzwNmYS9XCo4ZsBBV+8ZrMS3+dUTBvS04eYuc9Zi0C+bZPkMePYiIltN7Lwy4w
ukKwpqxcr1q/SWdKjOrN7Zc81Wf4e5Vl7zpKKgzEwp7SkIZa3eIK93980ZMj2qhyj8vggRib8Jq6
l6hWg1eHLWX2ELB+6cj+OfyfuHmDFYEgcxFtNUX0TYkV6VNuv+5A6KetsqFHeOeG2LwFkT2aEYCt
8qtoIkjN5GAzRR6/2bOwLopwIbyy5rnGbh7ezigEdSQKotBhvGzyeio0EX9Rjm6ixeLFm67IV45P
HSvLiEnmJT8YbOHeFxzDlvXe+8os+jqIepaZ5WZ9Wkhio57U9+9NKHlOKtpGWAwq1QteECkWlrdw
eD1m13VP86w9BC3Eg7T18vy2OjylG5oSHwjtmywPwKOhgpHXVnDKjQ+WW1hz7xUW577x7dV5gdzd
K8akzzRjJqA+CthDoWaZqjvLd74giIS6FEu5r9oMdAbY26m9QkaSAZibsV2dfmhms/GA9j+mbiUc
117exxPmmiPB68v2Oi9rUqG8SuvUiK+8m1AixW6UWJlycf9q3AY9ZxzEeaR1XWs731FKySQs4V2G
KoQNX1CYZKClmly98oW1xPuZVEt4MPhljRhw9YiJaUYlXN1hItKgd2xDpTfrr7GUalgk81Sy7UvW
Q5UIvwPJzTluFD6Jaar5uZIa7zBuVP/p4erKGHmzeedZ36h2Sb6XCMNOBoxykykWtnYNXZMna5Zl
b83fDIhDVJP2p5jEdyXF3VzKK1Bx26YxrmOR8C7cjt+k+s2uKI6ICeKRCobFVz5oZHuiUzjPknyX
2U5SBeBP4VPaK7xyuyP7IWUEQsG7N36kpPQV2fFG+PNB1iQNV2etk9BSEdiuuJ6WMZaoUPXxbz9W
MQBQxHi+QWcMxg8ZIW+NJuge63uO79M8sv+0lkTjVHs6i9HoSF3HnSADZG1HI5Vl6n69UXMEgai4
AQ7icOqZKWPDlAoQAtnmXarm27vwI36AZ/iJAcWYlj6Z9akSZjtOHiX1QIXoG6TlhBzOj+Krofhh
m6dK1SyS8e9BzwgUd68a4Y0Oc8y3orpL+3QD2ln9O+zqlWsKr1ALiwwUdHl6sW+y5i0AuzgvDyYR
TnTp07jZDiIsyKtHpoB8y3OjcZN+XGdjIoSE71rXSsIdKsArs6hGz6cXgJB7XF3oNkNoGTAEIPtP
wOTkVAlocuPLCDUwer5wdWcEILHIrhlUrMHW0RVpwDMQFwDW0RdgEJy/ajQQHjV8MNXqADCshq4q
Bj52DYza3faIIPIv8M+CmHRCmfX1DiWscHNtoBp8Q2oxO2zbePPt/Z7exBeSqc99uR/kdOtpyyxW
rbyiJiivYL23yYoV73UhhE3xhG4C4vnwoWYySJpUwQSaiMHiMBWjkenCY3fsJD8YT+AapFssJr7G
qdbvirpQvTMYot+wHvBeRBeft25d/mlnkwXt0Ta9oaojWOe+fFRB7GmDbc/Z+vz3ggS0CaLyxmuA
3f+M+fmKoyw30RBiS4j0ypxNhK2sFswLMtmOnOaw6F+D2zguyfv01teJA9XD+1zk2HFy4RTZLEVH
cuBJ2hbZDe2Ax9iylwhKLijvVNlLS+4Mw9mgJpYmQxelnvCgoAQ48la0ty2Tg+mHNWjRV5URTKCV
1T82GYqmf/rn6gb/z4UW8WQg3Pihh03lvng0+Ec4BVL1+jszUCy9BKuNxke/ryh9epCTDXRbKFse
qLYScg0elBQUs0LfZBTzfhAh+NH8irZCRUy1COYE9eLIg83l907JBX7yoICyLnCeMWsIU/zNQYGN
WEGbPiGpBwq8TOH/CuDGRY84RqY3gOKJY2W4SFVT8X74cmCqWf1b32MEE5AJ3Re9Ei5+SzLGN4oI
/OmRqg9NVxIst9g6r2BIvoMquQcDolEUdh3eFd8imv27/jPNWTiJZ1iczo2HA5g5sPuGhEVAk0F1
ll0wQvCMoj7SEEwLDRdtEN21gW04kG0Yuo50/IPN5Vf2QEfSEsYyIABeDwEkMWv9REHuWIlZCM2J
w3p3WncmX+qsqMjr1tnfmr/ft/1CAXh1Lfq2o9eNjwyrc6NRfBA53AMA6No28UKSaMvu0o1+fK58
Z1ev1NeYrDboqgXzZsF7qK4RH8Y9FQHriPrcgVsBwV2afwF/HHZK1EtjyGYSqMXADTU0k775SPV0
MZjocTe3TasD81ZcOJOwJzm8GTSLsRud56rtVpsmIm/OCBnQGg0nLQhBQyQNH/+5R81pXLq5GPW8
ZvnigHxJhyY7oiViunQLkO1Zx7+y298l/Ngm7c4/XgFWhNXy8E+AX9VpvBJpdk7VS8R/iA/zqQQa
CIRhN7ect07UZFnnfiquT2jWmLhgfzq5che4SPdNKIdkaVHtugFRs1jdRBlY0BpaVhmSEJhXvB8F
7CkLsePFjvp0AsQfiaksg/10KWr6fW2LsCecaTIxMGg/ChyjEQrtS9CfrqbGpzCRYWgXUEwrfXM6
CwAL/z4ZiH6/2gDjyTia2FsOROEkSq0m/ycljOp0N4FXsjTXfnQ/jtc9TyG4gE0eSRxzyN3Y3f8z
c2Fe+kv1xrtc/OOqT9rQpaZrdRK0RRLej7EGhhoymJ1tKgpYrQJf4dU4zaENodmhj4R3EJtHd7IV
jG336j3Pxn8gcD+DQoTxkIYj0bZXpnRNrNn2BPOgTAh/Z5NAzLb7bThnBqhXO6WE8v/XAaH7Dq3x
In+4c3AIjX2z5eOjPeqUTsrFGVz/zT9Rg/fqk2vBlW93F2Gzp+qTQT/Yefi2ykhZSIU9j2qF3jFj
pxFI/Pe6E/80lngJfGobGBZzpJpNM8PzREMeRpSHFUKUkHvqVr3LLsx3j/cQKscHdyuiZgcGq/Py
bE2QVyUh/yw0TvalU1T+wr8/T0VC5Ddy2LqITg8MWnotbTtgo1ed4ZL+oNBmaD4x0klft228J1XX
X1GaXKzL+3nwIf8OBwams8DTMGIsqZb7ga2u8nBxDpGrquWpfD5m4831kOVTWs9W0iNOBmZzbZ//
LI0AaX38w9611flExiHuxJ69Z6B1CBj2Iiw/CJHQQWYsJFK6nDurwVnBJGrnAODcjLtxNH76wojy
qcJrSlt7IZL0Ud5406/j4Y2sYZB4cHfCoCxVuPz5iMoFMtfkSBGByI3CODVnWZ/mi3PKlbHvys8a
tvgZVratyAEY1mddPsbCL0c3hF+G0nhjDeh7yCSJWK5acmqMAnzXnawcGbqf3lBKbxtf9FbH6hp3
WQJI+oCeJAjONCIGZuvll12A536gv91UNesrtYxJ0aEMzQABlNxZTRD9FssPQuILnX5nnRbiZ+l5
MWkVaBwuTPa1FOa8t7F9NTfExQV030Hx0BEvZzl+CmQPlrmXfp99rsAD8hsrlESEME0kNfQZtErD
l3qX2BmhD9pl0fJq9LXedn+/Qd27iP7AsWSWSpwrRz4ENPjlc/Ks4iQE1E8+AaOIthQEnFNHsTH5
p/S6gnO/wE4ECV2kQ1jI8f185Ll7oCCHK8QPoF0lYIOh0BXMrd4QuaEYIe4S7CHuc8D6q3oT/9nm
lnQxVMNN+Dmp9AspzkPPugX3mR1hosbjCR4+Cwu5GBbMWMq9O4WOdmcJEjPMgZnXyYZ+M9KLrTk5
5A047sWmcfbpsZaIjJr59iOMEVZsxVnHlksr5equIY9Sv3cJwQCwNPSNOfi1slf2T17gaSGv546J
n/BWOa6R7eQXy26l1h2ahAX1+EIsjtWF/Nx5/NJIkSm9dqYviyXmp7geXds2ACijg2ivgHMtP35R
+DDynV/AmxnD+pKQM8XMbckggR3/q/ViEWQpeQXURbcA2wC3kdn794MftpSlhVqVVeXLqEwj8WPz
lN4nvi2ry7PeK5D4finbbjidC8IcpblAk4rI/dODHmjHVyQWz9Qxjx+4RuBu6CM4LyMJIVPbdc0R
0H/3scQbkPWmfmgOsIhgmVm41becBhYOUM3BrEcDEiIR3UTk/26lGv2g4NZ7Ccx4ZW+7cLKsPa72
l6bnUYewph9BVTJ7CsX/CqK9hxVAqoBIHsaNhDXhSIOpesidLy9H2fPqCDpbbkslG9oHdPocCffc
+vzmTu4BB/8aC9CsAg6W+jX/OcXdYdSatCYC4uPWW3sNg1BBLUB11ZKQgyf79GK8/ajm56y9eaC4
fRcWP/LftiH3qBI/DKT2N7IT5osmeJ94fH+iEInEqlv/iduo67Dp4iK6SPzk1QcWMmldx+iAIOcd
ehRLSrJfoeeYokK3gjIUD94IBQ5/qABrbS0FwTDCVqXKvH1eXhQQl2d81lkerVW+ZkMgui/P10px
KSB/R4TUCMqIc7Kr9gkWyaYVBulv9mIwGB8bL3UFblgMWgQBiwiZx9UloMCCSx5PJ5pTxEtKf7J8
V1YnXGcgWI8KaaJ02ivbC/p26H+/f49gWu69PIMWflbQ2OOn64ch+kPOewEsXgsQ2c8ObF5Y/Ke2
N5REymu3qDPrrtUh6X0on/oD3k5Mk/V20slrzFqLNytzO49lKneehOVvtLV0MuAAyZEInziVuigJ
X5Ny+yXm1I0F/TpRTb3CBV9gXU5jy3qTlk3DlnFQKqFo7K2vlTUb8YgWgWAzvEVBMunIxS+O8wNP
8CBL5icLanYqapjPN5FTMwMVYBv8+JpoWS2/6MmedWQruqbLTEvtwJUly6VzXL9dB8jQpN+OYLzI
/V85NXNmNW+03HUrJMDYYHDholjKP1GQCLvJ+KXNNqjHIube5R4D02apm44WxFpp4XpuB7JdPxXg
Q2jFg/eZE+xb74nd2Frh9/JL2laN9lCty1aevKFZ2JMjDESpJvVMVRKTSH/aow1dNxuOE6nZcheD
TuaHqoBx6OwyBZIz4wh87r8BEKXotLk9aet+UeqlDNmkxTdz8lvB3qcD970IyJpf86xuoQNYtbyY
8MImNJajxIVz7V7S0DRzbVFrEeMWw+aq3SmjTlA+v8iPTajHdYHhBWpMP37/e0dJwhoLa69u2lpN
NUIyhIKGVIwmNuLEg+l754X+qM78N+03Y2+BiF2CQ/ILR2EUWvSPc8P5Z5oq4qFvGEhE5MxZeO95
ePL645U6gH+1dTDILrpMNbJ8qnYiT7jA9lYQolRZx8SA8Zl7KC4vYeYbfDTXH/IQwQiz+8oh/sVq
wmCEFj+nG4uue4Mg2RZ9VaP+g4p4M6uPsTXn3DoZu8zVHDkA7eZz0NcdmTgOo2Y8keM4H48BJiPT
4oUwR4Wr1ApqEIbR/aLgU7clhaKK1gRViyAaPbvU1grqv2q56IWUcnjER1/z+jo1Re644kFoQOel
4kzCR0dhSFb4YulhnZZw2F21CglkeR+xXgvRn32ecHpGmeLRBiJtLBQgm9POnor5O5dZLpsp95vz
/60OhjhzNVK1C+4XnxNEwQMBFku6+ct/dAbX6YW7aiWPe0nI+N2r62Oiddi97rIcTVMfOtHbOPeW
lZNoaa4/Ma/kOdXJF366ao8Kkg8cZpR3ZAVmkL0LU6Jhln3HNg3IqWQ3ceSkaGB1/Dn7YT4BXwp2
5Gf6T8RVIktAOxWM/5wGL4ftWN+zqeSna5vjZLLmMz6VS48OXJD505fW4ew6vlvp4zyaYo43Iwrv
qm7d1bHhlCByXvm6vGwzXV2CP6s+UL3AP6DeIR4JCeq/t+vgxmkokmeShyHmdq6oZfOqmnC0Cclu
gct0GzwO+oEFLks2th7lN5VtlC/Jwnn5AKEWErfTr8Ai+H35jbfLSKZ2x9/o9oBYZjPapAh+w5ml
mgz1RpcyYzIC3EWxE1ZoMSDL3HcpiEnNI5lTYneqSRxBsXSJ2C189Grap6n7/WyWjK2vNHvNYdIr
dGwa0rHwMwLurTMVvhPwATXhRYmcAGXkMwRxxhhhJmnynbtiPDz4dVwaj/P+Y3Svm67JaOx8Ott2
Ta7R/T2MJucxi9pV5VeopXg5o8xNce1JwlH9u68NpqTDvBcfklym1gxKW2j/GXcMImbZZA90SLN7
mCzv9Lfo6SuJZ8I9EontwE3RsAnAlkgwUpJBBUD/xB6wQ4kU8NNHYQIfB6IRc6mXiZuCKHBk7/l+
9zICVwCgCkvnLFEzyI5dBpwyaH1Z5IJKc1kAPTi1yXh+CsCunK86PzLU1qOhIxhAoJ1CRPCqm9S+
X6bXWyT4OYL4MVKY+MKzac5ktDUqfxsmmzuYP7zHxiriSD6Uq1kXsmwx5sFknFy6N7iPVIoC5zkg
YbacCdzctbHkZOEkYKQlJAC68ZlyT6lbpb1DJRz34/nAZlHHBGrhwUv0MKVJUk+x14dVn/QHQmmt
tefNjEh45kh8Yr0jN3ncu0HgT7ayP8PIfTA8pcGOvNUuwItaXWTBHBkGDaZ60lTacyjUwLDoLv0+
rvcBwMqSU8HzP4SiMoEwwPqpRRGa2CjJtQyK8T7BwgpHyWL7w/mJoe/MyS6s2YuA36sNGYQERW7F
c1pAzkCYSW7k9tMwrJLlvbeJNN0yk8KwyKnj/BJy6VorfuI/DORgzvGImu26jCH3jEA1GC6CiawR
pv5Ys5Lfv3R6Ojbc5SHIqZ/TDlP8/N759dkzfZd1r3yHOleqz1wzE9YnC536rYw6Gp4A6o4eskqJ
i7NnjUuL9J3YAcocK4Oys5n0pbIUThmTAh6UUmuHGy3LBHVcNBQvwQ4S5Lnrz5l9KFJnbXUUEJBC
KUsBkUtm3/CJ5xOa7AxQbp4kmW442c2mLHY9PS9TIrGhm5ZM1W0y7NzO82RsCd0NOFeAsZsiOqkU
ebgKFFueBrz1LN55kFWHteBIMhJeb/5hYr+hXVA13HmUX++F+ZKi39/lSYxdZqGh9bCE/sU7t2yX
DoaLd1ny4IzIuue9BERAPL9fPbh06CY5kpnPwipi1lxb3emkox4fGddUOC31HK6EL7qTd5GUG4+k
Olg4AuTyE1uvNfGOVoo4UqvZu/ggGX/vV28Y2QKJQqoAkRsahjUdVdNHc4ttxQBYZcVuv9ezCc4G
Gd7uh8tmh+qYNGbIoJK6r/R8aGgbQn6Mpf5hi2ocCwepOTBiJ2TR+IXGYi4ZPQIWSapnfGP2QYYH
igQnMzRiPueN2kNrESSnes52JQdkPQonw45cHvmeK5TINgKqRcWWcUZ7CB5KbHL00sgq9Ms+lbDX
qC3hunYW2ELCKgFyrD62/fcWquO3bMZXa5M2AYTWyNdBKEmCZW74ZioY/LaqObBluj776hzYd+/O
3Frv/ALwBzxsgC5NTKr7edrQEz3IutSv6KxRsjg1h2XUoPK8CUIXNxj89eKF9yBWvCHn/zhRVYbZ
WG5jVdBJ90ePo6n7JbvKWgheISEBEIP/ODt978/0QIxw67V4YbbHes/JwOJfiBlbfsklEMpEEkYN
aLkCALBoUoukYMCKSeiyMu4zjcMU3W6f1xVJo+U9QgJt3XnKPIjRdfPIVsJ3CJ3CnfS434p1Lw1x
/8Ztu2rAzznU7tqNFeFURC7zSDY36bMSSS8reud5K9p9SlGCCMAe5xxyjOtetpCjb4DLr28l2PYv
zOPQIZBdmEZOn8fN1D2fAEhOducvbpbk/3bZdKsGnU6uONpB7Y5g4FuxuUo/OUir/Sq2u97A54I0
cZpeU92dAf5EYcxtX6ghpMx8OhgJqvAFY85s0/JXdRwrTY3exIDjf5JyIJwW2Q8JSromqP6AuUYc
UsQhXDlyUqTUnR251anhGckmgfUJo7E8jnsaWTgOfIal7v7XdpWyXjIxjJmdsohReN7XH1zpROGk
InxWShPT8JgCqmzkBmHqhILQJIoCt1oTDssnqPSvchdU7/Hc6i7T3w/Xm7QNIL5p0KjDSKxfRZSe
GkHicYOQGAbsGmm8SmGnTncuj14QN2De6pu0tMeEQgtZImoDem5UhzXGGb8b/BivEDxFPJc1XBAS
2Rg59AXV7cCoDe99Of108fG1NYLSXaEJ2tKPG1qHOuliefhCh1YHKvY9RyA5pHd5CyS5efqzfm7S
UzRYX8p3Sf3A223gO7kSpKLGoIO7srfYugosgOtKLg7iHySlahgq3LIqZk092ynO7ljXOvK+3bR+
U3PVgynHgyW1V67mCQVW2R5WjutnYOpiOy1lzPuGmdXLsbsWwH1tYYg8Id+9/kYiL1DfUVg9oDZ+
n96jaZRyt8DFqgy3AVrqCGvMMoLMbV8QrsutO7j7QwQwKcou1pNa414Ss/udv1g8QPPKjK5tqStj
PeyUKVL/J3xLvrDyUmXTLwWZDlB0QdFn9GUEh+R+SSuSbgiYf7zWRSBLBhztiL2OWjbc8PD9TBKS
967CE+Io+W1H+tgCho4DfliNUD+jy9rk54tmJodt5QJJ7A/9mYdjFDFG2MWnYDQDgbUcrMZFEQDe
cGXYDGGAsEqp53ICwZcRh2Y1TE+MBIFoqMC3+v/hYQmVz7Fd6AsMqmcfE1Rns1BxcGQFtYqW/BG9
7+vOFzH/OpaJxFs4pL3KLjb70DlxxY5vCRiWAjB5a29tpp4CnG+EwvOHwyoOj+7pmw7G2m2kYjWc
tRj/wd5iyE1iWm2uOIG9upeUtAtJi5k6c4hcG9U/KApxZGbe77D477mmJdO5mgsWVCXoRQ9BQPQB
piUQnvjwlC4Xf6knQXAvtjo2cyOxeqAjmE/W/yXatXgKQVkeln6x6IYjnD0A9+rruA4zY4Qa+fF+
9gIAfjrE4Lwkn5zNDr3oyUJZVl6POrjRa7FacBakAnADgiilxFfIWFfN6bDZMPs1lw5nIDjBKrOB
/YZy0qgl+kRgQsu7ZiSRyV+ExiENFqOxmMGlqHmRuHcyqpvO15fJSE3oU5q6psesaW+9MnLrn4MN
m72UbQv7mI/VX3QIObZ3kJXUCDz1mT4CStcGvdhe9LQsA7egvC38eefBaZyCsxMeqduMyKjuqLmi
+lmqXB99AJnCqrHckJwzOxzQAUTLPRxVbfz7w8ppcu4wxsaNwMma/pBgU6OUOo6urHDKEcohTiJE
7YkqWZb6o1xs7Wi8Q1RmHPTJ6Y66uI44Y+a0gbof86XSFvoiNiGU6tN+tVhs2krgwmEjiYbhtYwH
ULjCbnay442W97Q5z0bCyAPbcuTMBK3JnlYGYFIH100XULtusDBkaxjjbkoCLbJ11qLVEk40xJwi
B3TN6XEHQRE6CWdbE9Zc1rf9kQymKM4Gpr+BbUDiLik64VSLIUPQx2dzltrv10ylaPLE6sgmh0Qf
vT01oU5T8tpX4AtOTTLeO065UQJR3wmmWYBREXbyMQPEEzJli9JJODkhjBn495fSZKvuPRDqAyPG
+gm0TmEIA3/bQ3HQHFImcY59kpnBd/TKGK1B+gN6buho9LYg9cZaMM2ZTq8p0HKe6O0fMuLoC2kC
35rg9Tpg1I1o21Usz0QP4v7FT216EkPvnsbhg+Nazgw3Q5Y78jE/Qh6dIv45JKPxw3mpMqQQf6BK
bNFNCWgCWoUeYIiKKMhwyBC7WhhYz550Y+aQw0JLGCAKB3gfihnHIUreQsUtnTYQp+0rtkuZzG3d
ORcUCjadM45DJeCtRQlDeClqcgHZ+GEaUivt7lYnLaVmYYs1GqRAinO2eXBTgPOLjJlImx760k0t
12ZFKL4lSYK8YBbXoCh7DbIudaYQjbIH+eayVZhGczd7wILFtoTiQa0G/1ypd1poXmKlH+p1NDh5
mikKkry/QacykGKiPaZ37s41qUga8ku1TctM7eJwI4g3+QPGevPFKpjiFNwJtBdyHYDX90TXCmE0
Dig7RgpBo0svrT5KjPO+TQf+7MwStdt5kTChH8RVwSuw/zJMrPD0a16BvUaHm4E25pA3naCQyxNy
nZOjFnxpqlWJypMB+GnW/yVBFtV5I4Hy0W9B/idHYrV90NivW9Hj4v25BUPtflkV1sbkIyiThSsX
zc60LPm4umlvy6x4JCAXbHDcqoWQE/IxvwLj2MImLlyvw4kdpNqQ1gMaA3VQDEMcXrUiWtoxqwRF
C/OWATG6C9joNGOd3MNCKT8RhQlMBUyciacS6oW3mNhXZstx3e1aIegEOgw+9TTn3C1Qa/QACmDk
Dy5rEICC0J1biW4MgzQOroX9gV+f2KjQgA/OV07fIN1OjunS9fa3FxZJiOBFZTJlShjisCCw7VjI
maIeQb3EYD/c9IjHzwoxK5WwXxDg0DeIAZ/yeQ7XH2iY41jFpcORQeyk809LeLybEpkWS3pCEcn0
z48JSs20D++0Dm+jg+yZ9h6EaTKOYEse1aarXw56vDV2OTqPmriUztTGD0ZTnaQQ2XdBC2eK78x8
RBijXSqGOJ5YlnQNdW7so3ZHT9cKCD/UxBi+n4rRf7Y+PTLPCfA79XiqWoXE3nXKPQ0lzSWsibc3
tGfAcsqPUTVPhr5NwFQhPhSru5ZF9Rz7GGckv1hfP5ejcIPIlDv8aSCYdesc/3t9h+JEIN3KEbUK
nxG6omxVKytSgVkZx34Vb65zDp/C5YImxs9P7si3pdOWC2sBoXcNGzdclWMonBlBflBJPJdAtjEP
zHxXfMbD5wxLNJrIQcutrm1zoep4DB8UMitcZ/XnfMy5x9P+o+PxS8yI1QfXwU/w0k7oRip0eg3l
ySSeg/YcJCWd1of/mVh9PRULaSRfdPBLwGiQIQL86m170Bft3GyzPIiLgRfirWEH8Wu5nCMKcXMC
ob7rNVMV2+z2z/OqmR60CYF4Vb8iuT7qADYPJGZHf0T+iag5bj8EhExwIuifWaAwPWiAXRy6pBnr
sx3RuQQEX7O5k+8C7h2P+rDG2+Lc2Y1wKqqzcV6DV7wKik0a0nKjUnlwrd5JGrrkrvEVuDS6Vkh0
ylGDnw2YdrN4RhudIKSIDxCayMLf3VY7nSo846Se51qfjPfoIR4gf8ez8+728cA/XSCxxe/tLzi5
e2VCK0g8XhEdXQAgkKxdybLIHNo2zT2ZuRJQIdM+BJVLApX4aSKHH8jKinPN1i175dXxs9uCOYbP
AvdaaKWnxKMZUwUoRqmFiljXmBaIPl5TNrGLDnSgodmnPph3l9xDliRYA27VpgDV5oS0sddXuAET
nIc1+A+CsX5gsDaEjUHLKzl0Yt3J4ED28s9Vr6RnREFsSIajUibNL+72x42v6i3HlfgAqrLLcR08
VtMkWT+03s3AhtHB82A6dZ/Ikp1+wGer3fxfdYwE7kPCy83PEI7z18U9+6qUWQbdRR7c6MqAqfSF
xLvrKWFa6JpJHZJqFe1hjlCrBLcs5a18uQrPjk8bRs6dMRDPYMehmSKLFWsXeDuMkwpa8snfgfB8
wv9VQOHw/n28tcCuP62TXO5pbNseRFP8qS/7n8ICFY6nxGZ1QNw9scZOrXKTgT2BAtZYQgT7trfR
43HJkUGfAnESroP/8hPRuMiyJof2L4NRfA+GjgboG4fd5teVhA8146CzYRaeUgFaXvt1BwchwDKg
cX5IrT3/KXSmY2SFTZ9hacmRnMLw3/vArMZJODUW2erqdNCPDRINDubTZaPv4DN382l44fwkFt0U
S+9u7wXi+fAib3qQfb19Z1ENmz5GcIWPGP4GoNzS2CO0CJ5tdTOX4ayr+Q5tQu7J+E1gbwZdn6WM
4g8CSDyEDXd7WAxhNDym8fixj2Wa0C8pK8aOTCGw0vsbA/PvBYuQuUsYhWdnWyTpV6zWH2yvzZe7
FgxnAvx4KIbhyBPo4Bq4VI6jbnYQBhbH80kL+8IA2bVOW2J6rLurPaREhqYBJwTXnDMCSB/XdF5t
vitwicIsrrCyueIyrWNHWR+ydLv3nrEw+32Lv3zNdZUK0obAGMw6E//AiGTc1Zqd7GyKIqS6qeNR
BA9sklR9G+BVjJZqtRGeRd92qj/JGbjTxg6jJhTqhobllXKXhxj1eiqJ4uHm03sfynLi0BP/tWbC
8zyLGMPoJG5tOUI1eZx/bd3X2z11Q4vLVKnHgK4saEEK9AebDrwPvbWiSfUeo/Qk67TeoWR25lfv
d0JUe4zcHWtRwio55oQg2VSIV/aEP4l9I/9j3w1MmiVncnOH+TYHHzS8UxpPiXga/EcX0ftktY9h
UAdIbIKxUWqmTjNHwyluCQEJfkQkz3s85vAcFRagvR6et5O4M4e8COAlVMIRVCbpe/k/GiEB2wQE
+RNZBrTbs8BzNmKMs6YawgrBK4+kW/lT7hHXmtyx1QtfYKSG9QaITbNWmSVZRsu2tKd3T94uluzg
agE5EVdzkxhJz7Eevq4oQ1hj4/Xf08bsvkEFDJHF2mUXFM/z8NSjWaLHE9fcv4s0FnmSuWdCOEJ+
CW/89oRXseft2hbdyuaoPQh5i+Kpo2Y74LSaNHqN8IAF5zubmgAHF/EnGmUtEcc8wkXzX1/NDsxi
rRhv4+U181YGk9mClVd91ASLCtIqFmsFG8oerLGt5onymAUCOWAYsFNT42IUjgE9MLaB+QnGPKI2
ygdeUb063I8vhiCO+0Qo2G22dTvDQNUhxEIcd4B0XG9QUzEBizJjz8OLQvDtgRBeP/MZZB7fCvfh
ygbPmzTAkyhenfs/qIbVN2Pohxtd8JJWG10wcbcVBRhiQzdg74HsdxjpK1J5aI6XnDBxLokVopdj
e5b4dHcdMX83TNjs7h3Re8nSe38g+tLUaGr5Dpw/BXSAvvpbmMLOB365/XGyb0AoLlhXRI+drikW
d6GjuyKSqObjDgpPKbxRSrDziWCsWTyJWznkvxLhMiC+YQpJRbR3tQvEybqzLjF7SRMBwhDXEknu
mPoxqiyczE4DpetVokHqf3eGkdSKiuoNJR0biYug61KrmR1SqaAwrdkxXnJS5sfJ7V4E9JLw7ico
SoBlQrErbU/4WCK0jSYab0J/6bGxjsUsoVdEq19JOEAZND8YZlGhFes0dJryJ0UYZx7gf3qS72on
vWkHZHHEnuh7QbKnybxz4TfalYX035jRuKKFuWym1tF9b6HrASbkJgPkJXScHsIXCenMnjpAdE3T
1okWmN/uvBfUFVTzwqB25C9OjE3uy9BpmrZNlnk/gTbNd0acH4DI+3RfXRm6LeiUopMMMFRwjC2u
egH9ArMOfQ72VkZ2yJnB9t6CIay6Sb92DPZafPnqf99Gv+IaCLxW06PHo66irS64zoKPbw6U/abF
JCPufslUzyDBMfJCVqo9Da5UM/8T15PKFbc3fNK6jX0urJXYYcFwdRbEPKfQcDJbaBo8cMcRJE1v
AGBOctIr0MxPkAwuTQK+J6MSK8DPvBSg7vwWcIgFespIlK1DUvJ4uk+ZpKb9U8VVelNOoWH6AZ9k
l4mbK4q9sXuxCP9s1yHkm0kgkqC1U6cHx2WwOrsBDN4Av553+z8LABAUC3eQrmpEDMUJA01dnihQ
XrleBBOv+atP5arSjNJrQx52TkLeuAACE8Zc0JPdyREpcqzSj1Wr/e+g8ZeQHkudTd6mLOGgAYVE
05a/eaiXXxxaxp4NvCFU8h/l4H36hH+A3WufJljlYd+q5XibIEAaolwCIS2VSlfprwQ5kCyusXYU
C9/dN45nV7kgNW3aMMv5w1l+k5XgrinlVxpES3IVYyqBN2yBxRW0i92SmUT1lsn7B09uhlODPYub
MdpAlEUbt/lQ8onh0LMjm5+R8G7wJ/MJb9+IMxIW08VPf24OSRGyjAJ2uYMWcumuEyWcht6b6poM
P+iZZb9ftBJqFlmpPPp4n2fP+cFnGANReGOVbN+g5cAybKnnZcumzzPbkGUh6XVZm+FA3fRxydQJ
2q27YUNkL2ifLUL9ykMPcpI359jARtoVt+RP6YONJ7dh65e6HPa05nPdnzsrbZSJxEdMICPw9qln
B3x3Iuqx/P5WX7l5uZZ0UGitBG/XKYKzYGJON1cVJxZzjYMPV30EsjN+YFcYG2UDRPrjbvbfr9p6
wdvxJlTJum9rAvFqwpjkGo/g9sDsorhvymUL8Xbbl41sFQJOuKj24ZlAOa0pkJT51FXQn71NA1EN
qJHMCyHxlArProkYgrKijpJA3wvwHOsxTIpj9fuSvqczlHweSAVsXKQOVkf6X/cA9clWASjJRKpp
m4E5EZB288DDoROrf/xyPjL6wfnUnyidSYZFaORz0EF/iG9lVCQMzKO2hNXIEeTspz9yRUSPwDP/
qCh2TYvUqIYegKlUtn2XwoWR/c84rZFwjyCtRxQUXwsvgElwtMOX6/Ebk2lUIpuXBmFtnVecbXVT
ozX3j1KniowL3KQUdg/2Tx+Zm1U0kOfIuk8Ygs37qI53ZHuPoSJwMEN8icQkCDyGqUgOI048I4UT
YnkkPkaGYoLszDcz0PNRBUtwlClWjYXCL+6/MLzSRyh+Y2Gyzbq3E1QuT15u3x/Ei7hGCtX3NODW
ZsouR1bQlEKIU6NbEjk8ihESFDzh0vTVnbdTKYIGbWyJXhql9SUtAF3ONaYHxwxJWwTP8y1j8sXJ
kGzk9fsvaiTx9rd1iRuCYFWmqYg3PZfYaJEuBwjv7pVTXEhc8lwGYbDRtKOd5ZvDHPkR1W34qgRz
S8XbFGxar9KHnr5/fvJEY0Ztf6rzTmqPdubAjZCPm4ga5f2KPZUvNCDYoe9Y94/Lzurl+ISL51W/
n/BA3v1/4jdInzz4m9rifPA5Tjv9wWwVzys3SugBfZMuGn1+NPU9S/hvVZPyO0hnhgOjQyM3Eo0Y
R9BMG+0Rdmbg86RAAqGC6ZTDweC4p+zLj2dpYAnvI1fhwDDNRm99zs34BCLyQZqiVkWZulSSaJBh
BBT0GWtw3R2gs9GLue75sofTBPeDVFC8g8cmqZeJkYyed5EW+YdQAITGTWtuHTU8Td6oD4b+1s59
tlJerNIieeJpE5pPGDfXMRKngK95koqWZ/dbxMgv1DWVwB7kNn9Cl1xYBfLhtgwg8N/Oa1EIPhFp
ISAxh1yQismVivdYi1mLIfS8GBg9wKAU/0w6/RtSfukTSSa7BedWVJhsjOtZep2laeDy/DYpGAj4
Lzuygjk7YUlEEl7EOtZfV3M8C2eedfEuU6Wj6fRB3zvWmR9GVS7zs0jUa//Zn99NBy+yjzsnMFn2
9Qi37FMB9t1TwfU0EJ+a1dOl2h9qVHn1Cj+Gxpbt+w1kRLwr6qAcZebrGjhoZzJeZMKclaOsJcVH
qCsXNqDWAGmvGUPCHIYTY3Lv6R5AyGAU24xVJoNjKFa/2EI03FRtq5e6InSf/pn2fWiUp/6Z9W3a
6ZXO2SMYCJkQOHpPCBpAxhjrnYUg/mKRAs+qcvCCA68MsUs+Mf54abnHTGC09buoB3zyo6OLvLAv
Cp7Uv91xWhgjW0DwlnhVN8Y0LX0vTncmcoXy6Y+nqZMZ7BJ+HtiaDb985w5RewLDKWXQ+fyHdV/y
IUYE2Fu9AKGQle2IFgLDB7AjZdWmEovqEUNlzYikMFCqAm0GhQO9q9SSkU0usUeS8OXUnf0L2ZXY
61kek3k5Owr/kCi27OvO1dD65yz3RLcuV/K7mz1ASjZqui3IQ5QRO07y7ycbQf4tYUK71/KBhezN
9XnoXIXvF2jvgTE6Q1aeQ6VR4+ZX1vET3jLmMf/djGOwpY0w7A7769CiWDD1j69soIkdKl+oeGM2
Jin9gnvEWwzeXczA7v27lJNrEXRdJGtMW+WkYnMWLbMVqcM55ZMBF6sQSEoMCgQ+BZg1FYd3928q
b8zhceZxWl/N+Wn3HbeKVzfD+GLSJ8T0geBVaF+CaX72/ePM8UmpeQPJfOstGTeF1Cj/4QakrPev
ZAWEcQGAUC7mDvgQvfaC4/5rgDuWhNlEoOEdvm18SFC4Iv9L74jxw2kfs/9w87APxaVlz0BkoNBI
4LMIm1VT0tp16JEO9u9N6rDOqD1ftHziLS/hsqQupdl6xap6xmQeSjDwent/caWoRDSyMupaAGuc
x7dj+rPkd0NdXNJsO8XI66JbE2dbO+tFK0DgZCvGAqmknFVZ8Eo6mVOBRQced1Ttfzc6O3vubP/G
YvRlAEflk4VvS9/gOwtHjS+tWKyYRV48rGQalmHoIVm6GOA7viyHTbEMgmPIrBcycymaG8uH1PIQ
Ok2awRcNtdzL21oZmhQKp8KTkueXxYVA05ch406QRNu+OGcuTUdWnl3SUypuzvmUX5yg2jcOmo2j
Epw3Eiqxb9zKmbxznQUBVnlZYp6ulbHZmnw9UjmZT1Tdg5r2iMwWaOwrv8ArpwzRHRpvLTBF9CFM
1EO4UV/F/NB/Kd/iUBzh0Kqq6/Qy+rvIO9U1zdjaxQsA46+iRlO59un40SWQQuBWG2wpZKquCzPz
aNbiQhlCQ4vk8W61GJ8X2PIqAkdzORwSLIvM7W8856KFWiseSX9AWMIG/p07fwnuHOR5LSf43zQ4
nKvzL5bC1HXQRGdZkXHFmUMnD3WjdResHbrztOTgA/gm/VNH+puQVWptZusmtIUJdOpG3ZRgGam5
053bEWHuOhyoe8DpnTmBgjW3KJ2Y5K0SgcX6eXEz1BFmQjfF8wBM0eKdJO7sjXeBCY9EyZFvEQrj
9LiQ/9GBBwU5wbZ+XJuaxL/IeGYWQGP99fnJso1MWJnme25slv6dvgfs2J+qayqNhkYiOOAs9e6u
eOnuPdaL0uLgRK7k/FTHI1b5cgdrZ/lp6CHdY3vqIsX1ZBdbBoeHfVgwR1uRK9XWeuNQycFq6xNl
vXcARfGMHd2qfiGo+nXIaI2ObTkOI66I9OWuBvoJmqP+Paod6JKiTg1vvoMlWcN3fbUa08Vch0Lo
X/X4DBotw3pR0eBqHm+2K0IgvnMd50maPh2+eALyewmOReb4Nh5hb/Pr9yDSsVKY8ZvwDGogOuMe
zWnuXibwdZi9gxOSB1+Z49q/ste89Wks8o6QUs5gjSsVtzO+viSpB/krg05HlWRAuohu6Rp7T4Qg
oro0GieTfEW2cbrhBxRgTcOsOcU8YIFOQwPj+GE2wMtK6IyvKAoEgmqarqAFtPw5Y02lsk438/EI
+DK3zpzuxVu2AW8v9kQtxuLEXgOBxbujEnfxUPZ6c1Jl4ZXFfpHmdla30zj8osmdziCiOSajt4Xw
yV11P/h6xjs6yLTSLmDI+Mbi++2QZHsgXokVfpaR2bLWQU+8SLtRT8TJQrHRetUsBoeAMmIMoF9R
UhXUXWD1FNn83tjwvRYO7wkY4RHLFU3AxPBz+Kj11Spcn2oHR4H8jWDUW2IzuLqI7sX9vkmu0GcG
E4JRecwBA1g9OaS5i+X+naokceFiYrl+r59UGaJ4UviFYUUCI+nfJ9pgbL5Ja6J252dP6rZVEbUU
yc+4qO/iOfFvn6+QO+70HpBZ1CkZ14hxb3h82/8pdIcNeOJAbESjYySGrR7/2kdcUETCtLxd2kJ5
a+VAuJdH61dR1H247SbeFwICZA4XUGx3AQUKOEcBIc9qElfSLh17DQ+8XtV7gLHE7EH1IpFP7qd/
kSG83K5g3K5pAs5GquSBmus042k27UqQsPndHEUxkuizrVfPpZMxlpT6VusbG5t5L6yXkMNSMDIw
5+JOnr8Ovx14VdAVminuZVg0m6iBbjWwb6aDyeelAophDT9dY19WSSWJHCm/chj2un+cpWNo23nf
n59TM+XYv8v12le+eCQ9HryYGUOapuZOpYbCHFbDZo4fUImmtSN0qk/i0Am09PXN2zudTYWFPgdF
5k+yW3I6My34KPLktI0SIEtrRe1bd0suX7DPfCSaYLllpelI8WWX0GUhAb4fpGbEtGHgyheyxK88
TqoHAVKMajxstabVGyO4tCBfu3aksuzqd1xeLt2aHW3VevtXgb2fn1og2xM+AW+IGVM454admrjR
YpXDU7FiGjLQOEYu0gbSAnpehDZGInhb8EltzzClOhP2rX8URripqUI1gQRJVj4HsdHcE2Q69y7y
eAgaMJVpdopzLkp7WWi2OTCCQyGX4jdpnMiNSgEbBKhKdMv0f5q1ZpSY7Mu8Q1xGnHQZYnNFsM7E
JZQJ+ZQH0jxA+5Doxj5Xyq3tYJ6FDHFJYRCPoPVPrAhwQtMIg5Bxvacpa9kpQTmqnVW8uTdqhQr2
7AAG9XFKckL4A9oMjHBAGpjFNOeth74vHOwQ4XPZFFCPfRNbId0l/XFXwIfSWMPDuoEaOpP9Y4OZ
X1opRGfkmaQ1VZYN672kWod4jWFNZ2ZLGCyJDyanz3RHEN0i08JzLnwErEqhXk8+cKpFtM0aog0F
WkcX43dP5X0IsfZiOtKYDUerBo2hiCq3Eosi0ZgPy/ib0QhulJZLmzm42jfjIojPxgnX5G1XaO7n
EVOTOoIjWn70ZYZqc4z1Ab426aay0t5LgQRP4h2xgAtWv5fnD+a+FSrWGKprjrFQyxT6VRYSKRoZ
WOdercvbm1LnRe67K8fIVyxQFT10mHOyjbK+x1KriTvKMDxjp3tXGf/hZMXAfzkaJmdotktNkTHb
5OdwJe/U8NS9i/l+zXbne9Z/8abgoS+z5tM2RSwpWUlzlgz2tPA3b9xE1qhnSjSNJ6N1S+0q2YJR
of+ksgt6sJOCBlb6secaTp/kbSUNkRq+REmzNkmKQw2Io1BMD89ggi5lHOYsEe1PtnrAt6Orpic1
bosOD3cFjn9mb7cmU2znU9husfe+pVXbFdh/HzH+vRCGdLv6BCPKia3n+1ddaSbZ/giKjnK8X45o
nNQVI453EyxPfIV5Ti405p8VqrYPRKN39Dg0uRNEdnnVEEVN+KF+gYTKflWu3PQlkVkyO3bxaKgQ
/8uBfvG5umPOIn5ZU8b8q5rnfLQ5dFNwgqxuvPykFxgPC6wCTI+6vhpl2FFeWM1kq7ZomZQkVC2c
tErSayCW6IlrIX0Us0wjwP0afHBVdM2wcK+SaDOECe9leJ9YQQBMT+sx5pCLogkIsBHnnSgne4tw
TZpXnyEINaIPDLKeYJs7nIfNy2dPoxHotEDzhN4gx/1SMRsYLjUYlP125CJ4gMu7F+wtFhffoSMG
Idr/NPob+Hyef9EqNpx9YKMcKJRgAdSYQOt8nZFo8oIqc4UAlZstrA035kvSy3nN+zrjCBynxMdS
7tmuFJnWcXjtSfLTRb3KEcPHRKxaDAP85WmUQgvi3g590aB5b32jMgZxqtvrJDhNeNipfFqmPx3w
i4i8Pj9vHed/NB4zeqjMjbzKHY2jrE79yF8hkaiub/JyNzjYvSMsad8vi/akomEx+59P4Zi+J/6h
t1ex1A0CpIwBV0Obb+UWSDbf7/967DVNUKcc0x3XPtP4LBf06c0ikBHM5CHjfBl7EOgN2TchRXT6
bAGzrsdUMBIwVmjgPFqBUysQa5RhN6KpwZhBkZfT6OHowVK+HHxiD8lyB9C2FRp0UvXl48nzWRL3
/YI8zYSbve3n9Mv7Drh8ydFef4OUywBNakZx5DiiUV+ZwQnjzie6MkvYH/EEAGaI/Ax1MukUqgq9
8HVdGPPg+abrpcQuPSHTPR6h8Nj8grV7lcvBbd805ED0aUMgPJzqkP4gXGm7sHxSakzrzmRP9aG2
bhcIVe8Gw7J/J1/8JM/+7117TT86mj+VsMMZCaJnJlHg4X+u+DtZBCb1KJcn3jsZqgyOMoceviq/
DvT58Yx7efKrLUPgHtQbWzmWJwtp3fwoyzoGdPZAzgC7JsfKD/MmBxn4twMjYmmMH9qGv1sL1DHX
3+54pY+F75C90f/yqmGqnxl+8hUvFycd5EF0SS8ppZYjn0B9zry77CxDo5AmjoHWH+IXz3IBrQkh
ezTt3b7JDioIA/SJ7BYfl/XespDlsXJ72cuUWHRc31N1B6n//5Ezl+j3oGLJfoi23cm81HMS3UfJ
xvzmzrxZ5BGCorBBI0oABChScUw64ZL5rEVDc+EAtAyR4rCIkbZKwoASaOYFHx7Gppxe/UiBG2KL
mEOMhbCKgC1t9edhq/kUk2FW3uYitxQX9mIBN9rSS2MobnCBCeBp0qlRA4yuL/N0BhWaFTPh2HPr
35/FAKvGF9VCxV9bUQieFT/gz/9b6TFV02FnGsgWWVlbv1KNQcMvkb8lcYDUDw/H/HLovsav4TfJ
G0fQEwjd4St3denQ0bC0kXBn6VLqRqarh9kOJSrx0dR1EiejBzIeIiO/fRhMvd9ej/1wO4TfDEdK
HchHQqbsIuDNGNS573Az3Pgn3YPRmzOPEmFRgNr431FeBnLUN2uQxve5K4NpL/ShqXRlH88qxV6U
lbPl8q7cyZ0F17SMCAQUDwlfUx8QP3EaWWCQTRlkmlx6SCj6Ebu59bmJ3uQ24x3WpW0w/HBk9RL0
d7RDveRrbxNIs8DC3XA1Ow/7pCZRLQ84NKMynQZAR3FoU7lxNrB0bnRWg1XmCJa+aTW6KdhDdRq8
BerfAtiHEmdQL8ff1v3OSRQPJ2lzMzcjZBtqjMCIJqElIc8FlceLz6UVnuf62JvPF5Zo0Y5Aw6e4
ly/2p4uJV1gVT8b2rW4qkWbHyjq2mBGdBodwZF5V2b+McvBkSCytDmbm7qZgB9vFhcscA7fRGUOV
o3bPx3SbLEgrx3g6OUP9VDujNzv2i+yORgjFnj/KdSWCcJkHFd8HzpqOeajmfSaco6iEoqj2q7Is
XFfT1phYMjTF5Ck3FsZdLVKI4kqCVV5HUhkHm5B7OoqzUUGXpvCF1aYQMQGQHjNTPG7KRKkVAwdK
UQVHWtjrBRQOSY3ROE22/91AiBrKCO0QitYCqAjpHWeEf0nCxNDkDv820mjZt4wZJHPKMZWJ6Js3
y2osNUfjt7HBiPEXGokZYWqW0jeI8rksq1+cxHeGqHERQEnHTXat7eJO8nTX5CMBjo04UAOywi/U
7N5ONGn1cQh9Sm0d2QspF/6lKDHoqNYUttEdFv3feRZXQ5owwQhscYgo5ffSow6Ug4SklKlxLtGw
ATyV9UBaupjPdmLgYTFmCLLprmI0sAU+9fz6bvnrbqDHiLjoH3guE+yUliCZ0CXB5YLp8eRNDexv
wPzPNuOQDfRR5szhKDxSkOQw3CmroKhoLrZcZRLPWs+KiVRb0dBJk2IRmAdm+zCuAuBQ8TQmRM4A
iNAP2I9UFOBgerBUCWM8ul9cQ8120rG3sgeLtuJcP2Q5kZXMcV1qjW0ape29WCkxBfkH6BiH82UP
rNq+k2ng5hMIZ/4VFvF7duOnbIWRFBimYuGr02v6Y0DY2YI6Ah8SyfZENR6mm8MUstR3HkCjMTs6
HWhUgbB59mVLbMLzobOhiIJu2nDLYvcWZULNH415MMh2d/4dqHK7RbRgKdy84X4Avx+yxKOQn4iG
XDVLXfJeZhcl2170EwpIHcju8zl+UiHgisviRSJrc8rXlZk007oalv9yNS7ky1C2UDxSkcMF62p/
EgZ4qFv5u7lb/QOD1TdfETTM1JF2ysKv7TNJRZEcpj8Phbg+azguDF3jU71ks1ADiVrPsp+TVCSx
mrdDH8MYia4Fuu+2G0sffrJB8JSoKoNqr0TbXTbvmkx5X+IKsNH0uiw+e+WWUcHPPKE8989yLtJA
vTQF/cy7GxXzc3VQUEetZo0jqI9f9OIEExjJGaCMF/Iha6j2M8ZklwB2UzueSVFFgdEcTTKeF6lt
RoOhLa7RXPmsXR/41hga3p9UZfAbvXurJLdifXJgBwSijrL7lLQ8j6ym2wHZ4+7uXdHNKKv8F+nc
aQaz2qAkdE/g2zbe5zF0x7ViH/agV25L/LjJaSZZb6PpwD6gkVg3i6oJQyyJJ8jLJGCKYrsPmm+q
xk9mrI9C6pHwO063n0mdnzVYDOMco5cQjXFZHIo2HFhije7y96e7ZBQHiDvblpOkCd5wM+/XkS1j
JZA/nspq3jGzKgzK6q7lZkFuIy4c1BjHoBck1nsxtVVAoz5SvMw+4O6B4U35a6m3hZ0sFbwTeHCo
NhG38N0ftleDwTH3Tqjyv2O1clBnAFUoRgWonLHbhVzjLlq5PbGbt+uNFdNOX/SWM4F+t3Z1M8FH
j+CELRxaxy/x5sS0I725Ozc8jSURWl81TDanyq8tiDKGRWZHj1Tx32lWh/lUfT3m3/ER/v7osF8p
1wFRQ6AHLdLfGxBhqHCRZGPbYeBoZIWK4yIcaSgp43SXQaNU4pV7XP80q787D/crMp+8remyDSIT
x36wljrosRUtO/UDhRztgEnoxAKuIvwSKzdhmbAVjOE9ZH5itfNTUOS4lhTRE1bImh61u6eeg2ex
5Rbn7dmd6nQPqtUe3Hd/nNm1AsGKz5beVC2OH50WESKe1HSuLi++2t5M1skUf/t7rMLLa9sk9FJJ
dSfTPA9feZUnNgJr6sSaD4XCA++J1O15MG7GQmiwq7d/OnMQwmF8qqi4er5N80cOyLAvzu8m+QP+
8i3wvtxJbIhpWqVKMUmBXDl5w+SYHuilCJTi6oLVBtEV40mzzbwua6nONVzz2aIIPypYBzPlFy2L
cIYF9HirK/5kiP/krEtf48CWln8zRIWeVNMf5D2By4SVIm8+qrDPN8x5BWNZfwewQkJ0LaYQ2ruL
f5c1Ub+oxD1PR9ZonJkH4NjzmFa3KzhhY2isuAHB8plVrlPXNitLKvvbkEKT1344gBe08Rl0T956
Gpfralj2HP0vhhawHNCmXP5tmRgkSEbvS+88zVs1E5worscL5T6GDa0JB73UO0PbQMQWp8YZULbY
ok0N8auJT4z0mrk/IABHfR7e56SZabVDf33nPU04CbBG1YJkElBCZhMw/EF0XO4DnhJpDYdGd/0Z
5yBr3ki6G+E58IP1oF4fHjYBfgq1nY1zXzk68KwilsXLI7Dxm24K+nGkF5vGOb2xKo9yKcy2rtP2
Ry1DfGw4HGnJDZ17vHKae5epyPpoUdXsWSb8dP0zCyoBjJ4xSF57bSvGHFto6e2VQEGW5YwI2RRE
NRCvo2P94AvAzE49zt1sA+44MeleajCnk8yt5IlCkp+tIYhQ9bCMKoRmZvydfmUnMlgFL7d638fe
IuYeIzB5qiZ+LH2UEki7HmDS8snyzqc1PlgND7/nxeG1tNaI1ifIEEMdf11GsA4wQmz80wWTMFwD
dmGuWH4SxpkCFn0tcysd0DEp6VwJ/48giz3mVfhC6fzXDahbw6HwMJ4smHDtB6SZ2bCi/ilNrgaL
351IkhG1ushkP7nnflvq4ICWeeCszCzSF85A5OwEqTSA2b/yMB379f25BwJG1ZY3XJJhrdHhXZZp
1EnPaS0n2qIZpjfmoHcqRine8j4z2TpFzAKHDqMgIh5nLtlPMJFlBJlbhtLpdjV5lM+8t2wStKl3
yS6t7YUqISdk0eJyBATIghKetu3mTf6nwEaRLiPuiT7i0xXhb26IlDCKEYUyp6QsI1jSrDWjOtEw
AKBOuu+sDJqb2XTlmGdl8ABAiEy80ouV95CY2OU2i7r9eeVeOPPV5fM95cQ8IMxNpUQGbpNbM1Ty
ILGm4KQR+NntZ5LwqAkWHu7oFeWWYV92I99pe1MvfeiSHXVkG7lRQ6tdzEeAfNUro/B+lPPtk1HU
h548rTpnnbNEmBOjI07Uck5ZulCx72YWEfCESqKlIEp1dAaSRLL06mrH+KQVdgLUCuQVWt6YXuxP
iK9lHUS3cnKJlgqWA+WlMcq2X5aDJ3HRKuI3DLsr6V97j2ZYf/9g1jhKSpCNKBRb0w4q8RM62A+m
96RP+QeWLMVeYeAwahkcKJtyn3PwIMIvsIKwStN4MU8QYo9DPtb5q8yLWlLbg6v/hHqb912uLYMF
AsKC7Rc2CaVmNuZy6P/khLjZ9/YoD0q7pyyhYo0c5v4CrvnWKRPrGzr0nlm2X08BtvhFEfVEmL0h
aQ0Sb19mgE2vU/X+rjwoVEV5Ey1/985h00syptIqQW0LdCG7P2L0tdvBBVpNBmW1BTH1xXCmnCgF
49jRDVtaSeFf0mxyl34MrnVdEikrludLp6yAVKVK5OdDRggJC8BtxrvTQb2fNFp36jPqZ7gQ7dVg
SA9JCu1vjV7lba5qgOInHf7vOQqDoo+WwV2ev8NO3sBJeJ+fS0J+DIrIBDyY24Mz2ap/cRYIsXT5
Ak6UQv+F9CF3S4lLGKO+aXg5lZ5/9NKhERKl35hhjTmEJZYyDaoAibbUaxk5yLAsYEn+Y3qLogZA
hd+ZL2dOJ3paBzbP6AXIEGZ/SsaGjovZCjp138bpogsYiT9CM3zmvFhBV8pvtegjDD/yT6ExLK8Y
xKMZ6rJDmfF31knp9e++JMhA+owfeRnd9MMhGue6faFq1aQT+fEqsvbyvwKGnWPjAlyp406tFqv3
1BZU8miwl4U0AJ1o1ilzSqgAuez7Cgn8HLomwaveGOIg/VVd46cReQDTx2LXCC3+HwjXWxgDydUG
budcQonI9KL53lPxJQOPzjIqSdXtFerpxSBXMghNzGELN8Tlu+Rt1q+Oh+jiWovqZ/12iMlnojW7
82ZS7wZ9wibCZMiKuvG47AByM4T6Vf5ocnVlR/T3xpCVxfYJci8TpdjohcRxMhuhTRv1M3WWAn5E
TluAc4caQ6sEO1iD3uSGzkc71jhfBfRr7LGuhWFp1e4WD4HFeO5uPJPxsh2ULDpxxNs8KZCCrDBi
W1uOeK/ihb2FL/Y0f4hUT3Kx7OAuzcj8VqdDGu0Qn8zKtBUVR8hjbVsW1PBcnvyeIXxLQ04dQZ6m
4UCCJmfy+QR6GP1X1X7Hu3Y97Qwz5HSjA82P0NNDmthBe5Bw5OETTi1fhkC/Sb/+hmd/45gGdXz6
BDY9EZ5waVEQZ43eYgo0H6VQnM65nEFhkReUXSvgui3qvwYIrOqd9Pbm5Dp4/DqDSe5RP3/BgiAP
ym2Duv+xoM7fIdhDiCCWDC6dfQby1t5DfMiTcUqNdFftvPLfd7ZVCu3oapLR0PFnhwXYlSTE+n5I
ASB9MUvpqQ7Oza7QbPBMnL4FjyR0GQNtboQ7rfoTIruDHMem19K+WOcOObg1tSovPjWMf9Et9UNd
OFfqFQjGJRb8WO5XV4xrTMD7Pgb/mUU9i5EGh5QRFYHifnjlQXt9Dut+0vCOnP13oPfbq4cQe0Jv
6kDejoDxFj5uTS0jywZUl2JHseXC//XKDPCkqDqF1vLPzIdHMUAEzy2rsBEH+fk8z3XcyJzObZ95
fp1obc+wVFUSDhGPLuj3BieBrM9GFQWHeF2/ewxoW2ObsV/i7gic2wUTWU5dbCPtee/VZRez+4HO
v2cfiNlY27edNWojBiF/UpNR+nHwfItL9sLKzTdYKOoMqH6OIEnFImsXzq5m0w0R2t2wzJfp0IEU
xWGj8oGRA2pB9a+izyRRGKKLPGKMNyvssgFtijqGNjQ6P9uwwZjQ8Db9fU3T/NqaYC0CIrYR9bUH
TMgNYhdr0PktqXzXLpYJZ3EdW0Cj6TgsrD7rEhOHb9OHNJDgERVrver587vzrYOD7ZHfU5E5vixt
zBFzFjWDSGPcBE/POrNe0z96oEmAkwTqSNTPztEQFmORP90kLrU/7x9IOYg/LqKfirkRM6F6dQt+
Fn9SLNGxUbeqR/BKaW8ghRWYfZb1J72TzhtJ60Um9I0sZq4b+OWHUOeoPX5p11JXoxNh1P0ZpK5+
iGb79V1wk5ayqYr5kyfw7rbE+3GXBBRfoQVnTeWH585W570qSHP7m4l9UGB6ScOFRUaIE4f6a2bB
f4AJs0qCc0IyqxTD0tQjb1ZqA+OJo8e1CYAuxRlxNxsRbQhnlus+gN5LwgBhiWOmReMpjgZeR0bJ
bhEpfwHb/xhA5RrN0/fiDu3gI65FpcI7rTarFZk19Yd6gc6ZegFCglGPdDxrDlXInJNCEc6HP8St
v81OrnQoL5wiaq7Y0e/6nLITgjkhSFcS2RdLKzgLwU17dtJHDSZ557ukaq80DXvZyO+FFwPFNL6A
t1a5ZcgsXQ2G1JKkggbAYLkY+1KvipEl7zHpxu+9YEdHU9MGD6H+ndcLqVbw1Ur2SUSax6C3oX+1
kpTqt6nRL96icWZj4ulZ4/21FdfTpGGaG3hJKETye8HLrHDTsaOUM4n24DJREYJHqF9sJbfMQaq2
KudKb1iK2IInRIolUsKLgTc0MRlf8L7v1BMJoDDRGxhAuNIgY6fuefFPy+V2J7dw1XXFYOpOg528
P37S80MZW8Tl39ifIQ9sBZ0xVOe4z8FLsdwYLAYAodcqLpA75H+IqY0lcQZFYEJeedhRWG8ALxxe
Hmznf9EoDbXWMFJ7fNgT7pE6Va/acUYV0AC1deiiZcsjGDfp83chnp0k1jDf8sfAnYq7CBFUfWDq
J+ZGAhyJAPaoZIUPEKMePYALjTElTLkFSFdq3bDPaGnEdYTk/UHRLMQ6PTMQDpPX2Z2BLmoMeWAc
JCab3brJ16yfNx6yiQVPnupMlcdFfv3mXYGkT7+5ASkmaYiDMdAOqHw3Oi6LxMNHQLZCW9eH8Wtn
mADrlEqdq9zG1pq/caoaUiQwVw0NEYhFogxdApST0d6UFK5xKtSIGshQ5bcj2UudAzUsDXIobuom
ErgYCGaDlDtz7k18uOqFP3btDXFBb2g+CCaLxKQJa5HUzTlKaf5PN7wvX6WGvapCEf5VvFdzRt57
Y9cmnr3mM4JH+U9EpE44RbFHW4ASiUQ6ySDTQcUDf4vrtI5IqmVziifF30/rEp1il8fstd9hdgMb
+PX9a0DmLwD404dDd6C2J6uBFb/BhugKi8ShCeBGywYxn5KqDonwHQrVGnd8FWiBZ+Erojj5uruB
PiCyvdLNPjwefyxEn/u2wlZqr/IdplrdoeIdb60zGJIcwLJBuAGCv2NF3y/nbtvpnmXKjK5lfYOi
AGUfjgX5e6JPPPZCY/ebSklfgz7QgSTRC1P6+w/bxGEQMkuAdKQBnTk5WVJ7TXDNb6eOMYIf3Qx3
//58cZBrmW0uJR7w/H1VtMumVQa2Rv7E6wadk4XBl5IlePoYFQ+5neTOutOZ9TCBIRHMcKvhDKY9
UH4zhmTJ79+UXYG6Uee5PPAiL5fpbXiufgrLu8Ury5oKr//ORGN7myVi7ZKLv/wrCVeSlgqPRlQX
k8bMOG2RVySWhDZIVnzWTk9zKtea+pPeIyQs9gt3ZGEHsIKXxupiqrGiMQgpc2VSPBFAmHOSDpst
LqsHJcb3RAyQ8gLQIRnZeph6wpqo4hjKgraey8OOVKJcwZDNLMsVnit/d6atJlShXQOYoorxKMsp
MnD3LK4vab1ffapqv4WjsNyDTmrMx82th3Etz/ubGfz0jxWi6sckkuBJIWrR+bwbLE0l92fL9c8X
klqZNmJxmiXi56OBNbH5o+h7HMxgABlRQLXtvtyeXm5MEfQ8JuIVGV9QOcr4qzAhthUJhLsgxUMh
Zo5fxwRppR9kR9anLjs4ilpRdo1w21ZO7VeWmvprCLd2oCvrWbtbEVafjg9OGjd9nX+fmPVhx9mn
c0TbKyfZp89rn7t2UM+nalxtKXsbLWRX0Atu7E3pbTVWeOSa2+Ubpt+v7H+f6wUUIexY0EiYTmP7
h1KVOpP/ahSDjyjJE6yxE3PaCm1rtmwAbWDDlh4xQLTA6CYbiNTF5a7NO0KCOTzhlt26cf/jlmXr
pchjnsvoP7niY4ljWxfyRxuIcW0RfXAKotMAGDj8QVbiCqsAoknRg8ooLkCSokBANikujFM7dA0r
neF1n679EOe92rLFp89+wekdou5CxE9SAkGfJfiC6Qodbh2nqhbIIdMu1h0slmvnD/b8teAkTHZO
bT6KiYoB/ZroXR4k5gfvumMd8eTMv+2ppFvarMJVKGo3fBA4JRWlnvI7qlSlVp92TYctNPu5QGzR
aympZhZLotLDSP7F962jAwcpNxPCIpteJNxifpi+OJYXq8i/82g9hveYiJLmi/86fTTN0kivLcfZ
A0/KJ9/QoaSIAnlFP0ezaHcXZ5o4/GoC7RR/aFibjiTRmWpreccMLcrvgum5Uvf9BpjqeF1UAvWI
LB2ha3i/iDkHFxaPqBUf9gNYgERW6zTz7gJsPds6fumDWYvdKEWucXIVH9NYjBSN2HjC6uaN4VjD
6seGWM7g31Lz2XkCxTWUKdFkoKJc4nXdK0swczoPL89arsmHnoB24bXlksnFESXSrXvf3QvEeB47
TElkja7dOdjE22SxckODQgc45iELgOq95Jv2Oekbim0sE41yMjqASDPK8VE9JyNXIQUJ5EnezqM5
4ZhlynGJlzMZEV05ttlC9Elnsm9NQVfS5CydXorsz1lLM90qK9ArcL9vSY5AhRRcsvN/zfnq5J6T
fr5hO3DAmnYHY9zlyuKLy6+cgU9GXFGnOQ9zUi60v1scgABeruaN3X1eAsGZHZJQxYdQtNtkwlxk
FgeumBoJgMG9nZgMG1nx3Xv5wrGoEAN9lI8fNAUZnQOx6OtYT4mRS3mPmJ9Qf00WIZHl8c/uiGPn
DbH93/clHSUfS6L+PUtLUZw5KBHtL0Ha8GBceNyHBik/b6oL91iEzWgnpvCY8/JCC+opTYtMq14x
NM2j6uDMI7Q/gg0fL+DaxhH/bPl3faDDZ3J2qvYAj7wftFSPXgOnfO6m5/M32h7H9CZFPZpwyz11
yWP7gRoji4/GgLrRGgHFCALmGfqVhLpVWhdsv7hNwUIzhoy0mzQ/sRRLR5VuN1t1bGcUEJBXKeNl
mmj4TwdbtCtRfisKeQxv7R8QQxiKTETV5DR6diy1RHga35G6H7JEoX6WSDKCmTvTLRvRoWy+RFo7
gdo2S7HKFjPfIxGNwvHUIqxyAL3amNj7pKmVJR13NaDqLF66q6uy3tyJfNFE74uHeGiViVdlrwA2
8XskevUZaNp3nMxU5ZZpSrJ4cxaE9Gednk9V00ijU0VZdYjYceZylyyR+YVoL9XK1sk179fep+6c
2Tjx+Bng+AYpxowJGuxOfVzGVpiKhOgcBzTzwj5juFvmvQ6QsE9sI+2DF3rYhLdJ4j1Jyp0/E+Td
lqvgOq5j84M9M15FSrhoWOY/ErXxgqYAAxSdk1v+vizNerZkKRVkvS95Byl1EP6wxHtbNekloCuf
TkRAXv9rflw1utkFNwiLe1G4UuVj3JbcInIdWS9b1biazEUPckwKjxLhZsVdJWySzu4sKzo0k7zp
I2pmaXvzUxHNgK9q/Eii9eOGr1GHa8czhbeK9+5h2Q8AdVeS5AcNMuzp9HGkoA/mgFSTFJi2wb1B
zZv8DPLxtEl6AWFPJRtN93/xHcgHM/uB0eObX7o42iX8zoNN/BREKc4SCcDt00eIhO86YkunXxsC
/2nY2M7zhaFdDnAIhvJZqJP8mwKeNqAgBsqmlPe3TEERo6UOJhG9/ALrcSqVuh/K4DgEFjLvpQeS
wVBdJ4Putg5Z0pOjDIbsiFei9ON5bXEvh0nvsxMZZpdCn2w34Lw+V8n4bo1+jK6PGEv53wR7T9QF
Gr/eqVpqMTOhTPXg+fFxFVudOARfHdBc8EJzXpjI2wrVVU/bk5yTEQMXbnCDBOYUg7SV+uBkueUs
3xHgQymIcMrqXF9INU9pb8Sx9F6OHjWOX1cADjjNEfekwsiliWZZgdYPyQ7omNDuF+T1OIgE5tca
SkuFjHFL5rjV3ot7OKj2LAwHdDQrC+L7c/iaS+tr0KenERxdrVLqEeKy55T9YvO+nHLlzClsRoWa
a1oztpYTzQFoyckFSRUxfYEjd62JX+QHP9pC3HnCu8dm+wiM52/8fsTpRmoOrECY8XWOHbfNW3JM
YSH2HnJxJ+f4PZZZSri2LJXjuWQ7vx5Izi46VVXoNvkNy7JimzY+hL5McSkymVzsZ3oN/pCLMGff
/L7MFJoKzB3X1LKU1rO5K2dCGyOvYzxngYw8pDJ/LEMav/MLPXCSxcvqh7DLpr0KJv5tjU0IeqJa
q0havVUltgciv/JfytTtovrxS3dvhmFwBqIyqzHrMC8EbKBMqsplU4cQPnIng35ZhaJzOlILcv1C
Q2uAGd8DcmBRbjaybh6ERdhpbQYo1bPVYZ7hLL2uBwck4m8+WwcVFaoBHbNXPhd5w+jWeHivrato
RMljSiK5NFgQbBLpnZJegf28657ktQ4P5szniyA2Z0LoP1tZNaLdfxpHfPjpCOz2pycZtwKqnazY
wHdKtfXxVp0XoHDb6E5OuOzQgVJlWMd52xAT8DyPQ/9knjzrPPbXgVO1Bd44LxjyxFOGoa+gtVyv
vCvxeLg/Yl/xir3YQlaMghxSqo47S2KjD8/k8CvDlUFntZx3Ouw62e7Q3uubMF9FmvagHlM7us7D
fZnfPtoK6qNGKaTeoxMFPYZQQnvjadisqPTL0/J/hROqWRYoBVw71pW4YfWrvsdB/6Mz/QOle+pC
8R8m8F1iL+WdJZJMIL6JVd604Yz5BTE0gj3ZDIiLdhsU5T59mmJbAifIIpnoOhGZO8aB7JdNEVDK
8HVOF5QWp6667o9gR0IRP9YCCrr/jV/ry2RDNET4cdGo6feXMzcHwle3FB3b66sXXqBbpy5kjwLX
/HhIu3ss5DJwCFdCeLj8u6Uu+CwvyLIzeHDigHXCw2mG60HXGKT0g+CqYI8c78DqH33ocBzgSksR
iOnqou0HHnszsKDxi3VJvrLRoNdj4om1kZrfeu1rgZOYp4x8/xNJTIU33gSfYhMHBw3LjTbQfXtI
9IFk6A/kV+mq+NNSDo/EkCia+9scoVX7ENpe20gu7kLxyAdrRj6BjEZs7tSTJRZJrTtC4zIOixhi
2pLBQOw9vtbcbO1mzKsuzzXqxRIIyc8I2V3Bvr1ZdQGOSps5DxWBK0n/L8QVW8PWvPtdZqGW3qW9
qsC/K/vz8PskWZk95M3H+jZzHTNwR6swvJaGMyqyIgseJ/JZKulDeVAjLG3nmw9rJh08opccLBtx
9jwywUOCtaESUyyUqhlLShyr8/+Zxz5W91GtUR7eDLYcnMx7hvY+faCYje7rutmwwtHaPYclewBz
SiOTFb7IDwrcPgq/fdWJ5xsRDh9wKJU4lIg3qBy54sHkCQnMLe+bpzPGP1jqjYh+dEynm7asUTRQ
N+ZBHH3NNoE/DX9CgbsIBtSl/REAo630bqOUv5NaUd3pv7+ayTMLFRTCTPjk5dLuOh9Q5fM5xZGg
+oympfjQGn/G6qGyqnnua1w4b0sYx+EEZsVekKWLY4k8klQjpt0Warr5P7aLNoZJcBGU0Vc3w76J
LWS3IiW/jzJXVwEv6Kr/d3gJZOaRPL26N2FEhpjo7+4LLEEbaYbS9LQaI5ZVcpiImEZBH4PyIh8G
TB8zAdym+Vj6dUqurvRo5rolc5sKvSSiZGxpw4SFC0RGQLXccqFh0MtLSumcwmu1Kw3ccEvg/Gik
+jfANFd/THmWjbjImh5AgBolXb8u75OUNYg/aOrH2M+sxwr+ptVaLZ1jhcipytBcJ04CVGFo6+Py
62VTWb69iqJFsrSkqZtZdARGqsqozT2r26VlzbbL1eKiyO8F2n+sl2qnyOl7z1yYyQO5E0O8Bgaz
g+cj0SM1h3yw0voL+VThaYP/1IaMJyAvtsIoX16WEO/U7WiMcrfVF6goqo93uHCkMmd4AUqMpZzC
ujTjGgVl6w9P21S+PxVVnYQR4NueaCjthkE/LHXZo586/+Jjn/yraNP5Sk0dDJsw0cAja2bDuxpC
6I+8EcSBiZHfC08FsYPegYf1pxbW2EteudX9K5EY0BiJj2rHRqlwr8DXCZ0JTTUNPrZOIj89VlfP
IHpsEbIQzoSpRt6Hvp7W89EqffWBjMrlAlPsW/4uPrLwq6OFTPkbQUOQ2B3HoRkVfzmSYf75iYb8
eGoA+t/3hsEIWVJ/R72LOK/YWxuEFl32GB4u2DFAnLZN2XSBTc9y8Lg9cI2c3UujvlSgkhaJHZ1x
WQAtZgJAjKffqG7ck8b6RoR2KW7q5ROCn2SJxl0HqxdEtFSqdsDdcHbIJ2HlE6T79FhfuceaR0a4
9ZrvO41CbvrfZfYOX3Hg5wJI2uRnCWVu6pB/8CxnLVFiu6QogAOdeTH59ciYCIUg25fqW2AMwlRz
5ZUJPifPoo4EC8SjQWqhDvWkrajpvpUgmVMmLtUcmHBhPd6pqLgf+Tm3EZs1r8DNQegmP5/yhlb6
qh05CZtR8wLVRBpt+E1l8nDkZrUFbpqNxthL8qILa9aN4i81mfnZBpds/iBA92V8WKU/ZLCeIpnP
BDUdMlcZ0ShkbL8lrqSVcxSJhrhVsQbEqFGome1KvLjxgv3H8qPu7dRDfAIEkcL/GokYRaO1H5Jv
bAnuN0tBS5D+SZcNy6EEUIzdCVDuxybJUAyzrZvTyTT/NFJ7/Mri0Od6o06ECZqdNMFmhLbtgo+D
7waphXXWLqLrY9AECEm/HkYUqQKoGHprYgFlyTQVapJP8CGNs0P3rAhCXEyEUq2rFP/gesRmXdl0
DoCi3eiqbrfOQ6x9vcUyZMO09aR0+thvSWjt7LD29Ya/d3Gi/9WjpYaLAE3+rHyu4w4KJHnm5PZa
TY1J+TkwB8mpDXed1Vztmw3eMOlozOK6kpWWj8/YNEBAEF6axcLq5VZCDXO3mQQJ1/a6eYxUuLEn
wGuF6v/4TRZcylxF1M/h4hGtDnNB/EoSC2W1/cib/8uVQ8ySHZUNWPSYHnlBL0EvpcCU5MQzWBv0
eG8JYVKkSE+1NihOmd14E/0Gh84mkIMBhThERUhngeL63a8yzWS+PS1k1CHHA3IEx2zKTccoqN0w
mYNQWRMdPq3m2MDbjGXt0lLuuKsrl6vDLZzcRugEAjhQM/jRT0OdV03pxMOKnE5jckuRa4FsAMd/
6gH0dhKdY5F1VPZjPhC3M8ClXHU4UMQmc5YIRIZFQkZP7WKZ/2w7amLdgHnBehAiGMtbOFncBEjv
NibR0TS/8F1X1wTkRZvMt3xNvQGF72TsXudQgVu5COjKamsbjfULTP7BXc93QH7ml9QJ5ugm0GgO
cNXLj3nOtbTwC7mj1sAnsVv5+5SqLJ1JmwjBwKwG/OThpFh9VZbkdvBWWM7PRWncoJqjDUrs5jMY
xSGrzNfguBgEW00jdhYqOGMd53dZJqiu0s772S9UcXY8k8hQ83+pGT67SljRkH4bn/xQXdiLdNFg
gmLGD+qwn24hlayO6GB5RBLnv2qEPG/j9//3Ebxou7xHmnHF8YIomeQf3q0nye/B5BlxPBCOGruf
cNyHQrnGyuaG2WvnCTREuX3VQ8EKIYeQChRf6y3qniBynzgn0qXlxtrQEdQwwYqT/Y0lcqp4ERzP
1Imgh95xHNzldYbj50RGj03875YwxNNTta3OCVKVnoftHT65xHNhbPw3P2GXoTA96qUpLxLdVEMD
Q3k2lWbhd5sUAL6dEQBcYTNiKhzWrIEYmJ8ktfyhUta9OIuArplJNO7cbHl+QWIVBi3XkLmMiebX
zANpRHUYonGC58ymvKKEUUrMvHSj8KbVaHTVzcltVYfmf1X1IWmjIQyGdqoJRUbABDMHGk7OC0Uu
4yo8L8FkUcV1Rj18bLkhStMLsX36Im0toQjdfy8xBOgWTFPUMPW0igw6sFEpVeu4JyD8aRz2lsJ+
xodo/6r3K0la3E+eNiYKgFwFasdWMHGh97pc1C1kOf+kd4dcnj7TEQtdNVAptFMMOqkTgtCTyIZw
ch9vSzEkim4nC7cSgScXgybM76PVNkdDfkNHfYnKUKlBsz6lyXdgVlC7UyMrTVlUldQvufgGT/pe
A8sBMH21sl4R4pSMRMbkjBD7lYF11nJPi5MmofSi+blFsOF37zOWAAdiY6uxYVUVumaOh7AAmT8E
3Kzb2zR1106XpgBEUm1Z/69pU3rHHRboQJ4bOtmqaVz124SPW3vzAlq0BBVJBoVbe5P4t3uhgNG3
xUjcgV7YGJNIO5zuCRPV/uN1y54BGRHB1ERvoUJ98M3SPJODq/dMjmQWwpYAyBdT+pBqEhxbnyKd
6tviNMkWlyeIsSDTXBjHGijty7rrSF53B/JRPMvEI/lttMciNYUtlC47p0IGh3f4vGKYtSNoXSKK
xj1GogfixAstigtS7gs04psJNsZ7T3U/5D3e06yfZ0CeiyHMdfhelqhhsoTBhqp3gZKRsBgtPjvQ
R02CtKxHKgK4IdYDGkoSpA9Whou0qjH6kXUAzg4AkprUjJoc6X/evdPk2ENfiG0WszovDL4OvQYj
PkiqawEosUFnRBS8TaJsFU47ahMlTK+X9QXrRgCNgnw+wplholS08r8euRdMcaJ2PtFWJNuDmmcQ
CwlLYUg5sGFeIfUbMXueJPdRh/Vx9ibVBkHx3Skb+PPEDYrBO/Iv8FbqfF9zlVxr3Hvznl86GsjB
Lnq9VMax6ZQBJfYN2od7/uS90CjnZCULIrkTF/tKT+4yH9HuaNyMDo4Ws4yxhnvGIpKmGOcCN/Ct
bZPRtwCgJ8MU64ycHEHTi2JjFiHM9QyOVAJK5HY/Wkh6RG3VzewBZhYiHHH+Dkh7CK+AggjraxqT
fIotoO0w/30lSr4uMkIiU+7FAjb62aCCTzTFJ5p9fqDMCuIL/hZ41kgGQO6/ujmlBf9Y7y3sAal8
JhQppprm6ZRl6pz0oqb3r/A9T7OJoHsDkN1cOv4b1rZwIUQC+Ba/H02ugRLlufOZ0G+O45gFGIKo
9ffGs3THMmK87KWNO6A4aRtV/cuiHE58f1BUePcTZSuG1EREXmfqpM36vHuo49qSXpocaF7aNbTL
RTOMMv+82OWRfqDLrw6Wxe+gKIHuT0BdXP/9e5LD3ef9iDgXsiH2g6Gm6Z0ZWrg38eA7QuOUoHc/
t0DPb5oyHFu9SdMB1yl5n+YwUKm0o5h/u4pzQ/pH0JLPvtJLrvrPtDQN8OyqYO24BjIZT955OYCH
1JpheSnRYi8F/AadWgvTNNN+QjcdaIFgE9z5nh4SFxht2ZgpL4DQUjeiF/34II5di0MV1MgAuZ5s
+ncWZ8RC7GIGxjP+faCPDWL9xSrBI0+rP3Gsb5HMbNp3c+zvlleN2IBPH1hMvrvBmosxVYqhrpO7
Vp+SEfb0Q2pIPSht52BzbqPNQJeAS2drEodGnkYOnpv5PpOVCvI4FXnlSiZNXJwxsUCTnz21waFk
COAKX7qUV0YqEOPYCe4YTwjDoGC3z08O/9uPUfQd9TlzjLwff76gcjMFIRuGltbxmnvg1CPKyGCo
ar3ScYEaNcxZpDiyEHYlyDNhJ4AcE+y/Ev/RjJC7NdpDQApVtQskogtGVSk3JprNT4br0zqzib2P
DEeIXULTLC4JhCrGtZifMFMdI8mLFaUDw/B/cFmcxnHiH1mheiE2JikdCT65ZV04MVqL+aVSrPtr
GFxJPatKMh/zp5DfL3tFjOW84XYUMreIqDykAmVNJkRg1Q3GvsGIcgEXx21AEp+Pym08lxTu89u+
aZKHtyJVN52oKufnK/iCzbiDhUI7mfOAwC8waq1Msvj3R+JCyCfpU3AiF7QzK8iew07TDX6v8XFn
TCyrAmx+rVyuSK7CGDAv2/wsgEHHfghPQw4hLpmptqi911nsRMJBFUI9Mp5xoEPFuezFNX+P7Agf
RFUA0uoNkTjGNJ6+wgdpppiXzpTuAH3+LSxIzS83apfgmd6Z85Jk7WwnUXLRNfneCk94k4Ld1lbx
dRSonm3ILuOwDRrOplq4zsebVpxeU/UVJ/X86jJMU2hf3gIp0GNsmS7kQaQMUjgcn+zzK6TQUf06
Pi4xTT9fCkvANTsVHA9lhDU7cTebCxb+fnUrVqU6cIYr/sylMcGxgiZd4ZcrvPjhdD9VE04N2kS5
BXnQ5BQqiX/HghxIrdGhUUDg1t6huqoC0UNfvZj5RSj0udT/RmNoUNdVRvMfCR7z7gkPS8QlC96l
Yc2Mdvj+5Uv6M36H8sZYrTLWnmJRYf2EajdsD5Ju8ENTX0tJZZcZoQh/HXF8dmk85zHhHjFsoS1D
i8JlmNRSAtxbTaU+3Zi71+2B2wUDDZRO6y31E5SEl8dOFfzQvJ+ad7jNLA1beCLUbGgK6BR+bQOz
qfvMfNJij2cCC3YwqmR9XM2BDAHrL3rNLu6oKthEsfxpj0CTFIy+HtvmxxCXdOzVmyZKTgBQ1aZm
iYnilXZo5xf0hnqaWo9DzX6zP1Uz6p+x4OS555vNuTafq3vxOlsfoH8rtI3N8aVXx9vUnR86Irli
ohQO+rfMu8N/7VfhBWw3AVYNOqcMZs7ApKmMyR+Kd8bp0nADIorL+AHcu8ygP0ZLbq0xiuy5GjrF
Y0ypB75rlMh17F8ospifziFuGb4uZVwZaEzJALttwJlDihSiOc7E+FPwsfPQHMlg/Eg8J5isSwgG
6n63O0Ai7HHBOMFncx+FUyh57BuGjsDvSrHdRvTuFImjupHBP/uw7ZH5bMCIC0z3WECYSWvB/0Fw
gQFh1Gyy8Y7/0zWWmPFFq8yRBWz9JSN0ddbjo+mN8YGKUB59Wfz8Qr3mGFExIMO4JD3kkf1ik2qh
iPrZUvhq+nGDCfpP4CW/x1DTq0Co1wep+W4vEVxQ3JBp7bwQomX14/cHIney8rdUkaWzyPov21Yc
jSQL386H3hlwIMltoFSxf2mOsu3wdDuvGaN3FskijJiPlPWmq5k/KLEdryKBjED6LtZ28xXyYED4
JUPlOPsv0agpHs59s4MyGW4Drs6f94/yHDZId5APOPIhOzVVT+sCuWSgkepQIm9J81COFxfg7WxG
IJpYOsdel+wJyDOwqXICM0HS5UAVtvp+dE7DEoej2DsYNYFsLnh5gwgkyaB27+38R2BuTDV276++
yoqP+HZ1nhbXFqQV0npp4FuwVPRZ02e74qP3mksdPAejiItVNVocVVgEV+iagD8i6zbwRHocFenT
z/JSa1J+tv+q9GmCKLDbV9ComhU7lP9PoI6PAIuxKFWxmmyOYZmTESXNiHo6uEDzaNrgWSFGckl0
O6/D9QX/YoS19dIu4p5MH9nlD1fyenQ7iFFm57dMy4lfoHte7tmulph5s8aHZdYVEAPj8HrKpm2C
OdQzDur29q5s8GRpHUDlezNuLSVYJpjoUda7bxpHEgDSXAp2fWmJw/LjuzTcGh4BFWPiqdDH6IOi
Dbd6UooGo+rFrCYsHXjIpIs2fKdEhkfYu/3GrNDP8HKsNlr7j17kG5hJdDfffVgQdyE43OAdQW/f
7Z1L3z6qBQ4aDDsZ0VfnnlTPjypqdGw6+aY5ewVHg9LI49r2sfAAKq/5e4Cgg2f1SDCDFde829G3
jqqPxTI3/aj/ySTwarRdBm7y4U9OlHhMdgagjyabsdAX8BQyA8W0U4ebFw+mf4C5hIa40JeFGWPV
WTWX69PAnNK0MIaLduS1kADImbTyblNllRq27nhr7nzei8pAFKwpb+eP+VPc9aLBjH7moitK8fce
HxQVvHPWd5U2v4wGld15ffpSdZnSm9PGHwjp+cUAhWtczOdHo8BnHMAAeHWOYdheVSaQ53NUHbq7
+OoO/SjfY/p7uzpHXm6dMBHCdVSj6FnNb42CpitqRv743uYk9Kas9CUehpCUnR1HXk1+nHlaU/h1
mXHUmEf4Iunih5hTRrs0cJaZxvEHpm4PBdUKe9ugrQMOtUfI1TS2wsKLmC8U/g+yeZbcmZcyQ4Cs
0R6HdnOBTl7fh2W2IlV02wV3fNu71yIeRKX8zwoQpz5/dUKlO29WcpRQk3x4gppAuv5tyeRTPMGX
QKhjhLuAjQdZNkdp6HX7qxib2KK65VUWnm5NGb7n2cDrLiKz6WJhSG+G2rfOxn7+1GtLHodRTdVy
DbTfU3OduiNUHHLXmpBeh95Rp5h/2Pteb8VB7pfB4a6JL5V4wux/7kOik0lGc/i6MddxHIjZyuSO
KTxK1AiO69y889qME64mS8/nc6gLcJdoQWMHrKC/a0g6h9H+rO13My5Oqrqjngv3A9UrqRahaANU
s6xqvn7efiKvtaMPkSAVrlyUrVlze9MpHwBrgcEX+UXvSFXJHGTpfuiITFiN32Pjjolk+mL/O+pJ
7zoqKXD6er43s9d6JYFm5WI+l67AEsDyIQQQ/hL4ZsWFMgVF+ecytCa7uVQBs0EfqPk85WO6byrI
oySNJzW6QlXdfJLkIynyI2lf6exLfKZrEbcSLVa1gzRSP1HAuzH/J4Yctr3J2IF2Znm/Njjqv7Ph
dOigiA/yQCT2ttixyIiRPYAdTK/cftmtLrhlcPHZljEU2Fp3gjUY8efY8WvZsmXZlOXd6Ha+Uunk
8fkItoCIGbwwk1+qvRsde2pWCgcKGmZTaqhXX2ZmAbaXVsjF8x1hIAipzyb4tC4Yv6IIsgDYgQ0X
LIPUA5vBtfDbxhTqE6VmgktF0kwzUMS6hL5wccnn1BN9RE6T4lxJuU2XCBqYsl8CCNAAPZBPvodJ
f8pWVdWpTmC9fiKLwyI5TRlGkjePfr8e1XsOvbG7KMNbZ0tTUHPa0yDuLNaZn2VuhbTUKyjaHw1y
xWvN1ZAwXpH0oiy6vx1k8yd9qW1OFPyq1HndIqyWv0VnjlRhFijl9v3rEa5Zftzx57pGarc2/OPa
EM2mfXA0NECZPPZWIhIBQN8yZXX5FMQax61SIALLLL2m+dWkpb4ST3QD5I6RJsTxjv4pCHCIJGMe
g6HrRrybU/59F4hSxSucTCClrPqHM7mn51Fbfw+3MbNG2uExGtLQ4aELQMO909pWUqxrA+FRnTwA
dBKnwxK1/7bzhLgEeY4J0O1fcZ6MWWL0rKC80Qa4DjO5d74DVQQXFhjdaxMaiGCjweO31hH+YTpq
PttuT86kVC6A/8d/aHM+cYGg+L8a7tjYIdu04J92ZlJvEIPPSUd5EdqESiFIEwjoLsSDpBWrghxc
VT4lBqnpkEL1SBwCPtCsb0ADprPiH9SjOfAcc22aH4WvAA9t43NzhI1N5o0I4ncNapkJA0E0hV/v
pWJrYH004o/GQt6ilVJH6ltPuq1r583eS1oIFXDzMnM6WDBsjBh5IootPPLrO5lKo9XDXWzJ8AaT
xmlYSECAF7gNWM/W74haEGzpCEN9xWtXto3U/h+e/p3n4oHDXeatyUVY2DsLXewLIxKhJ644Ufa3
bSFQFJ8zNQNP5p7xlREPQQyl+lW8wklaVjkt/UaWwskfVrdXd3KL0WhWzxOoBc9sloqCZgNRssdt
s+fxVnTKfO+kEKW0w3YK3YU6tAW/V/CBXpJkcfJ5bSjzO26u4CJHUIGFAYfkpHMswn0hRcDfv4UX
/P2rspzCgt4Yk2Jw3LebB3XzL6CCJiH5hTi/q2VkaxmRnG6Vxgks35lhIOAJUAphypzH0F2utHB6
/+KHHRH0MEyRuUq036aIzFf+r+7oMj5TYYBesSiOiOXvdWGRI3S/EZ+J5ACRRQaSEjdFbNXM0aAC
5Ah7ftgXspk010gI/GwiwQ9NDreaaYj2rxeBqIm3AdgVEqSgK4zrG/i1HCb07SoG+nHU/rwS9n+j
SOrBNVJjoc9NiMRa45K4TvEv8BOHfvFnzS9zijGLRI8EI/NRTXq4otiaxEr00gtJGzrxbhLUJNlI
oWPLPp52KPdgDB5IKdNH/9ldJw4+mwI1ll9Krnps2CTHdZfmTSHjlQtkOGqA4OdG3N4iRBhRNi9z
3f8P1BOEei+gfv3eYBrWfWoOPe/pZl9QSXC/aC0qrpJUOkmcEdcr36IkPayWBQCp0WZ1Irvax5uc
Kjvf3jXpK0yJb3LyqS/tpHWxjFlScaf1/95TKyu+pNPMd0wpQGxxfCKB7XA+sX176qzAMloOZ2bX
NFWt4UmN2pphsVdyDp8BUt7SStp5UPzdNHvChiuQA20O3fHaKKyJ7/TsTordMOr7Dy4+y8jBHEji
p3iwlHhMwJ8zKKoJ4ALWj6BBmAgqN9/1TguUE0yVLoDeCV21a1Zwy1V9sQHPd0lzZBODjk6/bXUb
PjLd9D54MOqTPkWTkc8WipczeZOPMZn3UUFqmAyr0H7fOMcNuPZGrn+2xD4RU1vmzJAYyA5ZF/jQ
Z/GZB/1slzOheFgL/CXFWvK/dU+mgevoRHW6O44ecDx5oVFkNefOysz6p5OQ5ZJc3p3VuBFyXBdr
5kaOoARzqqDTHMq39EvVf4wbmQ9MgVMjPxy4bYF4CDCoyzlOKrbUEgrPOsh5peOnN6mPIphBDHEl
2zb8knHKrwfH/tsMkzioDCq3vOHFxi6B7oEyAYFd1co85VBos8j75DOk7Bzja/c/av2KrTzWzyF/
Z1zBP/wJfALlGToy9cvk6FWM2i4d6FQgHqxtdOV8hCJ08FHJaPbaqC5Vg7KumUACi+/zrBcw7pA+
IBSd+NNoSG8IEfQ+XfuD2FltGpjsi2UTBKb5vCjQIKtNyO4qzjX2uV8zwx6e31kZzz+mfaJ5BJVC
5wUJxK4ANkKmNSGif2zx8D1sxrK76CnV89xkxtWs39JX8+gAWr7B3mojTinihwwnD6VvKbJv6Xhp
BO8kNE09QVCIRHQ6t9x0KVvsfjKsgXGBxahLUebBZGMl9JNupZSDgKP67Vx2O/YoisXJTfuTtjZh
UrMefCFz2DcuObIyMa5ZhqFP1r1GL1Spv/6TGL3RBWcQZuaaDx0PhgdmthBfgDpCrR7r6areBXgX
31u8umSHiUsOTV8J2IU5u31SKCghX7NGLNASkN8AmXPQ9Ir3/JZsNIVgiZp+B6nDni0T7GopPLG5
l8CQXlCc7258K25Z3HiUOz/DjRjexFgaBdcG0DUn1+iUpOObUkdeGjLqtJmSBrEKHnZA8UeiSYPm
6PeKv3FhnbxSMziMwl/LMZ9InCkF1Wj4qiAumMKNcHFuX4mZPCHuRnXY0bXL/v55+jI5j9fQdsuD
THccwSY/0jwuF7I6jNBbC3CgqFL9LbSPmEVvov7vEPrW0T6HsJMOgC8EY670e1X0T/zTxFpvEGLm
HOMouJ9PDiCfv+HbZMxMUTLMz6BHr5i32wO5VHDUloH0dCwFRYxhzymM1BLtfurxQgKMn/vqyt80
8dS36WWC6f79iqqXh8RDXbPMcZcBiVGgWrwe7OO1RB3N+kPYsQ1kKu1JkGZiujd21KHGT+1cboYg
gqnVlzoI9e4TFlnmbVPV08hyoU19Fr37Kg5GJcYs73BRDX9r4ymdoUOLU1tVg4lxKl/cFuaQuAuL
mQ/iJMdvN2M1rgGU8MwYdeSFFm+8qkQisp1epiVjiYnaIsrVi/S0E45d5Pt7B5AyYoqY3xQjo+nu
bNMx50BpojMsTWFZEh3It56aBuQ0XuxAeOeUKKcRj6cwFh4g+M4OLukjnoilJK+NgQslQuU4dvHC
dD0N1LlpgRgL0VFuMF62g6j23QXh4np2wC2PQIXtz6JWvApCYJJ9LWu0tYGlD4s6PS3bkwJRks1C
er6yaCbbKYcEmivtIeQPBC2zWyMvTuYo5Th+gmEQd4Qlr9etjMXk6sNSaDzFfXi7FW/9066QoAUD
JY7z/9aqj4WnEGtd8K51UR0x3PJgcERguI5PpmEZvPsCZhPJqB6QTnEblVXGbWLZebCFqv03JNKx
cTP4UzbKOlbW6xbFMSjPUPjP4HiDwIvSgqnTY0dK75oIGK3oFF3aXbdyApavsvwfVjwRfI9rp/al
LIyI0lEmwBuSZqTc1ha33umMTFxFTQ2ABL3k2/7zsS2o+9iek0SDuLC2Jw+6k9zBgD/orO/Xm6T1
bzQhHXRS4dBYveFmj7y6EcLvU37mQDYtpmWioxnnRwuNwUIgYHpwWM4NAGF5RCxq2NHFL9/K4xFq
pfRWah2RuBAIyihmBmbQCBhWh4lFsOF/jL3SNYxNwQCJd3TMtttTRod+gPFKVioIepYmTVXKJbT5
LmzjoBsmdq+U9zP/EyrKpN9tc3QHLx5rv3miw0kQkrJn6tlHKVUbkkHz9G/CidT+kJqzXMKbM01+
yVzg+FaRMxJyKHjsQQvKuUBtij6ZpvPtMDleTJ8Y0tN/yn8+NQ8TFHr6wv07kbsWr3+4RfPsxbRZ
SOES3EPb3yYv40KFVpO9aCrdaEm4Awj4RohHVKs0IsN6iIL1MIprdmQB1HdyBMsUkGh3FjP4ZI5i
zolG6etu5LfpLZcuJ0EE+03wYOXPnapzCD9/xqQCXlpzkiLNhDvD5UnB/5wyVQA0vfleh5xSa4WT
f1e+pId4ViDAQElLrpUxFf7GmrgHqqWN2VBfCGlYLFmRlkLnGwxgnJ7Fz6WgdhVGWMb7PmJSmSpD
EO+0hk3iU9b3WDgC68/jt4SxK3jxIp3MAaEjJ6HGRDWPYU+qrEA1RKw4uom+3O65h6N6y8vgwEh+
Oqe8dyWkCorZuxjJvhIxv2zCLJdCGRqKAfH+CSXUSq+UX2nmLtDY7ZpBO4roJ0yA74VqeQcuW2a2
qeU8nro0FAe0tk7KwClw1ET/Hk5/eoPu3covRGIm7hormAtSG5EA8RBFT0oB8zXgzr78eOMAumm8
NgMN/PiVEf1Nb+qBZ+n7fWJ/Z60ht4OSd3tzl4lwkplRnKCazBt5l9Na3P9Gi6KENSCVHgmeXxM+
+jeWOnClCgrHVYXQYX0YmWEHrK2LccrQvffgITa/8PSMvGlRzpGF4C78e3YNHBlHuOqmW+dUvIxn
MmN8CS21uXlFdNHWouA0dMlcF1FdE3SA6StKIcQBwjIr8hQdssY0kHG4+bANGK9i/B3ErD6C0Sfe
kXvyetKS7GJoADhf1hJ0OsFeOZbh3lgt8bdeqwK3WGtWMtaBJjNxVyDlqFU8W6ls/ewdlcaeUDmZ
bdAqLLbQXF26ZxEeVDL8NTMxuDPbo8EH2SfxCqvx0OfARhibwPnoB8IbuTy5XWTJKx82nsy39x/M
O67Pa85GO6I1Z+RhFCMooZf9D5YWdy83HzCNWSMBVKtaM999P13BoUKgL+XFVVA3QwP2a/eW0fYs
HBJo0NdQW+lhWOoyjKCSqvxN//i2yDVgsmtRfII50Jyf07Yrf8TbhLB9JHl83pLwNQtRTT69Di30
k1j1O4DSRojtXyDVaY0acDzRdINmGvF70egQSMEvtCXM5uxMvC4hY58pkfxRIR4rtlb+iYqro7oQ
wBgf3ixYWIf+Qmv22UHadXidZpTvjrOTxD1W4Ml4WpS36iRA3HVVm/5RcZIE3EPdfOr/PffNI38w
DBLkeGdZPZxJYP5L73iCiFmiRxCwh0+Z2IXls5Iqj5/2A7NHVEbBicPYVWw3KXIQcEHMgvvOi+Ao
o/hnk5y5jno7buJ+JnZHGucD0V329u8V687bhAx6G1wyqyGgz+KSVieKFRHDVMkMTtFwGOGj0Xhc
3/HCK3RgG6rbHvl+Qq4i+nqIrt/uLa6s5pK7HTGY39DIsC6I1pm1Ctityt+O4w9SlQzS55fNMy2m
lbiC9XBRaBpD4qmzYx2xHiRiGB3eCs9PEPgE0xlgUrFdFj7/t0o2MTBYwDcABzdLAyse2CPR91qa
jIJDfQHkivjz5FDxfmfqucI54ZX8uoRafnyWDo7u6mlZC+SpxvpxhGC+5xhhgqVykcRorxlAp7A2
E/F97+7Tv2dxpH2ic6Z8NmqS/3aTIaCf5xUx65elA1ZaUyteGOveRK87sqcyqfy5iwb8EnqaV4Bv
DFMNWeDVD9MfFGVIY0J4ne/ywrhQkeY92tmhwkmDfx8IoYfwqcKhZ/Cj2czlNOzvY7TANBkE2gvQ
tFG3hrBdKiN8KTr4YevXIEjsXYq5+wpQ7xoT0+cA8wzWEbyA75wXWAaez7nCL1bLlVgTqIzNf7dd
88ZgooJY+gvfzG6cVOkRwNYykUAgvfoCIJOKJZFE6C02mA8+2AudgXNxaIcH9MtNoJuovjgACXRH
Z0VXXfxUJGgt7hwLgnOC5AEUMlgteQQOTbLsRAsFQLXO6oCkdwUeOqR6wJY1qWqIr7rsUgo5L8Z4
ZQ2d/f06ENiV+TTqvdnOKAuV0uFp2uDowFGjCEPfGFI4m19LIY9A3I9IoG5BjFSftp12ZbnHOrkr
NhkvX0SIkKVOX1BfcnYC5y+pD2Frk7QMWoe2oKNAsmXN1s/ZL70iW1NP1acbOd8n55ZlJytZ4aB3
xiZp9P6SkFCHRsd/C2TxSuc+qiUbbdqHYPvXt7tTQ5qcxaq646OhughekuJbtNuRjapFpuiE7Wwf
mGvGBT3NY9bSocJSL7iQgk/5KuIx/GpPzHjHymfaJXRBeh3FHdbf4L8r9rZcIqNho5zQ6+2Rr8LJ
DK7MQ+KapdCnYEANwz//7zS8Ts+rCuPG+CgDUlyKC40q8n9m8xrv85voHE/jljZ70yYRPOEJwjv2
F48O/8Q0CptiIN9bFyv6oit6FkvioLSNpE3JVYtrY9i7/YKW992Z+aQjSv8/1aROu6uoNJt07/sp
n2lQ5U+xrsrWynkk+ZtkI3h1O5txNpfHoYHxqf5hCh4psHvGwnfElQnzjnoW4YTvKMOrJNYNGfyD
IIXSvsnmx5BZcPCZ6PWJ2AWJx7QKwSALeyUvrDCUZrXOP3NsYoJYmHxhndwn8eiNd3DCXbPF86Am
HuzISotKXsSGsiPrXp0UCrqd8LWZgbgz24nFWnwR0GKdG71iG9QJhcrnQSYq/eti233b80TosLMN
M/yonT4Gv/MOsWlS0LUCeGaohhxTEXYlEwK+/zUCo4RmO7rVOuoH7Nbdo5zKwHZ/5cb9pLGXfFOb
TkmnH8WxT2NlPF9L7Ara74xPOAoTW276TmRExUlEtrvcI/hcaBzJQUP3oxg9k4hb/F3D2T4HUSJE
1vQ+VGWgKmNDRU2Qsj3FOW7tRM3KY/MqukXq03E/GnmT6qG+jZQIQMq3LZxkRLMR+WUsSjDhVT2z
NgiLs834WT1C6PmkaIbm4BMBxFxJAH7LQFtAQQlLnRv91xgbXomQw3E5x2OdtCEHfAobDGHzMDKY
4t5GAgeVnrRbc+BkeTU2DsADf2eDjMqMVvstNc6jFgUVtzIFX/XDzA+8krSwNl7fRv+tqtfkp53B
fJZNPCvI6Qs05XEacYcVsmZc1bABJLVJDIUgdMRqZSS/+Pqif+wJ2dYYR+U0/CP4vgoUNcySjtRa
v5OO+0YOHetd39Rn4ZDTwmHtLLLhlipKM/Y0DD7J1Y7agv2nhzh/MTYUoBscL970m1PDxDP9BqG0
2+bF57EMoE7iuK5XVNDvr2MSNUZBYResqdlUlaQRbkMThfRZiu51kWk2FGEXkGNB2G6Kvn8EZPCt
lki0Pme4RFpoEkvFyVT5s7IALUzH7TccXJPueddMQ2+VUm4Mia6FKcwK6XycQoSRH8Hlqw9e8TO4
z25t6pgmzpd72v4aUaCqeJBPNWLUdjSeoOowNDKIb0xddd1JS8HDDpoEpCQZZJJakTxVmolPB0EL
JxEBEVBlcBnPtTFOBnxhnIr/ZSNyWR9AfK2eiLpEey7RgD0bpC7bbwoNgHlEG62k9oK1QW47L6tk
F4OSOTEoYtlGue7dl9k0HDZHoGWKbuUnhlWdkcdbujBhxJOzmPTJaR6VpxnUDI2d/5iIbynFu5o9
blS2uw9ZwUFUKh2LHEWp1jACM8pNnOZbveCB5AtLu6Z1LVbAtnRv3Kh/qBocV/PzRQLMjQRAK78m
jsGYBV7v+KKvvBuPViYK1sHLjpdtBQNTuS0k+ONwQadjFySkZ5PGohYYiAz66vEzx+pdfDjFQxuS
SB27nI3fKRBnDlEbsW4Pw2fjDtc3x6OUn5/8QEu/Dv7O3W0yz6CEKKf2WEm8WcylQuDL9v4Um6Fi
p8X6yqNw+tXctueErxw+C5kqwRus187O7OD6R6B5kMKtfHk5imnrdLmydZK45uTRhfZePTbrfTrj
2RT3q7HEraijGE8rrSTjlVfaHWmcDVVllbrol3sjLJSqTCLVOKAEoGXOLQJjXYWWvuDAc2kkTwdS
kALWlI1nCL0C+seSKKkjywUAJF63WDfYmRAfCw/TjYUw9o3K2dmTP7IRoO3Q9hqsRg5VoU49mNJX
nmR0Ptuol2L2AcZBd9N658AntL7NC8EcE6rYHpzyWQ7bu8YntiAiiJrvZQiDAJePBRBq+tUNAvKx
gB1kDGJSQmv1ZDM4WFR1G2vQwZvaE9WNF4cCETLVAQd2+lgKqzg7rmucm+Zk0uuUyjY1ytMt7aYU
OPk/yDI4y6Jm77y0aJ9Adcql8dkh2xCjrFTfzgT5GJzM3yYG5O8bcB545xHjBEW7J7ekKeD9cRns
H4916dA1K54obtx3soPXMVyQVsoOQfyOrCyv+cq3vSxYpKCaU3WUk0rILIH2W0zHebXVqhNI3Gxa
3HKwgf0yiNbTMBSnutjuAW/Z7hS7v6N5RZLxon5XkiRsg+/iAsmH1u891tQBDmIoCAhHo37T8azY
Pv6iKm94zjv3GHV9yXOF+VPP0QTDv63KWEjGp/Qmdx6IA2MnsRYlUGV6tEvPnt0pjyRHHUYc21qO
4zdtFMFrZIJtM+TfZfFj76gGscnzrUwiJsmlE1435bwNbZagud1n9rmfqXn/uEfUOG4LAs5IpHuw
OcBZ2U2E4BT9Dt47iQBElxx+j3t3QoCbtJ8yYoeaR6n4ZtOYIIVa2qusa3CiDkSsFTS1rrX5AQrY
gD49iYd+IRWhqJgzvZ/nS/Tg+k+mEwWITURiSw/ZEuXPxf98SKMIVILjMSA/ejjDT9UcmOaV4d0I
cO8NppXi0pYxI/BA6Ea2Ch+3dP5fPyTh9n4MmCiAp8Gv1x+sdtgsutrq9iFUqbvEVcVBVOKIDiZh
FLXMSTFQgzH5+vDCWOSnbvQo96E9pK1ueN687JWpQe86129wveFXtC3m5fQPH7pH2yyBCviLePEq
mG9FepsPN1MTwRvr5dV4HBMqdlx+N56GvBcx7hK+/YL87GgCFPeidKa5YjQ60iD9h7qjBLIi7fK8
6YxwbCj1ZSQx0+MGT5QNNjHxjFw/ZE0f5HSoZYgIl/hB6MD+QTf5ZVkVZjvz2m4g8ZHyFkVQ7nwA
evApHEuh6VzphziFuHjQRh3NHXp+81dT2663SgDepTliN169V204O4txI6DRKt9d7OHnBlM3Uh6J
cobhm7zluF1wDT2wYNGuOTdrYh8lQI67EZ8OcS9L4aEvmZ5nqtG8kaTc4M+mXL4WE8eIErCcskT/
O+V2JJsl6p1eUKLnKaJncNGhdwZHJIqr6PFpXr3JkcNgc92THD2PhE/7qF4JV3SzurhLn/d9BM89
IK/JTK7cDhRr2rZsCw6utyw4/k3VNn62dotKrNahHUuNyAA9iB5dX71G4xZa7wcCUhHMxRIhqRXh
DTo6DNqXBVGZSIR3oTC2+3aPgMS/CbEoj88ddhJV9sYpfVrOIDtas4+kcG1J8fGKR9DLqikSyLAG
L8t0iZ/lf+qx4KhkV03yubmA51w+sAUT3u2RtrjSU4N6+uLl3tSSYdpDpSTYzRyEUVoQ9Dfa0qXT
B1R1CRZOqXM5bHCkltCiBUc73asDweUoJWa9reHCjhyMPEa9m8YiEiGyGy7cKpCGlkHTgQ/qaGf6
YVESS9yilruibhxSB4UCTK4R+qwhneLt4FPvXMde4DoAIZHuxXUn/2OegmOd8BC5XXYD7j2HWWls
Gtva/4eNkU+he1iBLoSbTWU+GORs3TRaAcx3wIsviN1Zl9NVGyNAylQkHPNgh+NY7AhtEuIGSPwl
Hhzr9wFlGNZ0zst9iz3U44r2Nz8fL33gxARHGtDlSn7H/cPByDV1uCWnoS/f46bEp+t6/1VmEnfb
9GCsN14ScN9DuPACypxmzkhRag5uoFsP3OvKQOwi/aKLk75RMZktTiKhN4v/kPP8F+NNfqBDsvvA
vhBbmz4/sv8oYPPpJGRtqxLivgWzigPEs4pg0hwfz23Z7ijjmc2JjTNz0CQ4lB8FVBhtjdM1bBvA
dRA4SClJB+Bqm1nLGfEgWCPWoREz8kf5WUTS+qBg6iT/rdgImUBjL/sogitYTU37LZ6S2pYS6Fcw
A8D3HvtchFU/rlj+dtBkKVFomECXB+zviyYU+f55QqWwnk5WQ0LBVJ8OKeTP3/LrivDZqkkQk4QR
rcCY5ZYTQy1SmRplBZj1g0FrqD44O7TSTZlNo8MNFv2hhy0SFRxwWupl8bIunYemjE9yGr6E/E4s
SMTXb+oK6KQIj2v42uNW6zzrUzkDwIjprJn8WuuAtK6BCKub2WjjplVxVnl7KKMphpz7MSGCH1JH
Y0QPyCbOqcQZ9uIbnBX7VhFN0mRwi+j7hvJeIjyS6nvAlPEm3Hye+1Msss4Cws/df5Qm6pYVyA3D
ZHnID4sz5UwHCeE7SKRLTttBpOu1AxNhjIMV7qEc+IHx4YAPfC3CioBjTjesSIa7fDhDFC1qmIDZ
WTAS3CFmU9gtEI1vnb6WHYSziEgs5P2z15BxdJe0fRydeYAIDVSDZRUOY+oKSIYYbPzZmB63x/C7
Ja3ND9nQ39zMS/h3LF4U08KOAYD8mkA1b0pEmTuFwxtJrN0Yq4aYZ2tGAEtaLwvge7EKH5lztQlw
CURzWVCylcEhCQNJsF41lnM9qBzy3pPjUtHC+iw5UlBfRZQtq51o4Qt5gz5toiBChUG+ACYOUipv
g3O7IGlulS5cg7GLrA5HfHQ+YB9dyavjjdqtGl7huuZ8/HsDyzeG4PkfU84lD/9uHyDlzW/YE8ME
trKP9bYffqIeQKhrAUV6w25vJaGhfU93DRhfUo4NxZFDe+siM8P30s/lrO474OoFQGEYUYECALRJ
9Z9oNCVb7aW7RoxqdfWWc2mG8xBqg7YXtL5c/HMhrVFiizimMLbsUvctskoDEV8MNtHSGqpDziBI
2+7T4o1SxDziIRYIg9IRanZa5QCoBqO+1LxygqgY3R0zDU4/r+4IlhW8R9YOSINvvEvD1L8DtgzF
p6XRIAwTOY4IqJc/d5cVWq+zL36UA4XQLFsUltoSaZ0U+PJkDG3XaAHPQeJQNGQzeJxvYHfbVbl+
SQwAtKX5gjP0Ph0L7HHHwX9uKB1QsSYNeQPMUPBPWCjv6D9b81sNNju7KDtL/gsEvdIzvNbW44QG
hydTInjyYPgS/zGyowL83ueTUna/ZMBcZeBZGPeCOdxtyA/Z2JMMxO4T8sfmeWYdfp3t2y02Cn0x
H6h5HXpMQ+q0sAqAxS5jqinTw37/O7BtPN8o56JjpL9x64ctbrgjA1KPVXc+flK5DImaAAZ9k1pH
RIjZY+hEYlrOLCWSSBfE5ppsANWd8TZZcwOYs5iy4zE6+uUYnlSrDsftWWvjdo+MbZTErN1dyrvt
aVMptc8nw3+9M6aKxqXMTY+6BpixWN1g3b8zGWGMEtMOEEalxcnZ2W5yfYI9HSq+bfJe/QFJJTnn
Mlk36mvUOVTgFqmrerTN7cxvyZrg1PCxGI5ga45IvWJaA/9cOD3m2PcJ3hkk5O3GCkvGzyenFhQm
Q6tlZC/qAw1PdbKhHyje2sxSM6WpgXsce3WE+OxKxxadwS+Re8pFvY76gTB6dcxZjSAclZpp4DY/
58abxZOu3LPDMz+rSpi/rUeqdhcudahS+rHY5KNGQ+UxqI7nWi2ltE+VxQXyah6KWq7Zk2i7xCqQ
GC39ecoMBLXvcrCu1YBpaUfiiF+wxRpnDcadIcGDRQtmgsyZDdvd2EbBDVs6zxnLQfFxdhXeyE41
57ZabvmtsTKbgqEie0xgFuHOiXFMaJtAnWeqgN709QVTKnncATdJREtTJGBLb6YPiXZCtZj32UVp
1qXBoy2F4mg10qIGE08bATFQjMk4/oMj/iKDWkWza+8k0bMv+qgnGt7xDIc/o/B7QvDADQKtwWEy
22tfTfQqo2UtubdfVJWMhxWArGz4KaSRJNr2/Ud1fYzNi8d+/vjKy56GAog0eOtMD828RBoCba6f
SWcRarzaoCQe4S0+zQcdGffKerprmPsZAWDxszHEb7ZJKw48R6VM3+VDPJBn/66Ic/LgLYcaSJhf
3gvh4ZuLefZ4tKk2kWELcE+kp6Q4yKaUPM/4RWpft5FNNGQBnEQEAy1Zp4C9cIeujdtkQClE+WRT
FKE1oTfpjb2f0VRW8n5vNqOa8v9sONRqd6dgZbe8jBGWHIoFZrm6zCf6H7qRlQQt47vMWEx4T+uI
/jX3PQmLP8OZtq4bhcpbqvTO0N/mBpBA6YfoM2V2lWVvR6JLBDa+DdoeEMKYvY/Ko+LW1Qyz2AXm
pkfowq2KE8h48XbJxiXGE86Y62KyEBypXSDFQCE2EwO1+Fh0O19sQ/eZ9qlJymxijgPbNS22ZODd
rROOIOEIucF/eKC0EOJsbIVxlN8VhZaw1XRwhwl6MJOyfUfgDyHBTMiYfUexmytkF0/jncHfBBFt
8R5yBNHsZSdn8MSsi/4M4rMJv4isYJLdseOLCYe/pcTDV9rC4vfAdA+iyjD2Tt7tj53dGKgFSb92
MObOaR5imxuLlm172I1K7WovmEVDqlbRhaKKehLJtenG0zStyytA7KECOew9mSY1Dhb0fBPy2E0m
XbEJUxtodc1xeA86lKow67sl+0X+blIT6eFDgGXSWjvMkfwXFFNlBs/aTTlvavY6ni657MmeSpNz
9YWAhd6Hq2biNvnwfjv0VjoMY+jDKCj7BTtIvyrkujVuYWQpMdAm1rJzFaPr7Z7UbD5IcGBLNlC5
eppupgiGYmEYjvL9lmaNoG8POUxrdrns6L1os5AQM7LB2EOp2ivRBYPP9xyrsZYBUsDty4oXEjLs
ivn/xmL6nXZkBVSZZUytvSdxw8kBW2RJbPM5Sbz1qfmfTkkGT6TiFzt4BOVHfbsJTW5hfnoTq5Lj
8faQZvqXpGGFfG7htOI6XK5Qgg4novylMvUQflXdXKpogMKzg2GktEKmKV809l5Y0zb1l4Kg96fn
dPIwN2TLBzPNteS3NFeeBKD8fyopwbJ3/w275yTw81Tsvvg8TJ2qGufYJ7aGzw8DU+afQ1KSe7i/
wpeBsV3bcQe25ZM85NUTvBpjPw2MNYhE234cQRm/3UkUGp2gjG+XRaMfhLwM6n72OGsIDuB76s0V
3kaqzPE7ffIRKlHEXHlTo6H9x4inEtVHf5bThbHzI96bEuCUs+IkLQn73Q+uJ+odtivQMuZXjueF
J+X6aHvWWYupEa7stwmGKYcQb6QKgEaknhIicCT+fcTeUhxCY4tZYHM3OJQ/lM6xkW3oYvF5felt
8MByW9TJj8mjPbHrk9hVWZA7ucOmHbT3upPflkicNG8UawE3HvwJ7iolRSKxLWV23DwXkXJbToLy
5+W2e9k8WeRmWQKeAs7uKo2Owmoeez8Gf2u8pjU4JF47gmSE38TcNq7RtjNem17KfrVT+358nCQc
R1a7jHfjZ815/eSOMcDrjIUGd7LnyL0IRoaxnTQkqrJiQPBqbKAXr9wEdLHKysW/+ToSTxGCbGP5
eeUvW+RDlK1mR1GTEDda5+cYWrIgiyhom4yd1ZL+a7y7TJ437NaZjRSMJiX68ZtGjdgCEg8jEPeF
Q/VudPZ11eWdXmU83trKHs8vOo0j5XY3UwEwgTHK7GYpzPM2uQtx+PyHzbhTJLjLgYxCSrj1bdbv
r+iUymCA4He2v8bkwbg1rTZKchwH8L7SjfxAHOK/skcIUioBZlG4tnO/yvRCoGKiru8yMSZBGlm+
Up+5RhcXD/d+7iHzXYKdDP55Qfb9VpiIKAoT8IKbhF/VGfcO8r7xtcY4FljHAYeF6/JE3tlbeIXr
ZeMfl4RbLstMcq6Sn1PjqZvuqUrzSce4hNQ+U9MpAONOqbSA+JU987l2epttXSM6L3i222RaGruY
9c6sujn/xqYcxAGW/ugkf2at9mVsleNwbyxyvl1WMaNTGapD5AkiRZ0KIbYeigfh1lZD9mxYE8Sx
HI4yk/rTzPGEUTrSVF6QH9JUaUDnhFTe5SZ8aTzRz6Tiv/+N59keLMtBXI/gDfJ2tcTUjt+YMV1z
WHEezgodZ7gZpnk89qCIKa+36oPbHIWd1arWNQvnamUDoIFZb0HuSwko4WN5usEL5YI7tArwUzrk
ieJPtpgBB7GzPgV+hvQCKkdxQuk3IMOSyKpaYr9aGsSNImpOdERz4zZkD5Kw9REy3EhLKtgD24Ay
KWB0xrbI93UjFklj9WAuXLX0AF5auejbBBOkW8Hu3f7mqCcahrt2aXuFpWgIQcEH9/pvdnypQcmP
qIZ3AiR84uBEOAxAAFkU+nWXGaJYg8swt/aPZgCdeuYGSC0kY/gvwFw3EF4Tx3YYM7O0gwESJnGn
5wvABeydgHC8k/TMeyn2H8DqCOM1gw9Bar9xB9HO3V/rm5vU4zjCwKklFholyMUltLL2+85Y8XiS
KKpL+CgWY8jGSvxYixxRciSFX623kAKh7zSOLILTT16K7FmCzpEjo1xDSyKoCox5brGjrrnX86c4
mU5Ow6T1K1Nxidr8jHVP7Vxi6ZxwoeP5ykkpiGUHQdj45toUcA3nD+CppiUBhkNtD/NlDq+rUGg7
69d4Na6ffCrC9us2vGbVumKDThvyhT6F9BKIs80zdIwqobjeESXR2lPeekkNMvC0oVcUv7kAgUie
PUXy9jhFPanz4y55GnxeTYk/HPYtcYDhUAnAFP72zc8xD3JwhPeGKXHKic+NNohGOXaLW0b2buc/
ID2yuPG0f6vEqRUM/ON4zlN752xlc7DqzW76nFzzqgkIK6NrEraFw93oIoAmyeIgT3qVLHc/sHSt
qqq+iZm+n++TwRFa5C5d9QBUZD+kTZzsH0TTyRCsyony6+1sOLBjcxOHnelSy5CuFe8ObBsWIkRC
ar8rTQzIIE+CBrhBNhd9xEpDvwJJffWy8PJalbPsrr+9LNcUrhNNRWgyqHL1RFUgCszUlMB16Y8G
1BRZuBzmAzeV52m4BmOq8RJCHzPGiIalN3aVM7+ue1pEOV4/EhGlSAObqo7MUHwJ8LAe+SsdJZ/V
wwPpZNO1JdtEr88XPrK6x5ru0wm/JskoQfjdr4tLqQuL7IPNqwxzrilVETMdHS5gPOYqBgIO2kjI
vzgWRvq2B8ocpxSgXZBKEiyz5CCLRNWIMAKOLFkHNoaBV5BLKhX/BbnsFM9J1Cqs2aIM6Q1f/eHq
3t0LFI1BQNmPNhoCdcQ0NeL22nzwbabm6DMVB6Ri46B1dG4rMZm4A4PxEQuDANAcK9gIjjhU4X8i
kxdzKzU2tyzRv33hEWzvZgIbFVKBnGht+jzYAvgreiO0lGr2JJiFXdgsoHTACvva0ahxoOmAYNa6
NhZ/CVAQ+VqvHKBLv3uVhpuLznLb+kDzy/+hm09pfjWmeRsofqE/Joz9J5zEkfIcHy/k1vQ3FDi/
tFxDdOH8xlaTeuviI+CQX3oenoFym/Dz3ztkmak33Ce9aOuznA2Z4W1x0mV3KWe+XxJ6rQd+W+la
QztxsBgVUmKUelSYrrhDlfzRkKhNvWRLrOPPu0I5UfXFGf6ygN5r+y+CPs6T3ouldmfNylAtOHrQ
/FS4Lx90o8j81RuWwYbp/TRX6qq7eWhxCFMs8TDDFIp0gSUzbb7XJTxePxtK+KU2UIp3E3ev2WY8
B+xHwrARhXjBLlyAZImbkcpttdjQrizTIg689SV/D0vnH8Pqi8XUFC7dDiOYAzUhIPDk0DqXoRru
5jxmwiRXQHGNz4Q5Z82tr/NJVjIp/vc3OTi9iJpU0K5KJPktWLKz8Khul2aYDgtwPoR8nyZzEaMv
WyTFE1MlJoTOTUy6XRuybmKVSHAp20HmjKqGi1bfj6uD1lmqRENtt6SwvJTOxXyH0Y9kP6Xvx9No
zTQPLHE7oizVzLbQPE6q9t1w5A4uO69wNQ94sQEfrM93HywptegFj8dZIyxwRt/oy4hQwnMd6xlU
hcA4RY9oa/0FXIAjS83mQ9bng4KP5j71h1E6m4hd4kJk/iOiF0M1GhCjYJaLK4lPgwmtfxV3xMNk
PWACimHdbZL7WdC1MFP9QWZeXyYrOwAfnFl+zWquRCYTuTt5nY8rox0dvqxPu7RN9PPJJv938cYU
u6gZLWUkB6T6+rbpxHHQceY4eqZD4o2ZQDY6i16whisjgQ67LP371WqgPcB1+ADAv4n9aHrBhWrE
ncizoJX8BF1owuouYiyFHeQGvtbxeISAuCq2xLCJ87+2dFaavwueacdqiGiGymk6mxQLjQQMwhvs
nYYwXkrRKFzhIUQumjCHhIlfeFc2P7jaa8hbvo08VEuIrgga46PtJbrC4gJAHAWDQbWuPh3AnSSI
7bwM9MgJVKF6LLODWbxbw3jerN2NFpgtk0ZGaIVWM+D1vmYiqgyDgssnE0SISGGA2Ccpfb4NywxS
Ik5OG8G1wlQPuzRUC5KAHvWE6PHaXRrJZV7GAM4crEt0/X5HjM1szIj6ymfMOVnkpRdeoi0Tmh6Y
e8vesD4MwX38rmU0GaKFiX2aU4hbCr3nUXXeKrEv0W6N//HmIUyLpikmNWOU69Gloni++b/CJI8O
NgezuUjS05Z6LrA/yTFAkJxQr3WZavFOQVGO79sslUh43Ihr66/2oPlD632P/KnypQ9aHppBhlmK
d32WELnpGp0cxJl2CctsOCtYxmd+MEgz8KU9wDju+Y+QWBwrZa7bLhRcFg+y2L7nOMESdFgkY/W+
dE8XLSU2Oq1zg463HulbH4pj6Tipx2SMTW8+7xFT1G9G/h+rgUuCMusEAySGLj9dx/skQYX57+4u
wEwxeNdO1IffYxteB+qIQVTWwL8Iyu5IaNyc70Dirfs4SvVil3+GTDaOM+4rIDSbue8I9WaLFdWV
dsp54ZFW2ALQ78u0/XF9dI69m2CZVBdldYzTod2v0C1ainWirhCtCLxQvYdOjCNwVbjIRZ+i763T
2EYhxffJbB1kXJclOSykjm5jRKbIWzToMEF1MPwzx0RErAh6zV/XKJ/SZkLVxT4Lu1cF06LxRSWM
9LZ2rZ0ZcGpffCxZ9YTitfgeK2kPQvbfNeI8zD9vueGzCccn3nqk1NQQwBpfyVl1KBzvX/tBbkT8
SxpouJQWxT+T0DG4R+D2rSjBppIi8tgj5p8yC1+/TJfgVMP34e03YH92pgRZpRk2sxpYtSRZeIUM
goi10U7MAok9eMIwIN1X0r5UQA1qgsWr5oZdEau/qyYsUFvyfWuHmAvei2eBhKgn0tNpTXmgO03M
FS0dpQ1PWvrkPaVZpnlymKhiNyziMJ8kZ8Di3zwQDRpSkQVkY+GLYE3CtOJopZFHNJeC3lLSjJbB
02AmJ/MSq9Fst/D1rNHegTpJgP+IULYK7ba5OTD2fiK+9LsaDznzgFg7Z+hw4RFvYnwWoSrtChSm
wiX4dihPsE7+syauBrKN9A/kvq02FASnRy8gUUOxAqLLDSew7ky/897S0i1dvYsLZW8j/VwxIGZn
bJNVrxN0NRguCJzxQO6JhWSo7BoeZm0M2jOt73dtHxCiOtGHNzzOTq6YVxnR/rZZTBC73PXTE8CR
bzpIX4CAaFcKyIxMAfYHqz97EMe4tz60CsxNwuSiIgTAFmGC0nTChCBrb2fjBNXV1YeLKkleKKMj
hqEalguueMncNKouLAl9iZ0GCuGrzqI5CwwA1KB/4y7t8Ggj6sZWtWNXC/NAy8oC+oiqrNuarc9b
VkZiyAt14W/xUedx7Kq6L4eXbMwJFNI5pqZe8DLKFybE+0h//6jWxhelfsZ4zxQ9FuW7F1llXOLe
M2SIY2iEIaPid2Zjohe6j6JJ43DplChxLyHzXxP1jt0iFbCfI+TfoYEbqcox3TczBGx+1Sf4MCQr
CNvGjT0vleNHqfV5ivTKVwtVuC29tMH9SiXDgGOCcK2yGjtCcWnvOiXU3nLhw/ey1gVNSQU3NUum
FWtSglBdDMWV2rB6n/H2honWXjiZTxltCPQZQ1/vF28ZIO/oFjZfqrYT4/uka/cj//4FqjeOSIQE
6hFtsGaIE4kzQtR7nAms2WS1l9vx9FfRTaZGdqjhYC+TZEScMz9lmzyH9lzSKmACDbghWIFOeI2V
6W+Dkex0GglxOAVxeQ3YNWDDcJInUNmUkhgSbW5MEESwX6iGwz95OoDBqjpI7a8RMe542P/NDXAv
d8tQzPpAxPUSdOryBBDehWTCevX+q/vc9Jl1slxrAVfAr+SV7P6HmL5NFOBZf/7qfBfkmEpacDwb
5QirOP5YpwrD8OfrUfC/ITQQmoIXoUQJP1751xIY7KQaoeL+tBc1enYbQnQ0/MIG8GTAB0+07XSo
M004WM6esYNnYUv4crWDdIpymh4i/BVI7e7Ph8G2sDbUEAneicK7iVxGogN31RvrQoEqMzegrR9Q
xGcO5dUN65D1ZeHWK1qMP3ezzR+JhZOH7WAW1FgCeDLfag6+teNi4wvMRABQvGNVJpNlTYvoPLYK
RoQIpZ3J0BHXzPCpQ8qhph8X9S5xTggseF3NipV7NcEAZaPx6bRFnddCIEZHotgJDzDh/OYluQ78
9Xlp/0NtVKtMuzqIy0K/LK5hh3wsrPQ5hX0W2Lxr7JvCp+oXER6LSIcEojqeVOsqCSHBo3nJANip
L1/5QBSsSvXkKO8o13JiRkImk9+7i5I8oTyerMhg86dkKLvD3iMzULhv1Ck8GLXsKsROk2O3LP57
Jbx2oRjPLzC8wx9bxoTDiUhpX+IWbScQyXTERpUxOgv5iK/FS0dPGx+vutXFBKRFFBtD2h4PGOIX
mom4XwLPgR6CdOaWeud+oCaMQSN92djZV5ksNjtXzxBTtcbZPQzWuuDnDXNximDWaljahz/3QpqV
HgZRVHCVGS4jvJz7JxpGuBLLpT2Eg6cLY7SmJ+2DmrEHmtue8YY9GC9b+XJoy1D8U45lnEjVzUss
ueQ8PfmtzlDGnrsCHZLXZjSZgA98pYVUbatG6/k8W9UXpuYz3vtpEovMgY/06KpXMZpc1jf7+uTY
wezv5w8NWgPZTYbgZN52tRGeBQRSnHXKv5FXq9bLKbMD2ubkvmY0c1tLNal8G44Ioh/Oo1Rxm4S5
AMliJv4l2+6xSyiReljT4Ibs9Bm9j1yM6xQjRJyzqW2melQxt5wf9pqRrHl+pn8UjW+UMFGoiL00
l3qroMsk5AeFe+V33NtiMvTsGyDMwv7m/Bte5rLEvIxqbYSjvor+kJmT2SnVwOLhfh5cRUjS/YrS
mzpmIIlISFXy0Wq0fEUIjuYViBOCKju9IgpMmMEaq6bd4cylnfcgJ9vBdgmHPTw55Lho3pZTQc85
HiylROjrTpct8fphr6EXCVdUqggoklk4MuTYICBu6CutM27k4T2NYsv0FBSTKf8/ZQ3TX5QzFfM8
7JOWBpdMNyx1kutUx+QZ3gCQVpbUXPt6AuhS/81irbpKRgdfWF77S35WIrfRYrVwwVAzHAHE2bub
BDA5m2y/viCPEDnmVaK8DMnjY0T1EmiPpk/JcQFrObOBS2W/2cTfEXSEt5m7ccjs9UepTV2NoPN3
1KXM/gyGYnXKitlldaQlnQ6VaYGvcPSJSL4xlCJVgmrhfsTOPE0m8gmmzSt76oVWaKd7kK+Ifm3u
qai5ZD/gNYQWTzwMiVa10j5fB7t7qKcJhub8lamBzQuOEQdo45x5s6PmWxFPyPLYRQZt+HKF3RxP
mLXIupC1AmbIyAloaJz4MkP+QwMUoBgGIdmDpBxQUeJNBkrnNIVp87wOHVxhBjkgyq+jXfGMfSyD
mC+ioB5btyCzLbsMfmkDABr0Wnt4M6etRqLIkM7zZ3DtH8D+c+4qewS/ENFV9eHGglFpIA8OJDqa
P8HHXSFmCBn83sJHzMXeB/SjBWRsMh4NaVqzFlmShDwwbiN+EWsCgI49c7bZ+GLAd3rrL2NDO8X+
dzE+vJnbTVFhL96c68aH28NlknMZkk2jVi9T1/Os4/54LIKNCd1q9pKBgRUq4ZUZngy7jsry7j/B
UBPsoIOVCYLs/pjYMAlwG9YaMvpW2wtvK922HRmDyUpMcrit9R7WBfnvexuO8TOYPXMs6UbZhmK6
IQMrpvheB3S9/sngNGt4mHlFV/nPoPjs3HpmYhKRoLHatD14jfg3hc9zjK760rruyWbpRkeHAOda
VVlh1zfEjLBjvokFvwIda0saR5uoCG4qHUkN9slDAA+4DKHhfjZ3Gg4cLWU2d1CyC4VrOjGCUIX8
IUqfL6M5AhivL1b7cZtO+rCRsMSlK5JfDtRmPFAz3hudLa7jKogJl3vDqWSx6TPfDfPsiFE3XJPI
YIuVnhhlHLNIJ+I0JYd26njfdoI68qdyEw2BIlTDAYjSwSq5Hy4AV1Cjk/0yJ37SXh1VzILmaLUr
ror2mpPTjsgZpEARFkiGY71OrvfOn/Gi120DwHi47oL5VO2EzOlYwuY+R3Xsx20yiJRK63NKzftW
SgdjflWwDRdUiKBco/sTaySB5WZWWS/7qp0IamDd1TyEcbKqtzEKELG2n1LWGaDvFGCYgcqc2Eq/
JMH42oxM1L5fgDGj6jn95NbgiAVaLzMj6cykzoqmjzz5RaMgie98NQB3QVsCcwIyA7jw8ZXgIg/O
eU6Oq8UrXNH2iuCyAP4FGk3CNlmwqPrAu3pp/mPBq6/+i6gKbV1zKi9OA27ewEgBa+y0RNU1d4Ke
PeDCRaERas5KBSc3M/T/B5gMZ0tD0NvfnvN1cXaAnaw9tUog+jk3TgDZWd4GRIq4XnKzBrFJHuwI
VuwaPhov84nvLnNDJklIfeJNBEJAsrFwmBmB/kowP51PCnbkItHCgsm6xLSvHJHKs/dOYTW/Lj63
1K1jpDSUhKXwxDNVFQs6YtcaTmEZ5a5uL0OM1OFutg8Xuozoh7wovPTyZGdy3hXpn+2Vz5R/xN3f
bT2ClK1dO0T1OyI8NqBEpVm4yi1boJ3UYI+G1amwBGOUyltDG8Z5fwWqdRab/yorE0bq4vhKcL2b
eg7hqQvnSvnwPF9KTy+qR7cU1asPpesFvbL5GnjccPu4LOaF1cAh+3o9wYCY6LIicVQaDDwn++5/
LEM6cyHCZuOTlTxPdGIkkMeXYU7HnTPWsa71ABbvgp+QJqQvX8Nts5hcoXLiXGXTXW0NqBUs/Ng7
FTEaY8fjCPVB8uZagzSxbY3vF1GjId+Hc2Lwhc60DE3s9lde8K8oylKZy7z/FED+1h98sj6ppQpu
D6OdB+YzwkiLVa76gP/aKIQ4t4T991y6vGms9XphHi+KwbvvJPXex24KWNszy0flp2LvL6z8O5zo
NPouxP6hdt88Grpv1NnCrZRP2m6W5AbyxBg3AutxSAxoCApcJSfLRVX//UreXro53ybfVYqJvK7A
sqhRx129nfX/9MeCX05tMxpZ/KFJOFNynYkMequ2aXRSutucnnGLAbZvfmyF/a5LMvYrSx1dI8Os
Xy96SeA94sBk5lK3LYdSHFrb/Oe5q4s//8iDppfmt/vM2uugCv+DniXCG67s6zOIFduSodXE0X+5
5zqjDRBWfXdS8K5KdI25Ck6P5bUUifxZAS+Fg0HfheXyJSwJF8/eBuvBwXtsxwNRXYMH7U6ECpmA
PqghzP+HK17XEEBpHLWzcKer1jGPmv2g5mLM2vbaqNjmxwuYZQY43hvCeT0u4pdVxG5fs2+SGm6j
3VtfappqZoDlKdTnSAQEr0wotseZ/seaMMs25TyyYAnwf5UncBMFpvlsx2yRBg7Jef7bzTpByrSv
adX8BAHaIqrMr1ZSKbQaP5SXIcDcF+AbTfQNSb0ZviDXbGDmTFswq0RLWszM7crrYc++t0S3kkBX
5JcYK07mACaIGfFqP8excOp9r4fDMVeyxRV0fB9Y6DlFz7U86qDzpCa92sO3+eGo9O3r9Glrj1O5
4bOe5RoWbkP/vYZAwkEZQDh2CV4W6Zigk6u3Ehcf4oozhxbpHJvYPSLicQrLov/P+kEDWYnMizfJ
7YEFemAgL0CsDJxnGMrxiOPWg7uvb9ZQx7QjtpAejmM/KxMUiis8eQdDcREnbt79cyZj/S5M38lM
7h1lQ0oK5fDlt3eQkCfDcjMAzBuYh4KcPWwiJpN0PzHu9tywB2qB3aYwX0lJSKef7MolxHbwe1Ok
aafNojW+UG+IqCFjOJOuD4d25OaRUTGnkEdElwcsKGVwsFtfp3KeN3CRddlpV5utAbuYTzER6mEN
y038XbrJyDnFQ9js+uXEbIKtQAWnoQcNO3dXXi/LpPM+gQBFY6U4cSBrcczIXwZ9nhyGK7Oqs9pu
DdYbJ5gU+A0N3nihgCsC7dXcoaw9hb15ulPc2K7nAzV1pixqUggc4PCziH9ydWa1qWAOsa1uVc/Y
BecJ5V+LTqK+/k2y/f8WSNfncI2la2BEI5XF8mpvl/VJREUBpBoRixx2PseuXWG7hz1ZBL2lVrCr
BP62Fc25oxKFRxT21EOnExfKmIQDHfj6EViqpeLUqsShGkzYX0ujfu2pNYaSODhnrGqTvCy32rOt
hfodQQMAEx3zFZVO0InQ4TdlQCbP6QGwTq8JD2FJfA4gh7AOlKo8JV2k6IoofJyw8nrYC4/DKQZy
8gM8/quP8IeJDlzMeaovSrbBwTSt1sA+b0xjxhxP4YEmDoam5gSLeATIApQhoKgCzDUMUSfeH4U3
eoDm2sr+ooI+a9f8kBhooASa4XNKR3qyYGBdR2XNR9o9us2qkWZpslPkgA/OUyUQaM5ks6D4tDLV
faP9UgNPDzIi0w5xG5zSS3HoZk/yyplh1GLWBPLSCT0RlxaI7dmpRcTrW/+HPBegQ5pcL0qH55Mv
hFuhGVSlfDpaSULmnJfduiMq4dHzy5Iyx6z5BE8BLvj76elgNp3HsvYaaibirhuriI1MFOSoeDJP
TNQqPqadhuDHjHgqUNt7VLiiQP6Zs8fvxKQZ7wGYXAQNXiQbLCKJhjzCkodg2iT4GpKUkTm1z4OM
9VU/f4u729SxK0uQ7AuQVyLOcZysMWHILukov0REULiT640Qc3KlNQXmoZPDK0iuEcn1gVtPQI8B
2D1iaVCkLybryC2zSFTzRTe66a0JGt/uuOc6cKBUHe5SvOza7Lv3dR8/fVOAT9UHUTZn4MT9GxvS
v71X3uzDAcof1U1IlVfVYOC30ZmPVDgpaloL9FeUx9qz5nWJl7Nod9pSd4HqhhESldGBIhcFKPmF
1hoPYiP23LGJjytRSLBx1V2svaepZCyrp8hjB3OMpvtcnTDjBWBYdfnyZF75+djHdh6IPOpvdSkI
NIuksb6M+Vi0trkBo2k6y/1skqcOIOk0mK2oavdJje4WBlaYMN7pBI0trCY5uAQ4EFv6VSo0umdf
O1dxMmvmWaQbi0043jVFeAHGBEB/FSuAqN9SA5nnyMtsYwpRmOIbn9M0T3lMVVsLo2eyUvoczyX3
tv5NpUOJBbCahwOCIiOXIgUQCHs3EYy0SBUzcuWmIONkQEN3XLIJtH29PEjv0MP67noMkEUjSgI6
7APoY0M5hFEop1iGe8fk55EJQXPwx/Cb4pemVWcLc4qyw3uhCq5npxB9o6TbikubqiJTs8G+wvmV
/yjWRE0k2X0Op6DeCzjoiLF38j3yQSVxarrdDiDkdLua/wlcrTA3mTIW0EJfZElDn0ghuPwDDWO6
b+VocaovUnEhvg9+J/F4hQIZqc5W/ABZROEY7ZLsVkxMEsWX8Cz39up2mhktwkaKkuWB3TEGMWhb
hOS2bDNZhuk9HFmZzm/ak3ThbkoGlC/Ahvb7hd6uoE9bNcjHMz2M4FCvjNIlF3C6g64+JbP28D5j
OXh1FQPgd3A2gjfB6FbSKCQ3i9SoWSFAdJ/yrY5Mt23pCcwttNH4R6XlXtX8LBRaY6MfbPGrXC6t
CNfIdOACFx4vVp4n0s41PavRDcxYn1skGCy2ZNsAjY3Z6AI69mo7NV1NKxmlj6lfscxgCVjjEBwq
bi6ciF6mVlM8WtGADwilr7Na6zYrpUDpuz9iu1fSv0EWXNjKLqHUftUxbWFWbI+nkSYx0wI1018M
ShrVVLfBxghZlhyWX7UUR6h4re6mifWs+LvoZKgZB/soWO3nQoYLEsAYz2nqf81XsMc6whCn0G+c
zMgzTt2rt7tsJeHG86xrrsZcetO5EvkxZpKBA3iYRcColCl9O+vxPWkQ45rM7qxAMmqrTnMVr9du
TYVw5STyeGHXtOfxy8bs1y5bK/csbyI3781y1+sfU1sKHSslmlUVN0pXGHPVRbpZR9oBf6aSWwFa
eWeda9yuLllS6MyFPGntdvWIJG2iA1UJHaBQ5xf2k7awqk85pooUM+Bwu7dADnyFRIQmSrLDj76t
JMWNnFNavLaTH6oA8ypeuJITmkiWhKrGUWhYyjtGeLZfQ3TFlbCWyucyItsd2V5ZDAlQ7DiFwOAZ
waUPANg7IFg96kGauu976Rp9AZxurznhDWaKE//EDPFG7Nwlu5hUPpsI0L8aMBWyen3Lg4A+A/1z
XvMKvrLWWrODhuhUc6Qf/N6aCo7b5Afkg0uNf+N2011mOy9qfiDfbVR0HySI6bu+OkknphNNxoXB
HmuCbnwsWdhz6tlBg8YvsCJE/HkLovuPpQwE+MwLUPbdtyYfF9PL/P/HiTMEfOIoW4YVaTYkNKZo
Br2cndgx9BXeglol75fAlW6ir/uq1kcYJsfbo2xvhUKZ925t8RSvU2AH1Sia1SoV3RQY+ZgGbO/v
tMbc/jLadEHqa0FB4IA8lfhKKYfPMRvMYxJgG0CqizEcjnqA8XJkFQJeEr+PdCbwyQIChSei3LID
5sLK3OU8feCKm968XOQz6kmUYgflednpoqnwmZlBOJ1n64x3fBdsWiPwZYW6NlW/6vML+ShrLb6v
v//aIGvgLcgzaPpZfZ6KDN4LY26FHwEYt3i9Ri3nA66arxkl88xgsv9CdtpeLd/Rs+GR7Y9/s93N
sjb3hOLGHgORRU95USwmn0NTuXeiCPwdKCED6/C37nBV7Tom2S6hLpF82Er4N0VHXdX454X0EYh+
cgj+D0AcU584xMiA13hKdd60irDmRGmdnuGon6auaMtT0dES8qyirqHdhWMpVginCultBVcvoT4f
OFh4hUzjT3Q0zqRJ7ppM0+1W66u0j9WgVVi8b1/pip6c1j6ElCOALqM/xZkShPiBwkPCf4HeEhzA
9X8NkTOk33WsZxYRMhsudLhnjB7GfM9L9eZYQnEivc9HTffsnBrwZd7ouy6o3HI8RoPOgfc59Khu
kOaIrbMF8bRQoYqdoJijb0Z5866UKtzyKnd8+4FltoFTatt7/fKEwgkITQj1OJVbWAnRi+ufx+RU
HuHMQv5ZA3NGGz1od767EJvOjlt7BE6fSLEb7t7/PRWTRjKvf705uv3zuKZP5Vo+jdItl3o6SV4f
9ioMVfu/c7J4bx0TtTVqXrBFTGRm8gczeZg6+jDZlFLf0FGtUBlPK/HgOyKCweTTjOZo8W66iVCi
M1rloOoy4rNM82BZcTncUaMSFjfY7g3J8kzBrcJLR9GjxCaq7AMVZRJaLigMdqiyU6ZsWhl670o6
Hfmg9TB+29/BPMR2Akes3mIQk3RNeOENamNWD/wuq5+KZJaN5s8PzYAREsU/kCs1UYAk2A3dn+1A
s6UxKCQGpDZ52Ngiz+65ALSWUlSHm7S/uGdSaAZsdSU33ZNYVzgu6xLipOoWpwhuZayipjFyKD2r
pqSuFE5Yzq98pTQyDGeZV66NDqFDzcrg6vW86U4G64pH2+FP5zd2JZ1CbYImADQx3FsP9/l1f+Ta
f6var9SyJ+JvwbLKCdPYx2prdD3kBktcD0hojnhvRtuVWLbN61paBM53Xv+8F8RdnZJxKwcno8DZ
CCC+DYFxqU6xfUq0oLu3XrlTtkHAeT5lCPgyv4UFHLDyD5nF/37IfmyH22EcQ6c/DPIYj3hoHlmq
lz+L0GBkyn+NlHLhXaAKSP9/n3cJ6O5WtBG5cT6yPEPEX0MuU+z1nuTy+Ou7FClKFM2uNV7KNmSs
dkmYujy8P3u7HG73ZJKm5aDP/CsJ4eBZHWaBa59ZMHS1t8XzgS6o2V3nLi3mJu/xwAWXyJMu74mI
cPstFbD8QJwrsQ7sAO2dcI1UkBUfQ50qeMK3yhwHSiZ4HC39pJuGV3aUCMkrazlNoFuz/SC4Xxxk
GinFT4sW0JH4zmrLQV7WwmJo/GBq0JnRzJYZAI31468lMGCteizlGLUPg3jHKCU/84HqCBLXnItO
TL59KZ/NYxtn51oN3wGMX3CL/wlRxgRCrvSpdL7L7DKE3mc5ojUbYIxlIKRN0SyQY+mN+2vmLuVr
u9wrfKMC7HwVbdflKGiV7jTbTzB8zEAUxA+jjX9OE4ly7mUwRIuX8WeMAenFPOWhnqSfplIdEkFu
rsWLa4kmxlC8aDRtg3/VyjkiQe1YD3Li0qwGZ6IC0xOWIgeyIgtP7D5f9aie7XcLnISVBeMGgODx
ntan7z7ATIqTwskL89IQzpkw5kuwmWwErEI21PH6Eqb4v8Vr1W0XVJFz00G14FXM8flSKye+4t9U
oqFOTU46BJ71uRkwclrjfW2ORWizC2yNwQAU37DdSl+CEmfLF8p4weCbLaZ6hKeneCV3Z11R9mKy
OIQ8ltYJB5UpTdyR9Knm9wZrBKEzUyYIA5QX7mn2hurt7e4scHWQfau/b1hqcULU46UFCU+41Hns
syyIrdovgdP14Dt5ozN/oPDm7IW++k0htSnvjxdY6LDuxUW6PmDjR07QQuF1y9Nvban+vBCpeatc
ClwxtFMTfKCy1W1WyxHTM/9Yg0K37lwBhIAecPQ/TquDcbsn7UYqxeDSS/c9tYGccOPe9Mv4+mdI
Y4iHkEE0eSuEsrKDVMJiCL39UThnE/dU02ckFo/bEewWlmgbhl8E3bHXpgWDqkb0jNMjX27gNVnU
R9UKH6G/Q5rA1RN26YXN+RG74kd44Qu6dMXIi3Gzt5otwgBh9mmHxGVv4UgLhRwwu+IBw5M5fVae
wgMD5g656QtZlGmN5iQJ/cvvtoTJ9St85m4sMzu+7f2GUFdb/+YVJ2DYsNnjMgdW4/Lk1RBDmqy2
dqNf0bRPuaCE00OHSm3HE5D5s2/Oqlz5c0AmVZpMrRfZwO4n9CzghoMh9nFddOf7nkMelxGvRo6c
By+li23bjAWsh0TcV3DKtYR5sIhzm7MC1zXfCJiyh2Y5EFMXI43KTHrGps+34OpsD5CyhAdW+eQ/
qdtmCqr1ByPj3LrO44zhj53vexXGrvmdhQEPHxXdwmEZcmDKVUnSwuwIHuwpNnsReSPxtmdulrQb
XSOfJ41Jm5OdaZ1n7QdoSHQkp+olwqYNzKbEQKsaMKqatou+T0Rh/M+zsxy+52o6udrubxJEaS1e
4tfyQhEfYHRBPvM1Fm3TfQmAF15s5JtSXy18X4/b01ppnXQmm8RYCsKqIyua+3VmUaPGtmr06qad
GvjMU7GkOhVllhtRpxoa7OC1dCXdqLNpgcoe77DdzVbsAPyxVYV1fVxnWs8vzlgXHBcEVYgbm+2n
JIOp4a0f9EaonJe0OH4IEklW+Hb7AZQ8WMOyb+UpqPTM4bHXNX8yveApIPUz1km4TDtkb4REI34e
ulCfIYk+FhONQqXraCfE3wcGP5KDEpkYTop9u9lXgDCe7uG5CzsSEssFW8F72Fo25nwr8Ai8OQMs
5AzuLQjRaYqnCWLOPIqpiLPPhJG8b91suLXv74oUwyjzQwd6UGdDBAJ/FFXV/IUTQ/2xVU0Q7470
n6h1p07G/5eTzqrhB+DUIYRgEbcBh3b0ouo5IftJFoFaSu/xTFkLvEYWq7wu0NB87gH3KAZQZb/p
G+sey8mOfMi3TkJFfSnWgdU2IsHAh5Dk0uEPSbwooxxMNtbfAfX7Jc8sMnCJSM7PZfUXXKgEFN1v
08Ga6o9Whj7kI498zkvBjhV2s+sdh3R4oxsr5Wvi3drlrzpL612H7mGS9ccCxemcoJW1fJTrQxQN
X3/FnlrQV4WzRfo7xJ2mCQcuBrdeJJtOJxw5tk4fLmPYgNa6TgBkgW4fwT37FLWshY/1d2otge3U
MSiCX2dA/UFjEj1g+rGtTMtQuuNo4HwTCDYXlrI7hG3DXNbP/WrnpE5fNi80KS1FD99s24VO295s
E5/iQjM5edx70/hjxv9JbX1ibCM6mRzdyVT4GjyAFG+JDu/rLgCMX8mhFx/bw/ra0/wcjA2/VjkA
wEFr3U1IzFXgQh/+u1fd/u5M/5SYXCiylkaGdsqAqgYTvzO5z13OyGnVHPCQnZtsu3BOBNfg3Wjg
wHHYc7zCCOr1PcH6M2rUFUsnN4cb7xM4/WPKqga0EnB7LXx6iCsVUDP/EIT+ExXAz02Th4xxTjul
9lVvgLYz0j2dNLpaEWAFpBmQG2gXlPx5eSAYio0teNeFQUP0xvdJr86XgM+cX21qQ0LN3b4NZK3u
I++E7WyWYrOfJXcu8w38nEmTrEaC9SXEMHUk4A7kFWf0a1vDjLLv8lhHFuEV+8p+tTT/bSB3bdLM
ikRtYPUD/bFWx06BiI4E9daBfXVJY+8rNeYRL9ahskm0lZ7x+HE63hV9NSoCopoc/9s8GSJbANYQ
MFw8s6rHWEHxHkI67zsk3amw0EImW58dRQYSA3l2a+F+hVqX3DWenZrOal0eglVvyw0PIinphm3v
woqSm+r1p2t3r8KmTreODMyrEqrI8KJFze5qUm3pvCjLgxmQDmBP7FrLIxEI1ZMYg8leMF0I4IXK
QuOQPX1G5FYJca2n2EmO85sytx4VNQtawG2OXZXYOSITL1u0SeJUv9VJr1CRZvvt0EVrUFH3r0Sv
2ubszBgj+YvEZLcQzJTh/47N0zRTHUA1MJzrqiw8xPtRunl/trjVzsY73/guXZdfVAo1Q2kBFLA6
cT3pVwLoMj04Tivz//0ifFUXd0WphNCWqPhp4wt+k6feKkg418lEuCKjXDODtDN892hYIUeIH1Ym
Iyao4jWoC7nSAeKKmAtn3nZBC7HO/VGrUuxoFPVVJ5/E+prEIwOMsldmDpJGT6zolGP2p/phoqcs
bOUs/F85zUWxcz1sD57nCbRl5LiCHNDjAWC/9yEPrmAGiZCeOdIrCSUJsjI7SdvcL5+ppYa3AX74
WQNkJ2JQFqRW9TlSQo7q5i0eAFWNHkhEZigbxEnLUjiYn0wLLRJTBpkMweKVItq0g87bnhTy3THP
TXAgt5pqLIxdOzk6SDD+26faUgP5GC6HKTnomPU6yzjkUmBq4u60zZC6t5Unbv95cc2UYvZ8LR7I
/NZfoezm1kdsoEZidRJbqSdQme4xhfi7ENTu97DPDTmbXITy0gNTlvQcuv5aFcHEcSJ3+eCpKrq0
HP2KVKmCpUvAYh7ku74AaG0ylZyk4bvZRx9AvzgBZLlBLrwj9CiRZqFeIsYUUNueW8UG77B+5pOv
eWZyWD3kY7B00ycAlDzLko9U9dzWwWJkmuVOtiax/oN5dUaAfFc6VPWrIaT9vxqI0F6j9qmTu/aR
3yH3rJqPk/LvaQRU93mQjofStC+zZy0vNAXYoDnfB2O8rs0J53gf0wxvlBLbHvH3nEyjyuXxSnNw
NLS2bIFI+4YUZLjaon6KkSXrXalQLBy8/Y9glYUsd6PSf6BpE1klXutqCqurQt0CluDSTlmaYQBu
UB01ibUL78ZrtWdfwpQ/jun7CtLj6HL1DcCeZmXA9d+b41YFu9tgy7p6zQBelmE8pvDu2avazgwL
SF+8woDg9aTgcLyH43VHRPlM8e9pptLyYWQ/vh4VA/Gn92Qi5Cb2L6809Jk5LkRi13Rabr6xMsW6
h2oCzZ0sCPesKSd1l2PEFe12dK9E6chsIJH4mhqzFX23oYgVj+2OvqrrJRPhqNBZ1aqF7aNlH+on
V3RsY1vn6Loy3K9qb5SuaO4H2cZg25+4uuXf/ydLKh8AUE4WXT0VQ74gmk92U2g1rymA7e9ANtBx
7WFYLT773BDmW+wd87kuX+3GIHx861SUn/j8HEs+GeEuRpNYIJjew24sSwB2ykrFxEYpk7btBBx7
BfDVkN9mo6sLkpGcKkxi1SrjrbEWMjTiblJluZgg6KaU8MUUVtpbFv+RMfJkhcT3M8f0OND2FMby
RKRZCwn+9AR4600H6o1QcxbGd47Fbf06QUCKuovVk/aDra9qDXAksvNpyXzAAXfAZ46pG/rZHJRZ
3Kv4JOQqN0/1VVXBerCUC1DhRW4BWZNl/dIRwvDIfoGYRwe7I5yfboNHjWTarCqnBGuWhlnAlICC
rzPHdLsDlAP1PTnhXT0G+qvMkslW/2KKVPya4RnoAhek5noBVvKiZhtNSqv2dm+i4hnZOioWnYPV
H3aMgbyKRm9n+3msF/FmE1EvpQf+FWmqLxUQHq1k6psyqfBaJZ9r3zEBQXFTJY7GZNSaG2Wa2W3N
+9ZQO6bYJt2krIfUFSWnJhZk5DUS9dv4r31nb8R0zvXvT40IL4sqFNdvwXIB+y8oZcxFSlf+HcuJ
qgeTbSItTK9jcmZJlmxY55Hoa61q8K5WwdYFajkj4knio7bo11jIV75AmNC9yNXg2vm0ytv6EZnd
TIYc2lemntBL0NuYD9IlwZc6fdvEcIqXKgp89/wYFKDeK0UVkdi6oB0t6UITgt+mM8/lMgm62Glz
uEjb8Tf+9hpX35qFlNEuyrMwyeg0BybxUZwCb8433VPixcZ0FEAFllx0VHtlnOT0rHfgk/haMTGt
DVqUUHyG3tS8uZZ0SRgexaiGtOt3CgNO70/DxzHNBh6EtcU8KPmuB5xZaFMnBLlZabavkZ2Ysl1A
/caUK+dbv+eyyyZuoyGgI/941frMp+e8um9ya9EP/7QpxnD0r3fD9OiESPUV7Z5rksgC/o+wQSXN
PiX35PRhiqevMoQkR8lbFsIhvD7BuFm7vm/AeP+qqzFk07nEO0Luyjc9dkizEwPgJkKLvIYOujJs
6HOgttf4FNwggft2SZFbN3lM2QSx30M9aWo9e1FhpIeU8dWXZbeBYLLRXAxQ4NtMYn2iYsxV9SPy
N6lbiPrFggq+YegnGCtWBfkWp/uku5jkwy3alSTJdPagFPJiWkVw4pJkwFjIIHrc28HoHRUBuq40
IO5NXt4ffGz1RVndxibjc64ByNdFAd4EOGwIFn1uzOSsUqZcjt2rOz3xaq/jRZ/974H/xvJ99sBG
bcGmVYn0VvZpprPL1N9y0bIemRTJ72iE73NbRCrTuedt32LUpU74N53TE1XwlCPKhGveP4sURPB8
JjCnoUI3WhXcTSAwaX7XmGe6fTzuR6wBLOK6G0J5IfZJDutfetbo+zmSFQUdj2Go6U3QepNzMST0
NEOFnyw8UCvnZMYnweJvuuR0BL19gY3ozAeaQtdLOYX4oJelimchtja85NSqvF+erznXqQ8eaSrI
jT8oz85w2vD/fuM+IVfsRJpkZM06a3wjKiEBJj8e75nlLSHFsl9eNuafaUJPR0gE3IB22LvNl/Ke
TkEaAsXBcakaDlVjyO3TKBsK2FNxLncPRL7/Fe04qzblQY4C2F6zQxKXyuOn8V4PW3cQvBJrsfHs
M8q7z3bZeLifgeNrc8BNxHuv7BUeOovYcqEmzWeLxILjqqSv5xa+EZ498lKQQDYFASyMy6kSsQiV
gAKG+ztwDgchcFJf+DLU0fZYaDQOqaI/sSCPr+ar0I27uxv1V7ZzPW/smjpwJrvdHY7574PImOIB
fQQWnrY4V6VYSkg5AUPhD1Ou0jVafxoCay8egV7K1vq33B5jpQtAySF0w8IXJacecX613e69g/mV
75zaygP/yBVg9uJ+qnYulndDMi7qJt9z/slYdXHZKudsRgQKcM9K0bQ1xWSq3wIfEgJOBGb8+TqZ
NKdTC5TZ2OzKeh2bApy9869EB3E9N5ZVe7kWhaXoMDuYErP7RE4nAdRGS0RXkHZBl5Pd1UepQtZL
2Pm6awqZQ3aiWXo6vWUrozaq5gQJCQ8zQNltxjhRGjQ1VpMt/wv1vS0uIQxPEaIMtfEIB60oXQTn
FRs8RyQw6HYkyCDKuuHTwMfzq2uKncLo96LLJgkwTY4MEx2IwBG1+iGbWJp3OC33+WwKwaLgko56
tkLOpNE7HkmMorvcaaQASYRaGQAZtdxE7oRRoOZjQQhFk12fuYcHNmgmcHgcj7S3uCKbEzm6SrOc
/NPJKs0+Ueg3SmmZvjOcKOQTPFMdbptJUAzcvM5GslkRcdVDBrTm+GYxCaGiC2z+3uMC79uyE2VI
iOGU2MPEFDINSyoIOzdXOXJmzt5Kqok6ee0088gIIQbi3AQIozzbs5s6k1KrSI6Lz6qcsxyOSoP1
hePYgLjyvRiRnvEy+jvMpG1DZIr7d+8DApgEPvXsIT5M4bbQnzLtxB4Te5uaF+eUZkiSdq+KUm8p
S3BrE3p0WOr7sR7Bu23vJaCEbKw1P8GhaRUkD9jum/Kwiojap0e4LeOhtQFIP5yzPG76cjBltR4y
t8GMtmOWPQihjReBCs2kmnhjyrmvUQA/CE/c/RCidnUILl2+xpfpL3heZGid6XWReZ2MDBWN390g
WjiPd1szFO3iT0lWymm82Iq9gxDfy1lvz9gM21heLo+ROhIQTrZJtstnqmoj+usR71yuNZzk4kQK
J4Enlmbw+yJ8YPyQNDdXrjA9wNGvUdPhguhckHvUhE08dcnolKGLVAglpcCWSo8tn7AtQ9t13RiG
QxZsL3obmEIjPMWMKU5gJoQKSa7E76LIzqA76zgnEk0CwXDIfagCHTe8NtNAM5vV7dq6+ydkO4K5
0fuhhWM84Z6hNgeVZw9mB56bGAiMMl9nHjmixZcsbu1TJ+Sp04PB92jfXois/IvzrJ54S7fnpGdZ
Rku8xhI+yGK5PM0PsDpt75VlvlXUFIj7cGQIROIUN92cFCaOazG8I/NXYU4GTCTbQ6uEsYgWx1dI
IYsFdI7UKBl2U+EGeRiDxjyZ9RxevtKQiZic4EPAaSRUMBSIN7Dwvx2yjA7bvYsyBnPvwdPmePcd
LnMnoPBl3E3kMcopmkb+PFTI+X5v2RBn89lLAgBqt+SnSVEEeTPCmsfz7yQ93vO74qA17GD8g4LL
xWr89JRUoMFkIpXsHmDmYvbxTY0uliaIw3afm5itgbu5rkiCBQfTSP9vzYNXi1FLMl0kTH1+xoDs
Mt/ON1LxJfZ0c5ZXbseb3lcy6VAauE6QWnmTbBQw1UPKBfETCQZHJNARAU5rAaiCIZ4PpuvMXPW1
WnBT4FD8NbcRso5EQPIx0GnYA52DcknJjv7GyP+F6EwggPoiA5YQoNFHZZSojsflTtYgCz8OXz4a
3UxR9Cx7pnLG914CaAsvwfsjjToXY898IjkCHuuXJLClW2ZQU7OjMcVh4ggIjJbDuARXCjbVM/iu
S7UVvBTUmJ6A6pmAUJuzOIWYbjaXjak9DrtImB6NmZONipnVuyzTWCpnuqzrixVZmzrfrc4f7UWy
CA9dYzA7lY8qQHFIBc2ynoXPFnurPsEJkF606lWqhwOU8Q4cPkRZMOoaZtCcF7w/4GdH84P/cwkd
3Rx3TQJXXPzsBczO8rwu2hOYSHkz3zTuO/BABu42Gah4fiH9TjqJFBwv1J9UKwF5po8mzwUz8Ile
yaNOFpFByOYI54zlSIMFQY8gR9rWRdhKrfqn0IjV0jCJJ6jjUgGtMUkiFHi/xWGoVBJQdvQneCKr
lQKCRXaYDMhWOenkZukJD2C4xoQr2dQnNbQdN0sA/7KDEUlutVxkzBOliWHwQ8DM+57g2Qa71Cl0
2nH2kXFQBOeFIoOnoINuWa34HKpMzl38karODxMhcVIdeCDbpZLEPoMP2nUx71QVFYHEFgCjiHZC
CBlecsvbuoUBmHbxEXwzAZSwHd6PE6C174HDn7k2w/aqB4VWmcu9AIKx+Rcb3mUeYu8t66XZb2Gj
953X4S27VfowgSOrhYPRe95vkUhhC55OdzS8TK7dfkgHBnFQ5+O5jD9OaH0yoIyEria4a/OYBDgL
wIOSBSej0RPhjdsA++j9Tb1i0l17YDWbiJm4PhHSUNhQZegFHfeV1R8zJ55vlnxMNJI8nEX8TNaT
R9D0gP4J4t+UAIil+MQcmaV+QMBV3O3k32dzzV3BL7C3Dwjzj+z3sxySnlI5Vkb1unj4JWpUyweQ
kND1JGcuc+dxOKC0drdEzV/6Wq8R2+DD/DOt5r92qZ9Sk4JVSNobGN80B5AaQXF4AV04AZ/JKuNU
GbXCliR3kBhSGi21dzS/yGksWcKxiEZlW60EdCDS0AM1/0AWNB5pbHXQFV8U37cD2cxkpdSS37Ng
NE736922mUvkNXkck9+09RiBzlmGmz80MvfXsCSrtPrHIjLuDRTx6f0xMt5/0BwptS4V+FUrSk+M
voT1yuIf1Qe96JtJ2/0cp3VLDhl2nRvTGMZYJJpGplk9FwkBHZgFGoWh6WUwKC7tPIxBAG/om2vN
pB9by1im3CM9jXK6Jg+/otbQZ5ZH/DzKIgNbgOZdRYb1o3aNFmblrHrLfAaaLwONLx+ETHA4odtu
89/xD6RxmoaH0Omz9iSVnKhUJqLunyo/JqiNRdKoCvg9eFq2vLm7BHC9erehYVfyHE8/1DGrQp9T
dzqbyPxR6JB4oh7ex3LdxK3M6XnBIW2oPQP9daG83i8tV2ud9+nKRuGRc9hhBWGDErKVNa7xUQ7d
C8dy6DqssN5yMkzYJEnqFYfl4FTl/0BekMoNeSzP4kiEIWduanVlb0mH8lqsN1MLYXVpgq0QvG91
zaV1uPTAz2GwafMRbaXPww6jDU1SgIwTtjbPji5aVlGkfqV3sM+25AqpnzSLZg7bykuiYLtRiliy
WJx+mx+DYbQbeN8ITSYpeC2rxnYWvHIfgRZO/pFSP5elX2uuBKvuYz25rWuqLmemNNrirNg8mzgo
L/QFRMH7jbq7Uyn8YieLJ9Np6XNV7CiR6r8VesrZYHlefTcY6FPhfBQe/NUUlTc8oyhSG3j5tPRt
z+9UyhWrZuW4xMbCcyN0fZ9fnH2x8EKU6U/lpNn6VvGI19Gf20b7cbLeEBPGivg7NcDd9hDUqV6j
1APZUIWigU52ytLYb/XkKpMKqXBhZJ5ooR/mV7SRIEK33dKGeZXADtxNIRzABosoJ6wu8CUxrcVS
4MDFtmmqmsDRxmr2YfJE8OEpHMc4fHsHK6wU0KJ4F0Z+6dY9JRj43NZz7myXfxO6NKLa+vgVVaSZ
7wtna96Z9HRxqEec3xs+WAOke8WrWuH9MxbhkVBFsQ3Csu5PokEcq+H6t1euzitcuzIz1IXfgnh9
iOZ1MDpkV6xOyu1Gy1xX9m8LuZlvjIgPo4zzdr1PiJh9IScTio6xNtEL7GsVXTYlM/bMTE2FJ5jg
IqJnm01vO6hxRMWRtVTj0EW8VkbNrleNVfSPOodV6g/bPAuATTKNwB5TYLkJbn/KLLWb7p7XhLmm
RM5GJ4kFZLA7NHupfOU1f6GNdkFaQFWKVQon9vopRyih0AuxjsubR2Qt9wb0Hveskter2DH8KuNO
joqVaKRXn3SXfuz5EjZ1AEiKdCMjjJ+REQ7DDq/IBV+d/YzJAVLpLJzviMbfZJGF6cm0Tv9bRiKH
mlqp/23hNMsa+CMEPOF6thM666rxnXobbJKw3UaDrjzbLylbMSheiSf0ued9ofL0ZfJFyVhwy14m
n8IBVT44uETrfRb9AAah3Be9QOwcAuPt6pScPy8avJbxnwzs9/SDjzIcAX91rQTW0EloWgbwP+YD
g9BS5cYXwfXYOi8LVMgC5aBN1SmSTfKm1q4b70GbcLyC+f4eIQk9aEHGRJ8i4xuLpNjrI9HEr0c+
f+cZnjnOzrwalN+2hdWRyR0Zpfz4IWaGdKwFeE0uQbiefLLdRC4c0mOVeef+UsHkDUDomAcPVKbm
0wj8vAEiaP8OiGRsRrF4tKrnuyaQYinQeFvhrI1zG7aAfEjw2OFAYwQR+qE8jR4zpmkLkLKztUCA
yQbpA0OBLD/4/oSErS6Afz0AQF1DYm59byPkg2Q9fJWEIDocgX7SNnp+nyTSQKeR+x/ts5pz2LpE
1yQIHsoLOIocC1WNXsWHt+/zrgtujhKt6WwBMiUVdG1kJkbUaY3IM2SbfYem++EpTZzJ7+fO+nla
u6FLCphmLZFHn/qwpei2TNElEdUF9rT++gv4OUfi6hJ2ZdVkzR+3a4nMK6AulB43iXVn7C9p1wlg
e4O6NyN+VdwuB740lJNDO/5XhT2kt8HqzZIx2zw3cZ7TXysYbALUxmcVUQg+2ZYZW5UGVGbP218i
tC3OKuSleh5DygwGVTkz9yE7stHHPGEozV6s8VekNnW8rsxg3bXnTkid14HqjC9X+cge5VcIcNDF
7GQyc/8qFtP7W774WMJ6mv/yPptLiYOLv98lKJO1we4LljPWIYtbQgH9X+CKcUlDJ9X/CVb4eXFp
aZ2h3FDGTQM2fhEe8ZV2Xk0nrYe6Gp2O8+lWFERo/Q2LeopKu81RXaD82cM/8gVR9JyVGbVboFdf
VAh2DJyyffGwkdfAt7oRHAgpddv9nyaSh/PrF/rme3imMrySUe1SM6GsmfqKK4d+SYi+8/COc64P
p5OTB/Z/Qnoixv1gojwqrEKEBrZYeTrhpyCFuF8YNgFZbK/qywvjkqDQNF8m/1ZTosFyMrDUXHUp
o/6uisnoPaapMRopyFVrIpiRFKzjzP3AbEbPsfprsEayPMISbReHYNs8af83hbrTb2rGxhFi0igl
d52u0jHHuuMne/X1E4euFEw8zvWxu7UimO40dqFRaqt3mhuyIJiUFV3wygfPxd8dGYd/Gc1xSLFO
i32e0XzPUdQy0EEif3E05nt1+sqlWHRGJUiG/+abzljFK4s3jJoIiDC1E8kR/Z/o9POcW6WPujMM
CBLaKc2RM2HYql/t9LyiYiwZjUwZ3N4+m68zvQ3RdiN5+OwNXQQBCpBiFU8G1+3xGWfS9MDah97g
5aaZhrg/PJcslwTNFAn9Tp/xFD1kEYJ2A1FYuKug/K8hCpjmYayBMyLWvJsefEOMXu9pdrTIq9fj
4IC0f9o04R3tVQ3Jnah6x1l23S6KWDxqVP/PHwJjZ7CrNneLf1lGiIuw66SEgBf1e4c7HMPeGvqY
ZGH/Y2y4rX++8J2gWfv5BdPJKaJ4oum7tu3aJCcbWUZTmbtc5QWp2EM21e2PmtlBDFAbZuaLfi/g
JatJNilcXElcKEeCsNGjFxFteJG4UH5yBdh/SUGr3j5+fC4yz8gMyIBy2fZuxVrDAxdgJrtVoYBY
6fBECOdz5u7kTPf4+d0j0eDDAgZPKBFrTUSnQldVQSo3M7qKO/WMYD1t7zyjk/dfod9UO+jS//Ia
Rq1uNP3Qer5iQKla0dmdqfuxRz55JumIYUwsVEqrGu1jAgI6RbC3mNcb1M84RxXDy0nZ2rwrUtzE
7OfO5Je7K+LUbp0svXN0R3G6YKhBPtCW4/TEKlqesjeuehoFdZDc+ANO18YYJss9uYMYwwaxN3Ae
D6I8GCfZqcsUJV+vSIyjUHFUD/C44FDz0ZXjHCCof5s7swHb9bCogNExUoBg1RzOVDOJXSih8DGz
NKcppfCA5WyvgtIWdxRnR/ZbYIp3YxhCjCgiCJlGUzEdBYf6eHoMGLs89MOjnqJWcwa36KFmhv/Q
g5eTTgUR9E0JPlQk/EyNAfKoJ0/hAwBeWiX44A9tJzImtklqq3iGUebFluargXSdmpBNEkcnusrk
fXFFOQhyfnT8idTVE3LFgkthEtSAjmBVFtGnGYK6Eyr8Fr4WdIrxVgjlMEVaQ/FDNE/sIOqK+QgK
VLlTizMXnXkY4v1BFmMLd3IlG961y0VbpbBr/RdVm/nf8NafO6gt2zvmarjknbKzZHg36JrAps5z
Z2C95euni3+l4Ye5Eg7FPqjNTTHrMrIJINoNqoNQouIs3p64hBlvCTpeVL+Y84czoFKGJov6WXkt
sy1fdsDTYrMvSONS6xds0vLuU/2O52yplmxuZL7OTNxzugIxQzFIPBDZCSW/6FIUPIFb6c+KIA0P
Rm+E8fPcShsc2z2Imf9SPKqiAqG5VA8kyZxOIte7HHHXthbnY6XBOZBBaI5IaE9obVcU9PWWiOhk
nu/dCiLUchqHdU8yhNfE7ksefX1O6bgHz+1wjm+g3pk9xhJsH58MiUojiSR53yCAo35htg0skqGp
a1w1WndZtIMdjP2Oi8O3kujnnzijg1K4SRitaCYoTnb1q7J8In5TYHZNwphrN3OlwT3KRzK3Xht8
xnaJBWyaX0pFsvSMK+1S6tH589V44XKdeBzcaKZG41VLstZcO6/B/EVAQJa3kKfm0tEHi3AUWDOO
QFtF2oCrImWB5f1XG8Sb09h0TkVv2rrCRG1tpEEjKW/dqdTvHVu78FMHyxMR9b0Xs7wU/nW6I9Wo
Q99/PVGz9JR9fCsAqGm5erqd88uw/7jUVmkPN0uY9MjpPCzSt8Iwq2dJQR5MuR3Am5btVnzbGWR3
EhxnOnhKUjasehqa0CL6MAgr1stxnp1OGPoH+rW8/0kXRBxn7aydiYY4qItZuKKlStJPvPqVs3Po
ewlPpM8gTQcXyW3KAz67ZR8IpIEG9SHsiba0OTR4UsFWsYleFohhTdRHQbOGUyYXgp0mc300aFJ9
KHQY9zMLvBm9fcLOLnI9f6f8BaGe9XglDNTTejt5HW8J81X4pCeV4FZ+jqMu1Evqpd5x2EdbMbfz
RpqpwuBhLY6sqt/22K4RybZCSH1YcXNEVrhfhNlVWFWM3jemaz1WFwoK3e6H0IvEO4T1Nu1hFTCU
aAK0wuWP3ITbo7H14XSlIvEtdP5cW+ayyzJjLi/AJZHaHUwfB1xWxB3mbo3o9aEle5+489xMZNmY
39dhKGEzDMDet8uriMfiOJ/Yq8c9yJagSW8ZInvzxy0MzcY9tsSUkB4E0rmBqkR6ieLejLKGCDAl
Yh8ijal20pN6FwqiuDLmwpAmECeC2gk5s9HcPxqspBQposXjPAjK4nNDesedjIfh/yy91UOPi7lL
yctsA40h7hrYQy0InGQtpSEfh4cpeGP6XV9lK70sCdJUQcTCEHowRUTsThqjXk6YVijClPjc0SAI
h/56rxaK6245AN5KS/PaeUzV1w+YLv42yfLv/TnW8mueta7o9WVbHjruJbBYlt8xNDMtL3xjdnFB
Rub2hUeqokKOPgO9AYTF9koJiCCDc7Voxud0cpYEYTFfdikCpCJYh+Ie+7B98PgJLlec55BTZkWU
spIJE2IKI6Gky8pVgG9vOR3oF+qpej3pMBG8Ly6OaBqYURloa3ZhK61WXRyWDgQsz981eYKdn3rn
Dvirn3fbP1m8jfiJO8cxJtWNHCx+NgpT6oZP485jOutaSLuF7FofWy40GSovZX+7sGUY3TbRHrsl
wiTIrnUBIJSaMnAxS6kKoLolm1NMabSyk4lyjv1ZlFx394YA9J21PhVu9o41q8Htx+bfPZpJ+FmU
BGYE2uK5RWQ+8Fy2kdhuBX9WSuaObkLQlrWUgda/jyO8pisOe+BDwTn10Rj4gT/Lrz2zUswmS6IN
eUlvW0wpWKt4JDrV1PvJDKRrfcKL4mcq3q1VKiTGEJgfOYTtZ/AiKRnlWVgqlEBcDnKEEhttOT3J
veyrlvqke3E5idM5r2a5ZoAj9eraDWiUGP0BHvBrFS8zKLdXVFVs+jS+YGtCSKjoN+ZK1hggxUrw
QZ5bQneFWh7PkaxM60G+x3wxc4zmI2IhFCHYM3Kun/jGySofPlJ1VJPyI8QFR5C4OnMssy+/c3IH
6XOMVxdDuqYilpBbS0OoZ8dWI9DYO1UKYbwcIPkTsAdxFVPeKbq7joUi4gcoDhtZYXi8tUIPpNNh
AdqzjmivxLYs0BO0v9Zf+swlfekdv7S2NKCHTJhIrpWh94BJH3gx/RWSmAQv2HniCFC+jkdZIESG
4gxkqVV01HTeYGb7vbWG59Lrd18UZ+iTss9TGKJ7vATZp8Z5Hd8mr0rPGiekIDJ4973aKEXNcGZk
LJtAUe5IFjYLU3by9Io3CSL47kU9Bu3OqD4DwKXoR1JGRBhkZsPrJ6zaoWfhTowbkHZ8RqmIkZC4
9q9wXRzz81H1VZJxRtpLeo12Pn7x/HFXUk8w9PFce7CBm5O1t3C1KZ1vOlGK+x+cSLpwJDATGlVX
c3KbsxG2Lin523ybzax3aPBEEtYBXNhEvz/DTgXCML6veOW3+HEJp54jqbN4csMnlmLa/ODOLBRd
5nSRhfapFoQryZQdOugFJ3XFsqJmdUC5tMWpY41I9I7y5VDDWbxWsESWUwb0DnXs1lmi+w6eEIc7
vgFh8cuj0jgNLWekMohnvktWW+L4pziwGydUzIL8kHdgyCVxSn4Ig+y98gQxZSU/WHtlZ1AT+LVc
fw4lDgrodIbzmtPY3IRa4YvFKn53QZbmebktLGdFLQoFZDLJd/AEo1uU8oQEPLHuOespCnfwlsXY
iVKHKvSYO7XzMlzfFJTSNn3GI3XtBKW7S6ZEe44Ltr4EBlOcU4JbJNmjgGT1yBlDw6GDpQUxGWv5
6qE5UpyGw0rf47S7SY4+nlK+0CbwU4GOszfp1RnYz2Yb5vmH10/j9jfUySRGA4S+DAqDYPusWlKU
NdLY0pNgTpwbCf4rDlDTAFz6ptl52bJce/vj+JWu5PDeL72G4WMdnevsC+G7qoELEWact2VvMkVT
A4z38JdldOEkLxO0mPbh9eiuCUDEZ6JEcQdviVrN/qJp/rx5+yjySJkmoJX7CPA01lfBtdbw51YS
51whYJeBQ190Jvy3ZsUbpgTabYS1Obw+QNIqa8dlvnICOd0aZlV/zQFRJ4OMtUKQuL/iuYLiWgqn
SwciAeFhABY4/Cba3fBBm+7LB0wT9g1BPx7NbzAW2STolRKS1rN/KB0CjkfUxY2oqcx/8dbB+wla
l91aw9bsNtDbF37md5kyIY6BBfXbxnbi7iqZL1VDhzh47D3GiRpr2IZzO1yoILs87D0EwetDu8K8
aGRCPM3AF8H4yEJpdAFyZyeF+nmsjcPbXkPDi7UtRk3uYnl30bk0kYJMSg3sw+BFx84twgpknGO5
V3rfofSWb/upEe1QQt6jFmQiwla11kOdx5TjogLwq6XhNsl4NAlxSrZnpCM8mmLMrBpD7kdj+dEA
bPjkD92CEbr/v8VTIRN8bMEE3ddY9v0UAwbLo4Pv8jCVUKxN90MVWbxeM14ax3vb2yiL7AfxA4L7
VCSKnKqUtEzKs4WaBZP5ilKrKoLXblcgC5FJabdvUmjVmPsACuwDiqvioaGb2p2a8zJx6KE++4bb
8Wp9Sa6LE5eeDwihAQz8nlc/k2b+M6Zu7wvWT7vBRAxdN8hVRK+JJZSYPPxEpgC99FVvA0ISGZN2
N2cYRBp56P9j6rmw6+NRrt2WEoLpxSF1CxY+pWY8a64Pe5Uucoyn23iQBsk4cAjj0qq+R5nBQUke
ZXWIxRadja+lED4n7+EAJabcEr6pgE8mb2kVFm2zJ2f4BGPnz59J9Z/qiOCjxL5g4k1bgXEJFIXv
rqALNiiKQs1H7fx0zEd00eO3hJ1Sayzrn1gTxSGLNOQMyGH40qEbtrlUEyhpotIpnojbXUXAziuF
lhDX6dFQsm8r08LpO4OSogC+2U7lWXaqUGSx/S6d25uRF53EEoUku4n+iprCC8mbDcESE7VQKmng
fQ9nVJP8Ucv6atfKRY3ZL/b4vOsLx9E9JPy8bm47gJVVs/muul//wnOkEhoEh2CD38L9Au6U45MI
UuBcJ/HALfePxzoDHS/pGVXQNBKGci5GlEHFdrNT0MZwTi5ZRUtABQ0yiLJnxymhQhuY0MxYTFHr
HTAS1Y0wxbS0RDM25UoDMbntxEO2ly3eynHlP/HbAIXzQLPkcx8VmZVmpJi/SSi0TV+KlaX3/Lro
+KrT8kqi/BHJy2vy3wRZD8v/ScWB9+Iw8lsbrs1hOz5cs12E90wncjhVLlPIBEe87bmaDGMEVRXa
knEPurwhkqzOQL9sCRGxBD3NoFmSotuk8RuoY/rOR0LpROl8hLfNECoJu8TNknYgiHJTLIB09hSj
EAbx4WlNRvljgExglpWKMHQLZv96jMeaa7pMzfUgGTtOk3ITD6ubojVJ9vIx3YG7WKYZfGM3y+6N
R5JkhHnBMt/gFZpMyKknfHVixDei7Hfw74j65+MfdBXoGZuCRC9Fu7iezOwNh/JRVtxnM17jiB6g
8+gmYoJejqD6QijnPmSfXSCz+XI/tImVdZy7PFeas2MtjMMu2QFxd479Y3exbkOBHgDsRvynxiwY
p2VKefWzST64ErpCYzS6/gjBC7uY6vUt7e6fqCJPehcOjlfid1dGCrvXrMJmze4PDmqFbfUh29ax
4xoEgiEGiXjhPQAkXgs5HHlVjGjxLzdp83EFEV5/owPeACxU5HACSuTBmcLH+1V2NYoROijVzKx0
lTxvdQVlobiddPXjOziBxjimA2GjrttrAF08QnHLB9giKQPh0t0/knDycnWHyTz9XKfchReWUZtH
E1UiDNRZx8AnHg2DdxftN796sdVacbx59SnMueqYzf3fh3coKx3QoKc00nW0z9rqhcxwU0iZzoQ1
xTMUw9wCM9s5t4SZsipA1hcSO0dkpaKCx7311GZESwi1cKX6f8xgDfTl0rhfbwNDctsBEqxkn/cQ
Ol5T4ImE7uTpxBpyUEZK35AriJiJvFHHxboT/7ogJ4AsEhvZBUgGytNBoUlOxyNq/ua1ptGKxQ2v
p9ylvsdbWfHEx8XAM6qUfX+7Snw96zJ7gF08WX4t4aQ6yU3E04FCExYwC9U49s7V1cmmiVJ7sx+c
C7cQHeCYLb41p2l416xQjcwFqaX0Jm0lFeOd09QxqPpuqQ00Opx4cnF1+rfQbSLQLmPgLZVY1TB+
aZ6mriPprRq8N4QMdvI0lfocLn2U9GnCv6Xyv7umcYaKIdA4j7YTa38p20ivMbNnHBXddt9iIEcP
umWAyaTPpiR/99F0Bk5WuJNlHLlBcjUDAtc0+/fYkWTVgOxQdgljHx4ZB0WiB4e+xThE7iYjGudw
reFb9IYsvrDMexFxAJ/EHTmC5khPxTmxqAgfPtyOOXp5LBtkCfS42A74GYQfvSgX0HOejXllIOvP
bH4Pn9cSGoCKbbYLYNSmV1MNcPY+6z4QaHdUZMPx+Dmn44DlT9mfWZI85mPbWMep2BFN/slzqqC0
fvQylNWxWuGVxw5ilsnO6Hz8LsYLLp1AepIcxpL82q+r/B1tHc+Kx1mF+J6wCDZengl8d3tLTL/R
3JkjVIJGZqOzQqp1hBa4mUQ9mPaJ49Z1KLFwktxP/fDAYKKB4vIW15Lloy+x7cPXd15vjZh5T+0h
bImPR988K0SnZ3AQFxL3GpHqOl5AkwRgdAk6N5QBNlJQBs8dhEfHxUMWHUB4czKk6aIcKJw21T6F
WebneHc14k9n/zJ5+iEJ5FaW9rsiqCEveDT4YZyolm24pfcEp474RfTgCkpAIXV+oPYh+Oe7U0n7
/eLHvouIG7qO6TrslVq4Ui7eZOmq0S0b7xDIJpfBqbIg35g3uw8zEZVrItJtfBB9+bNSzyn1Z7ED
jNY7we2WbV+ppmRWrjCY5OBMI4MnlcQGSjFUdkb1PRSsptAFq6ZXZ0RPAw31UZ3dN2vyHe2vLhw2
29Ql8zna4rjgt+DY8cr8pnZvWDcFHHMsktepX+j/KqXNlJQifKYxWt1iKXW+8no3NRJaWT36HqR+
TYV/KLfpU7p3/JtfLkKxbXWLtkbLqQimQTzchAjA4eAORRrrwaXeDyStbfFgBhyU8bBqY56cuW4H
r84o81LUq1m0S6fuCVwSBydby0zPHfvpvGKWRjREG6ncZ7dG6w/uWdikolVJoRihhrBMtWX1cg9d
Rho6INYqd9ogC+nI4LokC6kmCaNiMFHLTo5EjUGmNJMvONgLk1i8eSjTvPsgOh9tnQaQts2Fk+Tl
wBl+/1gy+GC2fGjTSnPr2GWZKB8kz3Oc73iE89QF67BFxlsDWzBpFU+2nEi69GgaJqhb45xtB5oi
dHVgM7BiWCZXFWymC13WW6h6pvQeUm7BNqsSeCZGLcwu5RYOWixC+n1qAte6LCifg7RphNTV4fuW
uuJJlADShLr4zOEaoUJNIo65RNtZXDTsQq36rZ+btw3IdcsQDMJZc+pIJ3QUKOdlbvuATcmHL7zW
KJupHlJEWUQUDWQoCwpDNuBHek2zA3gRsUCmCQNRzze3XhnH9d+SXJ83x8khVdGAYtDCPl4Ympjh
4uWlCP1Eq3BG1rRZg+PwCIxiNGxMTfl3RyNfJmHsi7BuqZUtrk/43kuUllob3NOdCLNBoLm9sLK8
TTinN3EEcZFlewOVtZ+EG0TBJ74RKPYHcvmvzqAZsoVwcgdHXPO3rcxhm//9FMkqwTuNOr24hAH7
6DdzJ8C97REpO8UgUbh7NO+DdH3YwXh5CI+1ADRaiocJqfzAhtVqNfWkW7I3Ytn8f+uFYXf8Ltid
ktqefMUZAoKCuhlEp0f2NWajo/vyLQ42wW9cPTA+34BOpXwAZ7Tjr5ZQAgnTh9jA8Gxqi4Ce0MBL
atmQLnY2JDM7kpgTQZTwkaKm/tgW27pLEhVlNxFsuWZpiMcT2c9QS2HotuvNysuT92Io6F4MrFWm
6CEM+zLCUZ1nXOvZCEgAhfsM7UCE99Hxy26D1HzYyMIXKtgu4irir0lOo8E/w2mGKDOPBwgs7I6t
iQL/5GWPRjiV/NjkHaEvYJM+P2pZFviZfS5qO/PHGw5cEUzW0rA3KsEN97OeewOB012Z0Ag/qaPr
nYb/FlWHrEr5VNMEiGvYBxqt2djioJhd1y9/R2L8LdLy0qYo75FENZfzmAeydmUvV395WWYEz0dv
3OsGqRF6kcg+tB4gPlZoHF8g0AP0TBEeuDwE1J9qp9dHCmT++6XR4XLAgP6y4Jtgu1ZPe8ATIP/Y
szPGBTakjRWyJqswxGiV/j7GPF4nm/7TUBE9E0biMEJOGzXs2epAq8ULv4eZPOq4YFSPRf9nNWg0
cDqQsFdRgE8hkT4KqFvoI/GBqk/TNGm3roT9TbTi1xjMBiZLV2IBx2PWthuioNi0pgDAb3XQ5y+z
TOyjOJPXyRfL/7gm3AzVvFEK2Fj2mJ6JPEgY8PHcMhiCYLWxBR9218y5VtDL6MkmGeqqgeVPfd9z
1V2EOQWRn3tOa8P5JjTCMY491P/b12GkpC5Lb3ru3RLpRD4XNc5AVkB6/r2xbfD3ngpUnSrbExvp
vy02OLrEpl0o252n3Ba35rrouFoXDjq2ZP6SwrncJ98TNj7ua8DWc1o5r1O6DGNvffCcH+FvN6Yk
GRB9miMm8QxDTUHffCj8bb9K4jqdB6T1e+R1kA838FOZfVLxHOXFWazwNLFEK1FjufmJ43tCpQ5t
LJkVoKGA7d84MedH7oehBPoG/L/6J3sx6Q0XQWLtIhDcLGXC7vHtxg/OBvaJTaKUok2MPwdJO3xS
2hvz6xX8fwW48FShV9z6FTOeM0N3nStaBjc5dvN+cfw7FVFP2Ikp9CVgfXenQysoIhdJgsNm9SOt
W5Ob8KnTsR4a8AheQp/kJ3eufRVSxbII/zqATspb4jslrdbBwjFPuR3QyV7lTg51S7KqOjN68AKc
wdj68ksmpkRbp+wm9xtlRE8lGGfuGYjL0xSE6N/R03cpaONyRm7kgMdMzkWxgc5WKKd2XcVguJFu
3YS39WUaioEe2A0ZBglp+s9O/wS+pR4CLy8UAM7p4jaNLoJIq0Dww03Mp6KvUDdXXhrP8iftP+eE
92NhfxXakx0976lz/TpXzHwGiYsc+3CFEAuhWy+D5Qoq+dVoMyBjVCltji/SWrWJH07n0QU5X9L8
8QH6U1t6j8rTUcb6KHzpKR71mI1RSE+ybYbGcwiIjySGaVVfVYSptIf54tn6+UvtKARJS3+7Z7HF
m/cxaTH1TjX57QbQ6kwYhivREOKw5E5R2cK3HY2Hj/iDrk8j9xigDe39mHnz6usuGN6lfk6i3TOo
FkLXIrvLkGS0W7hACULJEfa81b8PkPHz3aHXPnBAGBASiBXd+oUwf8ObPuJmhSi6rG1uxker5Zfp
lO7OxdedpyOhTEpKPmVUQo+rtByh0IW0hQO49t3tuxd7oz1lrgpQPYaEym4dYUw7thob09nJSU5a
V+kom4CzUqyBs+Qj1IPbIZFA5faXRsmx8wW514QJ3MMuLCkELIfibIaIF3Ks9CxhWPoXu9fmnch8
s2xc66y1sEU+mIN7shwcc/qOMm6djpeMd3tXdkt9OqsoOJnjrVJD9qAfhxMwmmVd6VO0nawB7Yus
zGu9XqqoWjbi2T0KfIKvImLgcuF0+6iD2sathRhq4dwKSk/xmxy03NM+00jMEppRexuvhX+pxw28
Vs0lq9rS2QEQb10JIMRtUUdafRS3knFD0NwbZTFpO704QqVDLlk9whigoJa833xAUj9pmM7tvGf5
vh+hrJ1OB451/ymf6fkAdYqalWZz0MuK+MhU9CDZqps9m2jFcd3tfGmfdhgSA8999vlTuPUAuiA5
h9S58Fa4ELAkaUtC4rRelpIBaDQNNenhRvmSFRO5nzxgKxoLlB2BKVcMSWxHzmAH61LMrVtcMqmi
je1DVypbG9xxxexHnpQ7OiMs2Ez80co8hc7UuAgORCOj6RCqTLBLWNjBqLawNShaFV3QsNw6+QMB
/mdklhByvECivxW61+z1gqu2BQNeTU2KUFoTVB5lu5boWRNqs81YBfSpR1QCBax6Gm+cLhxXP42y
IeEd9jMhiIMnbFACH7msOPriTfg88ox2wLbsB8WvUGxPKfDiJSCKDUbpqG8sgZPlRNEGhzOLIVeF
cov6K7AAoU1vwGFVgdoUVLkpVa1zGdmsCicBIO+J7exFViGCTJb2fjgD9MSHIj5dbBPc2CIPvfa+
m09NkUSD742VtUnzJ/8Lg+DL62YOua+Vk7xbi00lzVfiamj6KzWCBsMdUnUArQsSs+gnYzmnHmXx
IAyztnG7p1D4OE5lRHHQNmalv/YeTSM/yvWW11trOJHye3HpOOidRIToVKWTw0IdueVnFDG+lfXl
VdRWz/ToybDAPwj68Z3YKTgWLDWipffWWWC5qy8dkemGwmGzGT8zASPMSCIntPrgCD9eW03hMNxJ
V11S+S0vxIQYzwtONxmZKGbJI/jt3e+7NmmowkPXTvEb/m367HokFd7FbAdlA6nBIg0C+kDC4E4D
erjjobLbHkZFhHoLRrddzMGoqo9DxXdjknG7SjE5yoQlVeE28rHiZcb9UzkLcwpo5xk+G6IqweUf
VBTmVPSL2seMMsLfTz3mq3Jx93n06HBXo1PE8vbkY/BUH3Lv7vxA/1m8KvKliyehdSuHLv0SBlNf
fsrM0vv+BKqcv2b9zhPqWZcwvH/t0NgpS51vziLob4mdVjyz6MqW8ILvNn+yb5M2XlS+HDGqqPd7
LUNFragURczAh8Yp6qa/07KIdudgGeAoEj+jfnW8eYbQuiSd9xxAP9CMcxeJ1iNdLZ3Gy/VmURJ2
4vn02gaEWSvgE/rGWwsKE104rZ7d+nbab5EDaPIo1yB5kWqcaMxGSeE7uChwAqT7aJP5dcJOJGPH
2JFiUUq3gE3qHdEgjVXH3Kre2vqMEu7aNiPPhdHwWw+F/kqwumABtsp47h/u+rNOJfcccgm9pxqM
0gYpg+uqy7txdmUFpVfpqKxGwx9OphBhYlSFYFtKwKrfalBDfD3ViQRZYGbiN/P5wzdthwCcK10e
DhVztzbPemRqnu5CwUA3DD/FONQ7tieohav+BWgda+F2Wf7LpA3J8oXkofrGfNqvp8DtcCY+5u5q
hd/vbb1RTCltUt2ME2bAYGY+3NsvIGpPfqQRvrm6KypB5sAdc0LX74KK5ZYgpjJUIExRjyP0v7ZS
XXiISw4EGuLMNjnoYjZyWOi8xvemD7flup1Wky95UkiZh3bMxyBaIF+jNW/wOemg3/Ru7pr7Nqhj
Qh67vpfhFeyLLbkownFn71B31v/5oWbKxDPdcX2FLLTlBqjrhf1REv7Ey9CMMmzMxUuhWwu37Cca
qsFRRggSj/GEMwrWhqIt5Ji9CNLIm0egvL0Dpt3PlpOvAcTq24FXAPGpP2igQ25XUbPCh/ashLsY
iVrsMZAPKjdhGQJ7BgA1t59aAE6LTqzanFjmyQW5TuoyDQbzQBs/jU2xqMrnIby25gvVOTrJKtdO
luW2wnLc/Uch1At5o7y3bqg1aDpYjQH+0PV3583VSWel3dNGD6O0DaH1PwLs8y5P7p6s7Dohq5gh
fLbSr0Cbwb4Lxwc0wNYo0MGXtkZDBW9VFm5Q5Q2CWTXWGTCxOYTiUzmQXraDbD0iBNOkjfKnxUAL
ukPNvx/5QiQ1uqYiFiKmzyclSBWw3ZIcC25TwdWsnnS6ynkmd/BOhq7UbXbobPqIlJVQRkwbas4N
LbSXWDG+9yTgJzof5tsigxyzcuXMxWWaSkUHkSU0Pmvw/aYARTnxL4PZF3aFj/kDDy7cIZzebstb
S33Hkgnd/zfPMHZwwLoI/MF21W3BgXgnsyFf/nLNNHXyBy0C6qdLBDc1yHvgNV13zg0U+/MVtFdW
UT9pjDMsgTW+l3E64o13lx8tSvd99t2ZQpSRwFkbxc/CGx08xnJ5hd9on7drD+jIimjfX8zr4Jnk
eSo98kG8LiaFCUcbsMWHXvNySreRvSvJHwXuK/pewSoZ6nzBblPnlnntcPKqT9LWAcNGXNjeLQ/r
0XyeS2ex5n5Dou0ZVfQBhsc2+iyOFams2ySUcb6Fns9LHTM5q8G2ULWwxj2piUaskJPqhdU8lea7
5AAOwJREiehWWQpzjW89mn2YWGrpvSSN14qog++FJSQ2KBhs94ug68e3PWRdm+d+gcvQDZLZHq4d
mOt/4rBKBQW8zBGCE4RiuisLoXaePEeyqiYoH6tnTXHfjulf4l9tV/BeRdcfmk36LY99Ae+FPVz9
YDzLcXuu6a19m4Vfuu7PF8V5PNqfd5ly6Qk8kMsnuX5NFohPglcOTi18BTc7ntPdwwSnKWamXGho
jbWJV+fwnKouZAAV4qzE911u1ylZ5L2LtILcJhWV4UxRAgk3IJo64iNczmq6Zepi5Bel7dQgdma2
X/kmKHMZKgIYEB2GWUGhsSyfl7fUfw+yrEF32BF9ro1bvyAN3FNNHVh2O2WeCCN7uwQRsD48lY7i
JdELamFjAiq8UynkxrNQVH5P71EaoUYXXcAaFnRz++4c9iBf+uyZrKVyseGIC22HEh3bxtQhHSdg
3jN3DQ54s6IyxLSvfuIMIHbgdr7KrG95YhGZmv7IIesD7eyUwOXnIIp0swwKjvUcQRiAhAFkALgM
kw6sHQ+TOI87MTWkJ+5usmz5bla+5pjA2KEEVjMDcGy2ji1Dqg9XCJ+Cd+Con3nNksVEdZDzbby6
08VvFuEqT4A7GKbe8CcK67r07aAl0AyRCnE0Pg7bqxPz2ZLspIxtrdmLqmi2oFmrOp9gzev3w9NP
ZEAvtApbfxtMTTWTrkeatEPrxs7iYgzNOAsN3ejuivSjg9FboPhQPk7ZeFM7OFraWpgE2GLUvxwq
SBAaAzyJaNrsWkoip2lajwkB8luIVTek1+I5ltIfQIfzXaS5qrivRGVRSyqfyDu7O7u1zXaaBdy6
LyFqDMb9JyMLmSk3wVzgF0XvCSAArNjzxceTaLnM9ZakhLBd5ZKROop/iAlJTSzv1XVws01Sr2yL
P0RiUkOgb2eg9b9chOy5QSRBeyNMDHT6seZaN//KvN7fwwB3opVLGv1a3XzQWEwgMTrNqrEepayM
5mR/Wgr/nxvp+yAABqlYTv4dpnv95XvgXan2lsrqKGN6ZnmguCGMzvtXR7ue3LmnvXK3QXorQZ65
hgOWhQ2I/Jcx2lFqh4HJt3U/h7ipUyY7uxBk6Z3MbqrG9Wk6hf/ETQ/zXl9g4XXgF7uSDKXsln88
RhtV5gA/ViTZ6s3NF1wNq4lLswEs43p+41FEphCptJOJ7lqDu6swp5+ojykQNSKu4z/dfd+4o8Tp
5ps0dEDHdVVSeXrUH+i4YC2ydQw2du0meg3Myi2MzbQHKBIdVUcH2da6NDzAgK4QwGbQTFjHhxDW
kYko013mmTlxHFqIpFpbSl0I3RoazPeLe2cTYwV5KkKj6pnwAnsQtEsf/ZhHj2evigxCZddYZgA0
4tj5ppYp/NyDjwgZrbZhDUNKXIkVsh7kscEoRA2xzZ/DCReahJVbzUwyaT57EaSc501uPCmmpR7A
UA1FFwJaTUHOHN/UuXVUXOBaEY0ju2wQH8MbjtHnPUxV+pZQ19ZIzKOd7IFcO7kOT9sAobVHhzfh
OUAmR/OKpLNZzUHzzdYpURX81g/fFNkpYktaXv02VYZhBSarLLiARzdFFaA5BXRQL+tHCh/rCcco
awDbFbvGb5CCdjfi/YrlAr2YX6Sij/SD+yxArlKM0rw0nrf367hK9xnD+NQZm9yOcG1XuvCefush
eijCayu42/+vd5zT8ScFoGuS2dn1iBgwiDa+zV40M+N+MLBLBdJBoarZCeAfkAXZDJNybFquS0Gy
W9jYjpNNYfdyZJmgZRISELFuRrjm4bA7MjPs0yitLLap8VjfXj+DZn9vYRa2gMInrffsPyjmxuoH
oJ82YA0MDmPJ7DFc/xQm4RTEXqz5YLYcGJURt+EP1H1x+O+fF3l0L9pN11LghotoS00j8aw8gXDR
WJuRUF/YwutPUL1nXt+NlO+ah/uuOV0vQ9mde77SBwjvVjdfe/iIQnLwPMrADYTiP7s4Y16fBZpl
VY7JSB8gL2N3/qCdZtOuR44ORaIMJnEKVXtVN5VrWqqcjZBsXIgdKh0ZfqSqDwBIKkRhd5Vw/nsy
/wvsOmpOkpgdqOOsYnxekq7gNUOCOTzMmZ+EncLpTevcf2nqykZbaHVj/lfopOyz0aPXs7SlA/nt
cSoJuU4zGn83zZ5fSd3ff/dMiztvhC170hixRCiAVdziYswyEAO1l7qQ924hYY5900WUZKgtCdON
gR8OKMd9GYShotiAkeBTcxhh1iAOvAKgMJYJ5mhfwkjIkaLGmuWhPcz11yVhwjAU+yF0J1w4WnhN
NWtEoamhDmefXFCyMkBiaEiONddiMf+ZiNHElvpeR6vySnijaML32+nC4VPn+/5OcpTnMKfj37Zy
r/OHIskGBufMWm33IV9pz+cDD7AvhbfyrFpkhTGNO12jyz4RDI+VeFVelIFMb3OVyd7cyFiyb169
Dx2LCsb4j2BGE9QDMyxGDeLbbUczVnM8LRAqYh02xeFLuLEQWYNNTfYbtBevNrjxQzk8aKACWGYa
1QecdZkMHBEo3kubSOXY9gkuYdegVTNXwX3+zl7z8sqpQ1YmwsSha5zNZDyC53t2Ni3ScP39Tr0y
erABGtQEI/rSsGtk10TDypWFKwt+N8yBlCr7lp3kMXZLRiAI7hc2LomE3Yd3LDQYNO+EYdJWQycC
+MC5jIfF4b42in4SahmJEbXzuy78nhXU4sRBskImCht8PQjdTW2WvIqTL9uMOu25qoh9HCUy/YRp
JFgD6pFitc1Moh/Hj5J57Hizzsh9E2oeRYln7m6UUjVKjobDhaZzybFjIAl7J+ScLinORV6CZeHN
5oz4WpDECaXfTUX6EI2qu2aEuAAQDjqBj4AVMAGQtIaS42KOwxJQFW9NuHUucPFJVZu0nussYNk2
WLGUqwG21kD6h0nqg976Y4xdZC8Jtg7sXLQUIO1h3rY3OTcV5FSQeZOL/aM18USm4zOEm6MSbU0e
5tFlXveP0yYBgcTTl3erI3fLJK5u6JYSxHvZbUpcxX+ow3LeJ4r/dcyM0tkAM5ZWGZWoJoKRIKwg
+V+lq5TW9UV4auXXH8boo/AmApl/HuPa1Xhxh+4Sxa7YTnxTOKXuFRKgv/+5db3DuqmtfbryafYj
j6nt0xouG1y4Yb+Xps0YlL5VqxZtraJ2HlUz5IueLe+jGzdA5t+SeaJXmNeJlTbyq3rKplwUs2sa
jk8tXEaDBePpLmWnzv74ZFfugtAlqejxL0cpUNGfRuckNzLH03PVcu7gY76LZbTcdMUjf7scpGPs
d8jZMQBxlbUhi7LyT8HQfWe0PLaCEjzdKGsMJRNB0TeeuTBXK0H843baxUZzEArii7CH3fWjrMks
/YiNaX47Sod4VJDWe58VTluzG1UBet/G8JUjzgSrTgeBJ6HXqoYRmPLXkiYZMUR0GrzSfDjTbFrA
IfZtNJdGr4saDiEAYn8CDYE59w0AnxP3fevjqvD3j33E5guS2lBDBnxiBbst7gQtEzLKGXN+PfxQ
lZUSafCYweH6WcjGP8b+EAqSrYXGVi1bWUN1kYWGaTzDItbSKWYwCz4RUUAyfy3tGeflmHNhXtjn
eYVxk+WhFft/v97YZUhB+VEFf5ydD0oNF6+uUbCMH+nKtYL4pGubsxmR22aEk1EJ+pxSeYGeXhRK
PCs+9U3i3dja59UjLa1ke4jj2UyE6joYzJ7aiLC3gO1XgKcy3DPL69gKacIFruPEY5Pyi3ZuaqFj
PLjRZU2Xu+LsmaAAyjFS5MN69Jmq7G2rzAXQsBLZxVR8C6YEXhbAZEgdOE2sgP97se1HAw4Ri/bt
PvQfPrtdmaikdHeYjBzBfNglnrrJH0n64s3vAMVfkair0Qdnpay7jH0Dmo0IJ1cI3Z/fagSWZwk+
w8E6MrZMqHbIP6EUJ//oKVLu1gLeou6caN2ZpbIivJ3t00G+QhF23ONTS7BzKKAUVI1ja04aD6L2
WKxs+BmEO2Nh0SVhrksTnZtzUzHLK/FWFQ7OG7tvJmw+ydAZzfuBqtDb0L9bFu9JW2YBKkouvxmV
OEhZ8DY2vVLJRDZGBi2AC013lFZwofy3PfIxpjWJ/tbGTQ2vQaKwokpRyPNSPuGKA03KD+MF+Q5v
ZZkJPNgkLjNKVqyFs/8mkDNNbU1/YfMMhzar5Zsp5zk9l2kBVWXalpKV5gaQFBRZXnqwahdadww2
8VYvIPvgK0RL73RTiDbGyK6PSkv+chUwW2+2On5/lQpQxc3rn4nhGcsICjovqablOMq7WQ0PljQy
W7dlTT1o9c53DbHIhsCRRBGUgZ9WAkOgXl50c5i33J+5SBUpi1RdvD4PWmv2O6BsQAMr/NXU09Sk
xpaUcWtztgo2HUaogMIeTd//Wx1YZJEA2URqnZAdxaxOMh8c2/g2CGeLuvBaO+hJJ8RAZBi+WDSC
2EMfry63l0TZG5n8xFYjh/F37PqR81s7tNOyYXGveUMilfv22weTA/4CskrHiaghQT3ciPlt2hc5
KQKf9J/b9JXlNqi3hSVuNhk3c1d+0I0ffwI5MxUhqnIN1UqRjNC5AuFAy0rA6KTqImbFHHK9ZHs9
2SOFD0/sjgXOIEbz3+WEPiKszIpgWLwsEyGBNegSaPlFeUdnXb9B+5EsEajHDidNFJtPi+pg6mdg
z6qlftZhDlNCg1XFoRhUVrZP5jmYCQaHIBPgQWCnzk4ZdxUIS3talMDedzHbNk4LXOC94Vo7PF7N
96m2g+7vd8Lle6HmflUuF+4XlCx4bahYXWh/UfzNnIr4yItsepeCrLZfBc4lNXGkDv864PelA5lg
zlpT3PVGzD7AvMsvYNGG0Llaa2NDjQeR5SPxrzEbKJfniNW7jnDsoQolVbBLK+Fs7+wlHTf/rRMk
zsVhifPTokTVwMLQ25rMmOxGrPwPcb+xBo90W6bgYU6CB/2S4GsfVNc2tcdlkJL/9KHBrVRfkTzx
ybez12uFnR2odWfoi+s5l0W26qls8fkE2odlC+sQ79J8FOk+1GF1rs6JII6IKVKQGrcfvSYliylq
awcQM46gkcKP7lPNnOg5M/AeEJTGlwaihiPRDnJjgp0V1Dsg3yjCIZALmB09boL2BpWKUf/eLwbH
car3eBifE0p5IuFEP3urrX1vKs5hTw2jxyOPOd2mFnvr9+QA8Drcdifh/gHX0jgY/PwK7PDr3aIe
2k1ZD1tBHtMc7QKV/36GisQ1/FQVi4ohfKW/228I/Up+4QE75pseRc8A2jV0E+RzyVDGEXkMxhXx
r4DEcUsdVHVM/bhsx3W82CZnho+m6BrdUHKQ7fiE2xjRMK2eBZgGdqGNdg0TQo2DmHeen+ItzVjd
YLZukmcuQKvoAtNgdl5Z6ZrxkEQbqiWs5Zlq83mLA1NfuttT4rJS2JW5+iiTzhierwh5dPRo3lSB
9O2sybgpXvg3/w7TQnEJyMlbUw4/6iwg5dRLzsecUHsdP0oQqjQXKweIZjJtU4UXdmJVBBFBArMr
F0ywfK2r2MOvrfxitTaCYZ+lIor4jyZgZDKSTiYRY/o3Hv3v1aR0Yxv2NDCGBU3NzVkhGbNfv45b
vgjj+XXQWyoqD6ePzGqUppAKGf6uYl9AsVbFc8MI1nJwI5ILhGyho5+O4ECKlRH5Lw+5za3ktZGz
E6WIHLCqMrDvymEEk14xRlZdsGdjpfalwKI8XYYzM+tKYAr9jOyRlJdzqT63n0HjqHlKddP2gBeA
jF8uN5N8lZ+TqI8jmR+Y15xS1jH9s2KO83crjYk2aP/pwiHhzhuBPGfVM7APEFIWpvVXI5s1FBFG
6uw0TeSZwcfxCXIdoAtgdxdApsIEla25BIjfqc40eopqRFtAymWjmLqmRB87xAz8PJkIDPxhbmpR
RWE8zpQDXpVIMycAUNLThVF4pWZSYKWKoqWYJr94bQf900hiTUQW8AY/p/LZoqJAqpJn98B3K7h+
VB6Kw9NM6Di9+UteSDxI8ofogMZCOSpvCKGeLIzezePLhIofI04DSMmHKqbErzxGiMReHO+R3Pzc
jh5cXHSlwKBoAooPyEgLyihfKdR6UaqdMikjI4KCrPjWh7zWtHFNSHKk9Jy1BU9TGMmssosVMw5T
8mYtWMrfZWQaxHSId4o600tlF1kzsSQLHADi27DY6OopwxOV8HpUYSLrCpZyNak7Kr17vMWm/ZA3
6wcRYw9WRZArSA4U9aKk/AUbmJKIkPq5TC6SE7/L84jkhNk1TlRUdvpla8tIzs1PP/+1xTLtwzgv
PcPHgP/jhQhjv0f3sekIqNcd5+ljK7wt2+gkLOL9VvNflajwso8KEO+WJJ4nu6DD5EWVwAXR/GLx
zZ218yHpapZd+T1LWaTpuQnDQIPLypUEFUxZw4rbeWp/nOCX9apVaAcv4y4652f5gEVgIxObGf1q
zdSfSm+0CELQUKoCpN9Xmtjken6p0ijsV8BX2UPBKNmnxGgovMpx7vicaWKTRVw0VFk+indMwBX/
sAi0lctWWcke7OwWReT9ZpahPgPq1RfiiFObnoVT/IW2OBnUjt46EsiM/oYM/qBzfm4tOE/ahka4
7Zr9BFFuEPO7UZFMNXJ6SLXbAZ7s/oJ6PsG1YwIbJdadbxEmoUBu0+RKOpdHcAYDVdV6rMuTAQSt
Kyo/FNN1t8lOz3NUq8EDHGnD+3g7gRTJZo6FqskyCdzQOi8EfwNrjPQKwuybJ4EpzwA6PrlZCFyl
9oLCIwc+h2HJ/1pcaDThDD2PtJfl4zTtABDMfkq9eWtlastLuELsi0X9PVPVLPcpFOogM+9T4QOl
02BsQdeAJGd0XMu29zoBwUYKC9o7IAvSDZ+la1iwnvcR9OfqsQECNiy88nadhKh0X4ZcJW1Bnt4b
DnsPwuhd6OUi9kkxLyT2ePxxEVEE3fn6Hi8OdUXi/I/Yx2O/xG/l3rTbFntylF2BnvYf1i7aecwK
x5XC5MYCt/nfDD7qytpqiXR+LUXvXz4W5fP5zCeee5b1NeaYfK13yUZBkA8RikdGCz1LiYzNPzog
oGxnJAIdNT6g1g6b23z+Bxfg2AyfRc5tuKeDqFcm8Km8XMyW4GyCXPG7/ASbc4ho7XpNks7LnbjO
1CYNPIXE2kKCIFUh6lsl28sMobhgQLtinBrikjXjsuAgqQY+7hJngVIy2ioAJLXA+pQTX0rUnJIW
Ybqux103RkUhCgnjEIL/JLqPprkfekb7BPU2Yc8vzEUko1uzWiCjoqN+qDCw7TcEX/ZwYKOAr2Wr
6YrQfIrHPl+0jmMhNbz6JVvZNZio19hV6S792hjW/MWCRgsH0RaTayHRWkpYXp5fyc4Bsy4tktjn
V/fs43c/+Z/Z9afWH4xxmDlU0ZWvIc07JuuRsUizE2XnyjMUZmSSFwmDCzLqtWkvYWK1OHM2w7Zb
MBJW2i2K9CRI1WD7fPGEVIUt9FJWNVoWiZ8oRE91roIuYVrWvpujpLz+Sjod9xVjykkHh+e9b2cF
ux4loK/5WOeM5KgLuN2FQfo+AvOml/U7VBS11WxP/r9X/ZJ1wUcGWNXRw9CV7hL4HBRVGl23y0/1
W+sB9pbi5PmMTg21cMKHJdhpQllcenbi2gRIPfK1DMYUt/FZCvtR2xrDKmCbJZPyigB+u+qWNbqo
T6G/8KwtEuM1HouLCD1CnzS7Oa7Gwb03v5N1kZsazxRDxXf54jHU/C1CDQHYPExJtuKzeMpACrv2
VUN8ns68y0NuGTtoFCSHD7WHhEaRNeIH75TdFfLL6EANgixxa8uVBpqoV9m6+PNmk8IqeLwKO89i
mxSFA1dYFl4yC43E1+TK0y4i0+QYttOT1sIdo+jvBEe0y276g16hCnqo0ynB9CZuoM0RHM2iQt2v
KuP59QKXITYJW3H14JI3nuMloNO2qPEqG/dTPouM5lYxl8PE/kGvt6dHd13N7TyP5phly3hCNirJ
ExsXKzR5zYRFw1CE733jWmZ0NEajDFAQmKLs3hVjtDUbIYPCB36AzdL0KddtrbapkUkqepatQ5OU
/s5C1lQodkML0L/MwoOFLjdB7Oip40cvv9YpjDyfKhKoS3grCjovrq/lU5PGgxtc+8RvflEQKeYC
RYuDfeIiJfLf3q4/m3Jqadqm3Cjdt94+VK+D35ERiRWj6FLva2WaNMJ2hRLUoISmW+0C4s117Jp6
PZso2plCWkbUYYEZ+OfBX93/Fs49LoP58on2k6P5CjEN3vQ+5lBj5RJ/cW04vvF7vb+rBBCOPron
NAVaWhBnBho7IIb6OgSjGaYw7GKyME+OzSulzCz+uFaT0qAKQIuTNM/0Oww1gnHlP3qX2Wu0L4XP
xiptTUTdU1S5nBhUUP2S7e2qvFRvuwfeBS9dU0H9+Znfnso9ZoVlFVDYoYxr4GBaHIqMjTS+IzL8
aL/Sgu56C4yhSzjkxvyk6W2I1mpSyc7ZJSP8Nb6LcSX1cWaruosuQ2huEoFzNDCCH0wofvUNsUpp
Uczl2unJ3Y3t1dqIuI2M05K2OidPZsxP4Iee4YvdF2yEabuc9aGqbpYM2f13oDQJ3YWjoQGPQ3iX
dCuqPhpIRmPFVm7ONWiUA+rZoTBtpiwu73ujzThuHcAQGlsPgJ5jwR33iObL6s1BBMOytsHAJtib
W2hmKtwQwd7BAgPqlZtV3tp1+4XywR+R6t955WI0BHduIlufgsZHhCugpMKymUijm5lPxB91Y1AC
sjGxjHoQpcz5eB8FDLelLAcTmkerxWrARtcFXnlGvEo3UTgnXgAlp0xRoR5CNFYTDpk9Z16FDWuJ
XPh34X+HFBdSkzDO7o6n3Pr+AiQK/G1UFGLSYzDZwmKrJtZ9XcBzYvJUH+pwgT8echxjdFlr1Jyo
oVYL7xH6gtylvbpofSCiPktn3G94pe8yTiErjT01fYlQPdVkMRU6oxgk7GlfRlzPpiNhHNPCtCci
+82vpoWpZkwnSL7rYWaPlRvxwUmbKrSRtUJoOF2Mykl5DZ7w1pxnwvUflL5U+s7li8zQdtnHjPp2
AH6CgHyY8FPbpt/DV75CiC0SrRTli9B4sxi1jVLh/J9kIDcT21RYj5qFTd7XSEVRhUhO12p56G3G
dY/jS6DRMsSoDFJkeU6Y0F3EO/+WVTUSQ6CGjHY/nDBSXp/ijdL+2DAFUeraV6DxMKdJOIctH7kT
bS7fk6VwZbPIM+7zPE7Cyi71OLljiRx5R1aCMqehanaOdZHElYtdRbEUM5RIIziasfCP/s8VvNJG
wqDsszSmcpt90WT2hzVDyOaDDdCXHpeCeDYxs2THdaFdelgBQxy434mqV5WRy4zFFDT5GQBq7/vn
RzPyQtD/mYtxhjLq4adzjJ4VkPwJqjraTtJiDiZdmPB5al1V2WWyKWSTKXLefd/GQ1fC9TxPrdBv
LJVtqBHVM+QetTzGKYUwR7gdcSgZhqxBLqAetyztv4t+yBqtK/OT+l9OAj5lg+vdTtVs1rlK17wH
Jp1dCnguOSiw1LCPjmV0Q9jCBUDnev204ZAyS+XGUwlsTOEMvVDjLdYKYTt0/za2R+hObzCX3XZl
vfr5dWVxF2k4W3HMEieH2dNgk5uF7+o9Aeh71Ng82+PPS28Bq/G7a/RAKYw3i7h+fNixXTz4FCUD
rX6o8SdhHZE8nGzTzzmPQ7av28f0ZMmqfF2aT1+W16MtT0PIAW6ivnIUyg+aAU4f61cpOVSntHL+
8mp/gir8laDzbUoFllSN0ogMkFKPxW2dyrnjpdw+czfkp43fWVNUYaDhsw/uJHTiy1RYZZB+6IdW
B9slX6YVlBlkHZVBcIhsgPanTXC65iwL7gGXDghTJ3l2uu45Nz8Uq8DBRgxIyw3B9jS00N0fftEA
0+widrNHC5Qp6LN3mGPITqHMOCWdPXMxHVNp314c9CaBMTid4deFg6rkrz2mHhq3paQtphw0WNZu
xqvlTvl+3HMB+PlAKlxNaVFdxfkxwSmBFEQYyLcu1nqgsW+/xFbPE7I/UTsLWerIjN0ZyhMbVNYh
vzz9OsUQIvNWDAxzYb+cZFCAQ9IxVNrlyD9keaAUuUD4fjGQ8CWMEUegFjiT4V7McR5aUd3CPu+3
IPjYSD2we/tzRL5FgqZArPpx5aBKjGRwJa+36X1hrs1ZpMCXFezAlN3gCwKWZbIqrrybl5RX1ULS
lDu8qer+DPXGnQD1H89dTpyCzK9lBAk3iFqkexD8ojA7DlgkO6y+EBKQczfj9NcqXO3LxWWwSkWw
D3J1bDdK5qgVuJqt8YpjdmEZlQEjY+TmPqV7RdBLkeNpidOsNAia2ROmAKFI7iHwWf4NzY7C3YLr
Mupd7qnppaZKknza9DhQ0HiZxXs2vVNLr9JzASj1HptmpeosijrgTeTY5pnDetoi2bo8ZO1Ty7Ib
DVIqSRTfVopzawN/0rjaAlnxttVaiOiI/B5X8FtBkYNrO4e+lPOyvz9F/hbpz01JVbDFfZ3bb0G6
NUXEvXa65ILA1vBaWo0BQLMeYHpjRUbSZbYP3sL5IsckKTbWyhRW03r6hJURGSdl0RAMudagwsfe
Wa6mI+v6FReflLNc6GsPg0blEW3Iexh+7rF/AUcY8Fhormsrz36FbqkPkLXrI39uA62cmgcJ6MXY
c99FpV2s5/tAAtYgcMFPTl/mFik/fTk8rJUbOTDN82HPMw8ihi6sK1zuP6Cqo+nfVO39Ucknn5Qp
+EfTzcWCEgVuOYfzFfx4l6HzDHyn2VPJhO3dZdV1mvgcx95jShfltpq54uHOGQG5wZKszgKod11y
JwGAxPcmKhPsZR9RhWSi/XzzLjmzQbPHBRgu9iuvb5jmbQ8GcwQSQ3Zs/fHEdTXagpVH6IGp7Jjk
37BHmQh33+VRWNKwo++DDpe1a3DxsQukDY+H7pTf30T0mtPAbfFdONCpMDUcseWLWngLvf7Ir2f3
PAOpGYBvuzm2IVxVCdZbo0Ki6qZp4wK43DJSepAxdklm5WimThW37RwowfKIMwcPp/pQPRZrYrTc
DYd943gNCeTXv/zAMl4HxF4r+aXptfoYvB+G7JeS8tgvXXND+mE9WCPe8gEwGDUzoOWngqfJGYfH
yPyVaIxTGn8s3ycT3CKM76Uo2wNP838Vt3qChqDbR0uco0pqUimqynNWvUzx6u2mqqa9FqrOCFB+
PIHJG69mMOirSzGpL+Y+UqmEPqB6hpiAlA9FcPY1xbhBqm6gS8EZn3k4jCrkFPX5fAYmBAkQoW0R
Rvl0i64D0OStb4CeLOpRktpfcIJ5fRBaNr9LmacConPdzD1/XOJjiOb7571QDt6RNZWp63FkxtT4
L3jkpeNA//qDVkdzqfSAu0dejIzy9FdxLkxWeixZy5398zbh3/vkjVq5Cei4QfbtbMoKJvJaEbqc
PfW3B71Gso4KG1XNu/mBrQ51amdhm8ST2+H0PDtc2PJ7jy1pPmikAmMQ5rRSnLwZ9WD/3aaJ1A8o
iLgvkQZNAd7tL+VuSOy8XuiL+T8d2Hz3ePGi8WZMEINIOKVil2nNOyulc9/7DYa7H/Qbi3LSlmKB
AXVejNpcbO7UYRe+QyaJEfXgE0k1edWBQS8RR124dI5D/uP2JSnXEsYM8ARVLLuRfgrpIsj9EpeG
gnt4QG3Vm5Y73d08ItECqyb70bpjknqmQh/WeARchZcylnYbJhuA3/ey8kYRbAChurw9SLR0206K
bObaLOw04e+e2l2TWhQ4Ba+AggDFrY0pcgPOaTATbpVAjT6t7oRA1f967QbkiROhLu7zn+0XLMkE
IQxMSMxcyngZprJFLyi/Gr1omwY2feLK0bc1w9uLXLEWAnYjkeubPlWOG+excnvYdiDUqFJH1DzO
1O6z7Vx4mugu2HOLwsGVGSqo8blADaN6HYJAnIsJv6LMEz+NCqbRuYGAA6nlQj4XevnKVSoIFrJG
ue0JnLhAw0s0ISLZJr0q8K6o+kWuVEc5r8rOVaMvs+znDcaTouRTBu+ED6cPqNwgY8emUr6GyRTc
GEVGWXh1+JoBBYicQ2J47Aq4YR+fJV1anOxVZ65bHVGx4pGJa0W6C9fCsBPNPfaMqM7c4V2dKLmZ
5odzQrukyGr1WDFiX9yhI5lS5unUFJN23wGP2+20TNEq2pnoqGv+loM/HGKGzrGnkgPiP6d4cgcu
O+tDVxwOU8JuTCg0+5r6LAR5YO3ry6cqbyR1Ai7SZXIElrn+Ax5tCeVYBfcLOGVcvF9RVONrt/0m
XWDeLlMJD0DEFoWLNODXAi9/BsDeluG71cB2IzEm1kghBi+dGsahAksQWFHmBvZswm1GrvtScIDv
q3H8N74HTCgK5qS7Z0SH3mGG+pV6HHlSu79Uaz+lexozS4ZthAWwtm5hY//JvXk2A8Cdf22Sy+WT
KbCIrYC32dTz/Zn2H9S+jBdwc+5hOSNbAlMBFeWRn/r3d/QovnPP+VbLyx84iikrtLc/1DmG0iLo
N+NS6BjRsEzS0TnMMZah8Tykutr6aTmC118juci5G6E19M+q4NHudm2uT4b9ElpdyDogd36b9FuJ
1ZnjjiwQnZen8hDal7Tu5lgs1SnWW0PLWFiDEQjThIta8GvoNZjpL9GaYSOhwy/v1UhyRBTJZ7LW
6CZLY0B8JObPSUazlMyCbzcFFcMFkHIHpyKNzxgizr/HFvFLUfCme8tcXVXKS19+HjiWwyf0GIjt
vdanWl3aqvhIJ7Aqf7gHl3Wx6CKaSyUjMO0y8ObSfLPaWCZzSQOJYXtNCsdB8ueoJ5VAhJRpOype
gkjgnI2A4h1GhhEpoK8aNQLvhkjZLwe/7GId/rnloxZyMPLmZagmpKO/D081a+Pv9DEAsA+6qyoX
xDR/z6NV6sbXGO06mttf/rWXYzS2zILFwfAwqRmdnroCr07gX7oPeb7wwsoCOS3/zHp/N5QvHW96
hqBQWm1ECyYkMwZzrxBuCWnU18KB4Cn84IUoIPv2M5vPuRCvcilFGfR+gFJY84IwvEYkmO64M0rv
1p7nRxO8oJfkqbFgVL8jWvScpF4pDskj3DMixdNrjzhKpXNyOO5Pq4he68AJlZ//yzcP23Y1gkeD
By+e3cPCS3pHySH7ZqHxrC7/GK8Dfs3Cgd3nv3IdcA/AMC/d7lF1gwtEPsZDl77AWM73Np3+XJer
gdUA+3mu5dxCM4469j6trDPZdcwKvIdT1zLyxnkvXQp1YZDEZc/qMQ7YfapB+RyxgyU7mxMPgXAI
e5LdnVmtxq6IPBhNwUIHB9fpAWAsIG0wocG3NlbF1Kw3NpG1uMqbFGvuTHuIKuL4PlYXtu1rqGMo
42dXfFnlT2dwZK+ZumN7j+OouAfEvSvtW/pX9STxieKSee3o5LWCaAJPZQHNtU7+5TQuKefKujUP
0l7PYW0R0HqTDWQ3RsBoxGV7Bi7up0XBoHV91sn6lXVs8rOzz0RtaQnnIocB3nXepSwte/HwtP5J
mBRJtoM+6sTOsewORVOt+mIMF/jm5mZOQ36ObbGI5KJURhTyW3QbJzQ0zXUUN5Os9VBfmQpBD7FE
A4qtPoBg+kqcDIVwKTxNzb6kyKqZSHhLy85klnJL3/4bh2ri1r5IETjkIeq+bA5lbrSHiERXh69I
muTGa7ISQ19xvHNqfI3GgCHep7KWayFMozNKh6QFNWY2jAMkLn8jUN/T3z20qqXHS/q9fSGuzM1t
1b8IxaFWiDNlb8BQmfotECFUgEJ+ag38z4vmuFt/jfjnx+fHTNzSD22xMCu3qR2CrYMmWRbiTtVR
iPwvNRWlUNEDzmPAhy3kPGmVl99p3UUyod0HOYVRmFxXHX3lr+WgTPg4srINtH3EvGmfcWUDuHsf
6++TKNsdKCrJSqbeUALy/ceObzc87/ybu5umZV0YLyP59cKyWFFmoflQ00oSdibIrmhtSxSNGnW2
a++9ePa3iSu+0td6A4FBA9+747DvRhGo/fTaUZ5RIdHDEbMTPusLRFIkWJmmtGNIoOjkJsP9M/aD
WQKSLYpoyXipsOcQrdlzxhMXWBR7pFsjSXydGWK0OVwwqynPJ1lbl3WmSwLL5zwyCDQ/NJOU61hT
DprnhgaBliFIfapKRJuug9JEEfYR656onlFSouRNRKlQYZGKo+udBF1EYhfovswN0qRuQKxXw4/L
SB+riULS9JwV0xXoo4aMa91szsC8Luf4HwJxN5WMAEGIQjqeS4+vAtCD8vw18DHZui0oTHhfExo9
v6RM1d70GWz76Sb3tUYbCkoCAQKI/VRuZEjuW+I+0O++X+wdpusytWS8wcUUt8VqcpBHfPZmuA07
WFl8j3KYKbFS4ovYMVQ9HMkMLBPF6ZxRaxkQ4NcyHvGL8x4eMuXwE+agEihBhyCa5w5CP/ua/yw6
+g2B4ED8MM7OZfinJm5YkAIrodGhtyKzt0YYSgQEzb6O/d01EufShK99BHniNMTeXd+qJSbuPrU5
ef0jH8hvYQCU9K5S0ToMVJ7a0zCtEYRej5arL7PrL134XR4/L9naguAoERsMtKuGhZfCsxd2Leio
cojNZJjCfdHvrJha2sEnweU1W+0P/jUrs9didq8sExgD1hQKuUWRQIbtv3I1WHbin29C2c7/bP2s
0vY2xfD6XCZE8hotQa8v8eVc4v2hZ5313qnuBWM3geoB0I5kKsMkCQ4nBiT9CyCVuZv2FhPVDiIF
Pi42y+Vn4EupYM2wrxB9q/5sE35xsNjjVV90CT7L5wn3vqsze3yNHmkco0/uOvZu3yeSNP5sYYSk
Tg8OxpACM3pPTcIK/UvTWHFapTXulZ1rmqk7nctv//SqbHOw0XvYLRrV8xFktOJMYxBpKhusLiXJ
La1kL5cHLgsTjNSe8H8TuEDD78ZIxvZXC9cDryXGYyQyiFaWLj8/3bQjWJy/YmG1opkesVrsWOD+
Cx1R4zgS8X7ogCgpYlApDQnymC/WgULAdPIlbdzhI6AeFgLaZTk2T3kOqoIFhC26KAjwNULG6rkI
gDkoTotuyJhlgoKHeNZO0QHdIuuFEKMiM5YLnPwqXbM0pghNLaPI0wdJS+KvE3lsSLmBWg6GKLr8
wU6JpprIGgwFgpxDt8wt4nR3KHvY5B9dVtIR6uc3bEYUQ05ZbOehrGvBYrcG/Lg1D7vqQjgqi717
jnxYmgQZYwWt2yHLBqEOzy4hzNSvg5SeiFp6Rj1C+N9GzbvsvW+h3OE0DQ86Ov/5tVPemu28FNNl
uGvSpap1+xhaKjK6yeXvmtezEe7Ceg4sx6f/b0NKXq84ntxJhQ9Af89sJhxexK7kScqeQm2dg50J
YuoyvOOU41mjuGkQ74DOakM72pjy76yAMJvgdZbkKxdcVHyTYvSgHNJlL5npD56TTr1OK/INYTuQ
+NzwElLj37fcUH/InqhY8CcE/g+6tOkdmfIddFe6Ao9GMD/HgPHV+P0b60Ob853TupBPJ/5nx2FS
Zv78/zi23D5KTaIHyODCRMcBOJynb4/kUxQV6h0QF/DOw3LsApprk/E85k2yhMBDChhTPM8mCVOs
+xDVsFoo8H9ehfjTLCIDZ35tScC4HIFBb+Fj1PLHAz8mzNlf+MbJHfszkYf7b8P5CPEomq89cFhh
VDj9Ool730td7bOjsy/A8N4eOqa9pGXnxstkGT/yFJcxWAiuvmlMU9dcOTiQWUvlgIR1nydyfm65
14pCclG3UtjKT2s+n7zoqi6eW6HAxbnnE+r38hFbSgPcFtAEtCLc6J5mOVLLRUF9/ottRQ9ZydrL
NqUJvgkDGFL0tpwUqmgbrRI6lGN5MwjjML2yAc9OEQga2W85XsDfPHvSenkANkPQrJKYEpptIuMi
JRKF8x2kvfSiQdVEUy6tl164BrdL5RSJixk9GU869vcxc0gPdCGSHQ25giEty2iA3nKpTuggmiTx
Li/kcUYRvty3YFZTEmGRRXRUs0xV1TI462V6x8GCMopvfwxI7/uC5vdQKptxcRZH88a60/ugr7at
KVM25EEsl2nCl+WzeOR22SvnL8Y4ukkHK7xeR4oysdGfWlhuJF8j9M1flpcqCGa98s8IuPZWGT2S
AvDOa+/bP0k2Qw+/+07LQyNug3tT3PkdUJlI2iLyCfOB1FD+LZZcYFa1QJQQdbUQf/rjWoWGTI8v
/PVxJO7DSaZ9Sq3fJhaMM8Rq9E5yRxuvdr/6Qnd8h1VLMldfcW0KdPzsXfNhC/NRg0/XnQOceOp9
9fCn7apdiEVcFIv3jlfSBQUGB1oBi63q1hxN5vA4nq5IMojBJggdUJqYQ3qKt65CJQNYrruWdk59
FD0K6HjZGS0/ygdXjRdVMENp1ExTishKVi5Ba/JUIo7aXFTV4S7NUwHTqKmFwX+m1wuLPyN3vTHQ
dZQY97de9CM4tISa+zJeCJ0q7K7qs4UYO6Mf9iTPsN5yzkbti5TsKFCFmrZXyAIMAtUXTLAJril/
ym79XcRxzYuGSYnEUBunaDpId4aUY9MD4DfiyQzwTPXoxTWqqtSq7fgMzD4G22zwZqElC6yOGRtd
YFF2FCqtKHyvjPd+coX4XgKL2a3Fb8OMM7L0Wu6ICwj/1vdORffh2bO5SuiiNg4ApSiWSJCgLqYl
Bm+Q+fGL+TfMuFfPxJzDdVrGzhWusvRwcSvby2AK753f5fE1FQ0/YkPVfU9HQmpo5ogrZGVJKnce
opqJrhtMXCd61nW4RvxcXNCj/83J8rqgavdUGT61OQNM4BXcS4UFHkouRjsGqk4ZDfn5dzroakPn
58hJmeys6FjWAAHg+m8QCtj26jOTgiAUP6KKU24nZ7iJ8h4IHNQkjdWnRGZ+p38knMEygzotGjcs
KL/u0WnEtq40QQZUtf3jjyBNMgpZmjHdyEr3s1M7Iwo7K2d8SYdoi9pyyDhZsVhikb1dj6zC8GMW
ngX4r87sAEk+ZpEhbMSWYyd+kZgNCBmKQ+WK/UjAi242VjbyikpG9jdY51AFk5WideqhZk1nSszx
V/+qyc60FOUrpP/RiyskY2MMDtLrkRLTHXhHfI2U7EA7PanUcLOLAI85yA6VsReMdVdkAgigFgix
EeanCR/VeAf9qO3adzzGlQbcbDWnhT+Tn/Xfq3gq9KTsZwKJAZ4E6iAYNG5/4ABuJxWZh4JTlvFS
P1n32JWYicFOjCUG1u4DelfKcCtxuwYpfv/6QyOFSoJwiMdLWpL5J61dfTPl+M1USMo/xPNjv6vZ
urj/yHyQ7MjFtBvHaJiBHZvL2tQmBBiJzTxuBUrpTR8BCYwbRwYW2E8RvLXT2rLTbZsvbwNcmaSU
51EyvODD7DzMGFgU4NwQUnM7iF9wLjBU1AXkXE+zWR3WJi3mTwrobSOujijwGjdRIMFZk2v1BNwj
6Y6wSS3VFt2xhUTzFsv7+mifUL+LsEITEXDtoJ6QGAM5WN6AYPqy9ORK/eoy2S6wxYTr5x18rmuT
kECCJJl0MfUFYBoB27fF4HgaUuyLvZKEpYyZJ1BPXlENKo7AO+E5Sh0Te45FW9nQ3luNBDJCsbWU
Za2hDDK/UX2qZZXXdnnvySC1a0eeEZuema8+mjj4jxNWtzl98RSH0A4ryBr9bprZkDb2vA/OvWUr
rkXL5zVHFniqukd517zvBy0d7uTbuMKFClmzP2W7nXS1TmikxjE4viMc2sHqCeJhUP719GtxFjsu
mk8Xef9XONTOjYIhdacRCJIFV2u5AOoXuz6KSduOmvYUJtNVd3TVNyIZtJZmvLa4tYdEuxmu9eYd
aDeim8WKW3hmm2nIePs+40vm0ma/eQ4w62u+dQXoJ9Mr13AEDIJl7MB6XZUOFG9RsQVWgf31QbA8
Gqo1CIx+2X3EpSzK9N7qFxrW7bMKPEfH6/LiTcu2+es08NiXQ1dz8B4GZucQhsmPD7J6IOttliVe
SrPiyTFpuV911v+HxN/yP8suGxpT5NYRgLlx3u5AwKQLM0bDLPv4GSnR7TnrV8HvzfX3ZfBoV9Wr
pfHYIB/BFsUURgLWMUdMNR5MY0KwCQ/yH7li0gZ13wYFbEIy54qPwK4qwzgoXaCM4bvr1ko7sWcV
pGytpsElT0J1dpTaxsPI1EjStts5olLBwZTR0MQwTS7MxP5PYNJNZcFQMvSFrHU2v6o2f4KIAG/J
ghfqLadQokc/pomY/v22uuo+xsNLJjsAby3KgsIf/XMOHla4kS4dtsZUyXhqiVRgim73FzzEmqqz
RWPHLJw0VHxh6zBCH4BW/VvL1dR/YIMhCO39ZT7Pht8AQXxrOSpCaQUs7tZfALT+H8j84qN8uVuY
lz/UsP3CruQ0taqiJD/a+cvcU87PsCqN2CVAg58ho911y+UZDJG1+eSnq1ZKJ8ZE9PXKQybjlea9
m4qyprMtmLho4jHPW1FhsGol2dSA7phOwIjLLpPNOPDwHH58Qgp6HipLdUqoRgOjqG2wS/Y7tYiN
/wIDq33uSTpcQcBu3k1tvZ6BHLdhw3PJqjLruxCLwKSOSyWP7bWlXeL16wG6VZhp0f7dLFmgY5Yy
5RypEO/lK9SB5fIyaSiI3Idma29wW1B9fLN6U3l03g827HvrpxjfqNFRvhgpGKQVfsESu2666PEk
ePQSRIn5kn+d7h6Jzst/qMrpBCrXp0J8gbTV4hsjJny2ykuMGTvYl7qCh5SratBFawvYYSt24iot
DgmJCPDD6QIWaUzPoElW0cRsjf8f1dZwjMGTuwrZAgzsqrCK1uVMPJq12NM10mDlzlHmyCEOvOum
gjwGg8NebMJk0PoWdnRfZLcMX4w9CjbfZbc05DpTHjqc5EsCN0StTzpO5QkGR8F3G4OEnYvcBEGb
NeSgysjt0VttXp9VDuZYzL7LOwOYVSsUc1XlgSo8h/J7jAWV+wn7d4vqoxhQyjcNMDVOo0579kuH
2U1PazSh7QST403FK4YLe3zqyMYAE4Bei0OMu7MugAgvfkPtZkl1arJwmoQAHGezJfD/5a9XzMGU
FHWyzKH1korddNi1Qx1ieCFK2jdWPAvsNjW8HZSX4s/amqzj2TX5GogFCDyG5hNVShOdHShyvqQw
Jp9nqPYPiI76pIHCLAjV0nhfTQuHTZP2T3syhI3gi8aK9V/SQBfr5qrFt4CpdGFv9x6tiTvBA9TB
mju+78Zpbw9PeP5qCpYFBfBddhW0H3qMMX5OaNQ0N+buqw9uSr7c5jwjkLP19zCLjLeeckAKtFFV
d4SO+CZdiIWP/VX2hJ/UNsQ2T3WGwwe6Qo/e6r5oEVOkh/QqL2SA88IExJ584j/uQjhamYJFANiq
e76gf6KxFDLQ1w76j+fMcR2rj5SjrWDbsYPJ6mitMYxu7UN0AC+EH1bCPPC+//tOD+dWVT4SxotD
GEDm/v3P2AjvMIsn/d81rAU0ZaDc25ztHkTzU3dgOp093JUpBVOq/ZlGxkc1MJPCgDT5xFWcjXQD
3oBG/Fud9uYkwTI+h5BRhpfGJae4NqIcUjyCeb6ac+9LEbB2LE5ULiTupsCzHKc0yDs8GeN/sOao
0/LAbMXLWb1HrD2yTuwKoVEZ5BcRNqxK3oIHhijBfTv1596GpDMgtCysysOxbHrtvDpmUOaKKlvs
1xsBLn3mjIH4WZO0a5kffRnXXXmBFmzkbJ5zI+btRVTazS2FuiBXXxI+yeMap1XF2NGxDLEPHOam
gDbAm3LHrOGb8nhzwpF2b4k8C+3v5TI3kYfP8ndmvbLwmMf2kebvKNKJXjBp4V38wMnySBRLN3bo
Nph6k/4CMxkNjs1aOx8nYXLX97tcs8T5eXQRL0SEA5uiwfsdAYxOaoNpwnbsGj/CcjKBNxZo1Dv+
pvCUNuGTLp5SV5XQFZDxEFtEfO+0qdNKvYBlByxZGNVED5jSMs0oZMAthy3+X5wvqZ3VP/MVs/9i
x8a3eGuQyxyDtll3hwWd4p4ysVayXeT9ZdEnyRZjk5CQTLXK8V1VcNmi0+RY3S9LbsWijVKFv/uc
xcXNa8vCJajBFDQG3Nt/ACT9cNB3n/vVvJuw44AlfewF68VrakM/ymTg5zgXTNFHco5jNKbAh7Q5
aj6zVVc+fDpY8cp6NigSR+c06nyJNVqfBPrjoPH7dtBoD3CUP36m3J5GtpUCd5Qj3v84qgEEw1tk
+/rRMk2P6XbtR6ZmNlOapNUI552qYetG+D9Idh3Udnvn4iqOVb3cMrXXVzXRn9ynF87DBO8kXr97
jhV3OUt7gaRKbOO6HjwWRIJVEUJUqU9/fGP9Ask9AXXed0ky2J59/4ee/uy5vRN07kcr1jlp3BmH
7kiqI+4qZgfX6dlWqN+4nCyUgZRmxTmdPUw1GMDIl/1HY0JLQRmDvOVHkPbe4pASmXwmnVz0BoTe
HlVm79Upf5qFda+jna73ZjbPvcDMmRXcIZuUA3U6ikUZuegejgI29OIvc7T8He1GmV9dqx4xijx2
d1ntXIwZkJxGctcGET/g692khW1a9M31mHXv6BEt0jFF5C3oJNvzlxDqLt0VyREwIHUTlTjxmBMW
6iWOL9rlvsx0KDyzjujmOI4L5RuNCHvwpaXdYaLm+vVuegiLMqflPkFOGg93yBJMZzW0lGLkXlJM
nkVtVZ4mbMYXAFPjSHzcD/xRLfDR/OuhcO1+euogGQz/PNRiwsS3v/79IQWJ912bwMPPhxEfXRPU
lQFYXbH75YHb/nxA8ZiHCGwKGyB4ySuThDTkjfgQrRqGciAcQZdUm4DcUkAaRR7xLQ7Wr/H4HskW
33bKgyaR8eVJzZ2BgrzCPGA4rttHSZSt8XjFhKky4MTVMYWh5TjQiopnRQq7Kf9VuuB4/lLu5dQk
YTfhw6wbXgGvvTM/upomiuxjS3PGTJBpzOi3VfLPA4WqJVL1dXZiQrXBdU5FE89G2gK7punWe+aD
azzfTqA6BX4ikFkI89i9GLgmar3M+0k1FWP1Sk6/IbT9Oq4rYLzDBSP/AXTJjqifIIZo9iQ0oSgZ
EOb5sp1REDGlbt7a0Z9IFhyB2W+2WmsYA5CQ2CUFTjdCeUV2w4ilHQx45NKbiiSnE3h19ZFqB2UF
b9IiwbB15TKAzzhBpIrj2LzhxqlXwRMeGPYx6phvYJUwxLO3sMWO0uSMGG5eadw6WbsmqStFSRQ5
U9mnIcm4x+M+yRSZOwv1/VQ4FQI2sq2N0/CSXebb7fc8i6JNDzyD7dgZre2/5vZeDhzwe/JEEsaL
wkUTWGRLGqnSmuCyKty+RvXUCqrPnalUX5SOJ6r258fF0DLvi7aPVyCnfM9/5TIaM2b26lSyC9Cn
VgbQURIkRUbZ5MzsWqKFT+s5m35AbrvNSLpQI4WDVpJCdlt4JyzWhoMryZMkB1Q8344FltHsBe35
cZe5f/KACybQlrxdpkR6lW21jCR7IiUJTMYGucWTD5MDFDM4exfVRtQCrHInGN4troQqbwh1sdaF
YbYP6NTNXK3SVbvhAPb56kwUik5Twcim7GyLcsUbJ5seIr7a4lrZZQTecBr9A6MMSwaGo+j9758Q
T9XQma9CsdhqwMu298DorbSn3s5uRdGR9tJBuZaL8GRf+IaFJZCXTccMN6bUTkYF3IWJOtYvkNEc
5g7+H1BVwitRRiD6ABpK7xmui83ekUS4mlrWwMLqvpB/2f69MU4iIS49uCdvaEtGj+IY+op2FjF7
CDkri0Yi58lkTrpMPFP9F4P4iHFiSW2981uhb5SkgqMhwrb7jG4FeT/C+58XETqBmv/apm0aQjhE
jvmpdopHbazDsRd4+290E8flb/1k0j7rAXmxbmSRDaDrM+CbLq+eCUgw5Ljn6OfjoxgdG9DyNvnX
QykEmfJS1hZUMbqOQmPY/94KZsQ7EJEUR3D9kozvQP5P2tv6yE+Mwo+B+ZhEXqWq1v45+5RVDK4d
sCf1O+U1q+xyu3a5S9wtSNJbiuNZfmgQYI6qf8JnrRgciobywCM5zxD9rchAl7ki4wbvDhW8zExC
AYhX+ugfA2d0oGjXDMK1amn5ZaHpm+AiSzkAIzjcQyHrveCLS46q/HY3ABHVmEq/bdAZI9/PDkxY
T10srYO+ZNnldzVEsssn0xvQOPK4ZdVsRXbk7nLExgwgoGaxXedgRceuLJt7/zp2HSL48m1Zvcp/
N2Tbot2rQhu84FiWaClYTmDBPqygKaxB9U3LzZH+arYqwoI8+3OuWJYa8tHm2+hQlm96Plj5+PNZ
P0NyfhSKf+XkYRsHmYPHIffdFwDe/+TXiElEVU4lJjV+QYB9hNzTBZIvNnzI4m3B28RATxbzeT1+
YWH2fiab8m8Z0jxmJbdGbhtdNsnEiyD39cm2lTAn0DLsPtwaADhClRZqe+dqumgmtGgyrupdUQ4/
6e4U7B1nYjlINs8Gb+pwe8PuP+tuSWbZRRpzaHGc28YUSwwxp5XSMrQtA/pY9DQ9ZQY/tc+zxoA8
1fvgaBUeCK+iEYlXKfB5Pjnz0qLhi6ecvE0ePG1QJeK42mSW5QnkXsD7LfidnSNhKr9ahqZV2NzL
aTMalahgLse2sLT1Y7p0q7F3yOox0iY8eVoHLe0V6LZviB7Ek3dCRVJvB9BPMeu1AojMi2fvECxD
lzrksijP2vS7tz6Sj5nXhwgQdA8JIGG13hCjQVzvoxR0tNXrtvq2YABucBHqZqiD7So1TGKh0M/N
rp1v5GO2P6n0xO+fX8ibWfs4ZqQX+WGZfkmhKV34m7PnqkZx15ccwzKXblQW4zXrTEP6Uq1cJqHH
D0kcQzH5U4HqoP0cIt7fsDJ4SuETy7hGtT5C33KtjmcgSDKQKNOlehATwnNg+ITCufpAHZJV9b5m
vvx+Zp12j2qDDW2n7MHNcUMOCFb4QPcQ5CTN8xPvGVnTptIE+ZeIzlpczwyGkkOrLtRRZvw3ehbd
VLYyLVLU9MjdcfG9HmSmTn8GvRQrCMCVVsgr0mfwchHlMwZ01gkUmydNdi5s8oEOtgajyNSnui9Y
2NWv7gONa71KlEggf1BG3vwcYua/WU6DMRGZz4CkBeLwZSn0ww79Xf17gM6lD1qvzCO3r9TKxEJo
CsRfKJnxw5mcH10o8qCzoeHGkTnj40v3IpiYv70Nm3QIMIW59VlrmlEVrPyhzq+YNO95KhvbEPKb
81nDy6VSo2khi616cGc9L7ayqhm4/kKfoFUERqCUnMQeo8B8j8CTQ5v7REjB5EgPzDD27Rne8B4o
0FCOIyP35ysASIhFhv6i3vF5DztaIbgI+ubIh548tNYowrMLtwWBECVYA1sFDmBW/gkskXk3RLYm
enlV/UowWnBWnDKg0bYMZdDD05/QSv5nnwOyl19HSTNNMKmSQPNF6edsnKz//Bhowwt9as2/EPp4
sS1GENhXsiG8asewu6Be7Dq6iJDINSQgJZB3HVzFFHKCY4qcMuQCkXZmC5ofXC7tqRk4J4CP/Tgf
whVlz7qclvS10ePNrTDUfK7UaomQrk6UWhTzSR3dGmCNPrmdJ4TNAf3SysBOfeRlYh0YwT22DBEp
108lQDeZGNNemfV8nepCJFklw7IHb2jjPtVWagKRR2QGcrSWkcEKni96qLnCsCmNi2YTFgshjg0R
a1Ts3IBz1Chi2Np0T9auy4hdvJ5aDANZvNwK3Fwi9AR2Gjbn3uTAgxlLU2hSYGXQUKBcqr2PTrms
O4tzP8jDfXuoYEbcZM/l0vg83h82qT/NUfM0Fmq+IWXEvQ4QVI+4MtrUA3tziekOzeRURkyC9nFz
jWJ+3UBr2TbropVUXmzJwaOuyy8qp0m+XxfdGI39tWxskbmHslRWHmJZTCZgfUGHolIKkdnJ37s3
hcyr29VMXPnV3HlXK3hKC2/B3Nc7/7SRVn1SxxHM45a9tSNOd0ATcVH44N5UJldh+JISOS+r26b9
qnMD8H3++IvE0DvXffU7iFVjjbMwclA3Kw0L3t/3RVwxOHXbzRU5pbBf3XdXEUZzEAD974cNhPst
wGBTF+pCLluhJJzGIEiXZx5gi90nxhY2eKejS5ND6AVOf7/iW5Fe7NTULfGw1Lbpqjn8zBR7lav2
qdEmSe66TPgSjdfAh1X5oBryhsp2GY9pKxv2AZsEyrJyXVjYOo24Appdrk5cZgrSsblaMo5Xd5B4
B2FPrg4AO6F9bvCUH9pnW7NJH5g53JzuJCWZgzhF9LUEk14V81oPptHCB2IP0RS4ymUEIEa5H31E
c0XlDBe6E7MmGZQ3mW837Zxk3Qu/LY1Lu8PUGy0yWKjZpynM42vxeMd4VZ+3DeZOqX9K5vSSZo2O
UmVyUFZBnLnW83SnhQ0QDkUZWH3eXQM4RJzXbfpEZgf/rCcTz8G6qtwLvnEF4iAmHjGYgr+R7BGy
Xs4Cs6ifQ4d56Z/DY9OJEEBn8Vv1AuhqkHK1K3HYXZaHGJfws/3yThzKseY20HEFOxwW9AkErX4n
Mj6bxLIxjRGSeIXDRQdFqbie+uh+Izy7IpyPcCt/PORJwcBL7TJ0O52DH41FKLJ8ZUOnn67aYT5E
RITlSVJgRG6ey1K6n2RxKJTf6ZxCXSgD1ZGibTkyo2mXGmWCQ6dMB831ImHAs2B0XPpdsH3Su+tg
1aiM2OoAO6uD4FsS7YyDgdDnP7ePa5zAY4e6fNv19JPAGYuqwhpa1W45Fh1lrlmcBzbVY6zWqAsM
vRLvAi4JtZQPj/mnFYd/KRLO100v4ZdciJHYYeDGTtA/aFiNUhBBRs09IrQuB2a3VGoXocWBIgvD
vXBkvSaeMBDhhGJhGFJvrsRwIs3XIFDApJj/AqQU4wL/Ki6cAQSvdisDyWFfZ08fRliEobRFQtbW
XMNdWx3YHTurPGqgagnZb8oL/lLPIooOs8h6MisVxE7YuTFtwTY4UOmpZD5NbswEz9C6eGiBdtZe
7U5Ui/+xa/QpxCpVHBbExv3TIUWoaLQkyXhRXY5MpNjjAuG8VjonXz5poz17sdOg03uSZII4chMK
AlZlgRPoHUOCRPIjrAVFPAVC/esU5OyZkJvrfh2iWqQ0olzJMoyI3uAh7n2xVY//bY2XXt3aZ3+J
d3H/v9aVVqynT2pHFR7VpxEOsBfFwSXmacb08QGX4aDLSE8eNa3F8v48dtnUEb643UPFZMFcc0oo
YljJi0lfOjajsgP2ypAHz6Ulu01Znyh9y4yuCe2/z1OYHrBh30xXXT374GuhtsuRiPtyQsNLQ44J
xALvuq/PP3Pqz6vDdyc0TekzrkbBmgWvZV/Y9osb0aiV2I0BzPTK9UlQjOtEJER3MAmsWxwzLIaz
mV1lwgzzKRP4XuEccgjAsuwekHHAdYnP1i5JOUVMbFSwlg2gMlQuw9fpsL+0OE/6SsCgFRNY54WP
psbCJhxiJG+Sr/lMtOPJ4UFmYPjTzmrp1uu/BWUQ8fc84M9rUliIsJDSfboTIeoaKLxFPVTwBLdr
Dl6N2tIXrMgpWnoYmJe0J/DU1he6hBD4fon2YT+sN3aENyNvdpncV6Sa00eocBHbJqE+AIdaVlAF
97YIPHBagKWnGl5sO9LHhpPPp6AJZyi4j2oA2fkkqWByFZ1ZpldfC/IuszlDyT/yZrb9gIJLYybT
m3goUBU9kx/9aEai8hNoJDXbrxX3bA1FMybL5TfwwWJXdZTeY262hhs0qptKfdUUvO2ZxiZpDJE9
k/Xij0QR50cOwfz0+FfiMZKbCNTUNRB8Qr0qtElX1t0qR5927j6ELm+8WvCLtmZ0OqE+hg0n9x4y
tf/VotcS0yC7YYiIzQrhc5ODsarfn7QBlIn8P+2PmaNYDZ/3q4TUpfHwWqT+OsbhQNjHPJ+AkBGt
Ba/vkIxUvwMADof4RsObPRYAFKbmrj65PRaAJh1Stw/s919pMa1NkH1BdwgCnRqwlChmoEqeLt4B
f5BOzlQKPcK7pmY1PuMb6iNF8vQ6Rr+7ZC1rrQwCBaJEeIYsRPHrtMouLuqgRytlupFfDldi0ER1
NWb9vC6xmMj9sVy6E9XhLh+miWYVepCcmGMS4eswaUJgHlvlwz+vjIBovOt9pYvCblgw8ck2egrV
s+g/yjyVsWQtFXpGWZsXCWbBunBHSXvZjNSqezOTeNWly+MZT0y8oZHS9zSGX2mrTqufVKRqmubT
e3yR+KSPQlVVpVGOzUiB24oaagJTgYJxpe7Seq/m2n1s7CaOuHMqQLv5tABQsy6Bmf/Cfsh8BbU0
zA1TsMBxPQKB3NrOefebcrWsSLY+VWR0o7opWTA6q+fgt/Z/Ld7b0nkOMeph5Q2rhwUkpP9hzlrF
2sOGueLfYe+8sPLkb84X4WIHReleZFgGQV4ayzWQkMhXp0NlRC6tghzrNa+c2Y4hYoP8IWVdwsw7
T8ea6mVHKn/8w/PvNTXzYWbQbsbcKYGJ6teKFBC8Jm+F7wHPrSj7rRpeSKGTI4d1FM4CT6v0Yl1n
Ip0OuvrrKZtIMtyHY9zeDpZpEA/Qkymdb3SWt0wmcfCoZHajLk7v7aCZN3jLk7wRN29nMrf+PYaN
oN5T8W3WnbOsmZ/sVpkfZwVWaeQBqNL62jDCb78lHOFfaX6s7Br6FXiWfscqQIVK9l8u5+szQG1i
9jTvyJuKYnEOPd3aTTRhiQsgb5oCYmEz+edpsAstD9ntKuZ7VUG/CCifezjC5RN8vBiZrDvphtjG
W0yjb8xReynoZQbZkjHU6DGAYg0jJAi6SORybYSPDZn+96EyinNdv3gNK5KFnOY0pDNuXwNSk66r
atnWj/wS2Qv0mtlpEh7z+vazlV3SYWFAZ3cby02iQDdnGpw0Xchquy1jPIzGXgCFj4Il63qqK/Q5
gmeBnEzAiQW5d8YY97p5bZvvP79qAgNy8vU94t6MqazkWA0ka0R7bDkvywxVKxWHknmvMZQJMrzK
6WTV1ERQY1jdnPZskHqxYfh1ndkXCmWLRsd5EU/cwaw/PZJvnHgYPxI+35cVnpIat3TVdK3MLlj2
fzLXO4F/hhd2kwV6Wx/nCJqgHekP8iPnAraoq/INZFl+EFpfw/F2tjJepoIM4Qb0olv2LwRxI4R4
D5JnFhJ0M377WNmIoSX9b/ynmTba2Qa13/pbxhtCbPIvVeUcSDDGReP3FWEQi5xIg2P3GpdGmerI
876hfwhs+9rvuXi2HnMkmF2vD14kiA0S8WMSVZNwWaFkxW+uVUW6v0/fS7yjxMYFfXxritdvxVOP
pnS62w+fUch4IDHgc8LnRzJKDL2gHEH40z3MicHrvoIbBYwKbdgl1TMb0g8eWrdhmVzmQYIwVJ73
rsNp3aDDFj+RFam7qDGWTY+AohZ/KscKGrQ3qfsJXTQ9CpmI4vt9LXy7knaKHLdcs2sfbanbAl/d
RWCEF8SXBxHiKN4EZRuAhEbyXuuAjmoaGocLkFzwGnFOpfMTInnCl8kqBEo07Q1zsDmCz1QCSrZC
S64fVKkfuA5t7R6j5TBF5GPb4IhXscGvhs4Z3aLbt3R1ndj/DkKVp3Qm6UkIDjq3Nq5DT+Q4YGL1
iIRNN5Au4Nax3QKEcFeQsDTKRvNvbGCGxWO05yGbU2WnWdjVNsoLowOlzu2o4Tcn0X4qHUUsxqhV
jSDZrQmHIILGk26wjWmXLCynRXfhJOJel3gbFkYV831BxN6cyGB3y83uMf4dtJ7z12eKyvo+H7vx
fxZBYvuryVqORXr8nP1tEE2RE8BYxb/I0tutDDzTDQ9NeYM36VSL7TMyr1ZTtS1oXz3lyhbkMeKd
207yRf4Ep4fsoGcTuLYL/eclCEytq2y0m8RP6mauZ2WrBGJxcPonaRoaCq9DjQ+pwePggT2mRcKN
ubvZtZS7eS+f9Tu/ypkrj1riafK7GWyrK9wCBLu0f36ydkbmXOJwN86pRUyiHOFC15SyqBHrSHtE
BuvRmhbZYsLEEFwhuXBVVB5N02uGvmNvI/15wvwxWdDXM3zrQc3NFpN6O36n5P/Vovz3Xm/hjU0k
aO+VthzHV6xk+1HkSq7crNp26M8xdT3RKJ6zZ4k5tUTLctdZ/Zet9nqRozS5ZqkNHtasRV1z/o0D
P1p4HT3oa5Fs1J3T1elnNj2rPtTtwCpYgJ4zAB86ZIREKqhyi1v9sQoxH5f4dWp8KcN2rWFwu8ij
7COOtq9j8O5g1QezBFrtUp5Mu6Xd0aOYj1Pn9i/t4G1CpwqRWutNZ2TZZzkbsTxwLayXdFeajxol
wqe/QfPk9snNsCHoSVebAIRwukOslYvYFyzvW0gkLlmKogsgj4OcHBN17uWiyYSGJbL0ZgDSB1nE
mGXp4Nj3rGfudOmrRFUhNG7f8sqcM5assCNakzvC+32wH2CEwcc3P68Z9CYFSU0PZ3GRF12sCZi/
HijfAAnHwI/Vg3V/tRTcGrtoyseiiAkXk9zzWwSGkomZ0ZHNApf89bQo4pBag6M4clKreiqDSsOj
ziHKxZWfNO5rol4mVUzn44bQaJORl8TkTqU/kQQlnKHv+Z6i5BO1wqc8CbR4u5dzT+oHpIx4XLoC
Q/sajongVpQOUVGUD7IFRbhuTWJedshX5AdNQ9KbZw/O/voq2qU0+V/vqDLMF+r0zLXX0c/RIIPU
+AxO1bufFOHyzQpHlmuHkAcTfBOL8RAjh70ZmOS9+ILUbovbzjA9UXARPdnBBH/AdI3f7mmmDCpt
ijp3uIRmQIJsmkzsMJ4eBHDii1fGDUcTXKDdM/nDGpMQFchtdNUmJ310gfZiqZmE8OB2KeXTBZBm
G/ldtw6BQRT1qZkCPxuX3tt6Lu14CCIsDWFqjBbKiGEXAXtwsvjRBExXSpqwMr0im/DRRUW++5Y8
p7lpWXkHhSMp9cdYbROmcQlOGgdQfUVCyyjBewAL7XtvXJTuIi6sxRnKoJ5Bf6iy/CYqgTG9H95/
Ws2SRorXXY15sUDirJiDKLWQXHf7KSoOnt5jWARqErzy+X+pJfBqqb4OXhkEi/+9mILmVM0j1yfs
xycW50qHj1zaT+AOPEflmlPnjohi1d0oUtSDGJgAGrL+reu1RVwwmgWD3yNPQEtkm9Rc10fmfE50
YIdYnBW373KBhAbboEeFEMjEvJElyS/Spqmu8vjwjvhKcJDQgU46477Tcd1tcZm3jNk2G+QHf+fI
n03WjIUn5fWM0k9L9fcXeg8iyjAUDGc13cbUn6P/Gf5vlNfY0aqysi7D1U4GQi83KhxLHQukUpci
wn1t3xJO4o/gkhFvbPzprPspMWv+y/gO0RnK/QlJiFtsUz0VDM+8ygWYEZV7FDPaPvkeNiVHrAZ4
q42TT5JOpBUm6lky4lx34ycxKMKd1oLPgy8mLcOWxT9bcvm+hAG0157M6yAcSzeGRsdcZ3miWGO9
lNEhUAdSh2Lwk7oVU7IuwB4gkcpvMZMVuKhNDRHt+z5Fb+TpNr7aQXZ1LBnc2fO9OS6ufj0K+Mil
Pwbfm6xzjeBsKndoyfIAunQXif6/QNE2QTwOi/a7kHQVAqmi/FSxYXkfeYOCIis+HzUA6Vtwz2Kh
kEkMLDx6Xj6/CnCyTtgWMzM40fPa/PUbqvCJ1XOqFO7GgoseOXB1xikdzE3c/puBJvTwghps/fYI
gzuICue8Sg4CKh2LrBcojAz/FCRxCgSswBNK3kVoEHiJESFMipyMvYFf4vhn4lWuP/q7Mrdw2xkx
5vCS6+NNUg3TOSE2aGLebwyMg796INeJioXlrWjTooKuKrZwOmcWZ2sP0M10KGKKBch31PSidnMo
Bn5fBop6rexQlNC31z/NeF3PBztNbn7RtGkGoXumAg23RJpzsjnqR22hJoqbXaHYhq5zjuEvWGDT
C797G2M3tNFaFqtweUIvo0y93UBuehyGZF0Lr4G42E2yI/q/kJCreDis38tVB/1+9z3TU+UubVe8
sH8FJbpOdyzA0lEu8D2CzRWv0ZPLLsQWIa3W5yMsNmdDcb/5qaaPeaPr0b6I3iEWo0iWUofuY5F+
Yd9prEsnDHTYHqqYJu9VV4bydyx9QE0hhLHDX82hqxwG7VWau+sujN5zTtD2bQHI2Z8D6TMBc7l6
/8XEfSFkfr41gtVoomq7M+odE1ujpS9rTpU0u63mWZPS2a495/IH/EfXEiy/SYIehP6c8TIFF6a1
UWMvoCJJwDqCigc12LCYzuz03trzWdb06LI32EF+soipWR8e8shW0l1xf0BWwTGTYeGll1drPPNB
bIHrCoGzSGssIQr4FrcM0zCezdX9vaeBMTIjaGhI5o23N9IjISFl7dft9NuXPoyJeYPvzI2anSm4
OGA1kdGAMjplBCMgaFPhX9Om3ESbcWLEynsGblkXZqVZrtITKLxpLwWJ1XAMqmqFoQ5FmRNrJtFr
cTdSGkgmFKV8WGHFZ7ICqocdDEBOWu7w2gSaLvJNTeDvolDyYwA4+nVgy0fEBhjY7V30xRglRv6L
sex/sZnryx/CQwgeAeAY9sYvKgUMnKVdS+5p3IqBzuBXquXeoJoLrNZZUEzNrImhI+g/k1Wo9DIe
eMhAQLmRoWgj5dW28or5DodMH6pd+W2/chESpay7qe8od9meLtzCps1kRtM7EXyWspRwXP5cZNg8
GT5gd2cwPn+X+oOfjZE72gsKvAx6Lnu3WITqCUtlWGHpI5g5C+rEopGfgDMecsa2wACgptxm+EU0
ZE5e+47hXfGcQI3PHrdw40+y9hIDS7SogH7SNB7Veplqg1qdbhTjVFtWbWwKTrKm6JB0zQXP+HPE
uLggLIXRouwkpFkT33RfCebj8zfplJtNPf9EJxUQMZMEAbVKe22HPrO1zGRlRGzN4jgSnQOrh3sb
YN6ZPOIGHte7PJBZmVyZSDbimi7Msjuth9xaqBmIhum2NnCB3hYp4XfKvqVrfG8JT66hyU6P6T2G
VuN4GokjTvgdnDI5URXCEiummfnfXqmbDsiVr1yUxN43wE74naOE5/8MjkpEXSZp87TqIzKBZX9S
eE+680xqKBaeEeXOD8yerzPaX4sbSdPML5qsnuJBw1fS5VElw0j2RgFdCg5IHOvBhBNsOx30Yoyl
vQHF6mL22yGr900BOZWlpuc7ySp4eXIxKr8BotvkkyLNv/Knean4KmRYIcJgXqmtcnoBvh/nr/+d
5snrMILM73MIeNq4hbx71Uu+z74Bth6gp9MTYnSbsMLTJbQQSW35grLdKtQe1WPmlh2mE74GOCvW
fM4/C5jCFr5DjgAmXzxDb6cLp3of2gUATSFDiAvZao/W45/NS5sg+92O3aGbD+GJdFca2OeofPsT
WguD+AekliLJiucU+wYzGCWcaFSBd0hMGxXqSUoQRDwp3PNLapgbFZfBUqU6961bW+iRfeUNuNP7
S9B+yu+gMhY53xwZrb3WExLMtuw5XJMODhmRsKW8AUpZmOTWOWWgmKJV3myg7ixQtZImxULv+Jno
RWeMCKnJZ8EVzyvCQtZGhN8W7H+VNs+xTs9TujvX6bYqActm8yMkahKGIDQ+mgBCXoW96pgJ11ic
jXHsdmE6B/BhrljeyZ7JMrVU0PCNQpvFDF35CRA+o21Oyfal53VKeZSacGLHzGhVrr6zueu8sAsl
RfmOBGNhc4iMDHwEMXI/QyAPvMLLMZGKDB7BJaPwcJdhrOenvNhogOWp7EkBQlpyFeExBlfrbxJy
lvWV+tXg1CDOw9OssHBwQFthKMPS2UTAts4u/xUNUfDbDv+4TeclVmRT0cpO8MDrcX62ubLIAqXL
m9n1uEX7i2f03uJKEh2qNzLwMK/PJx+PzMjTqjcVSqD6wV+oszReAeQFovD1vo4XtgQoVEuG3nHb
c43SManbbLVsQ1cJQr3iafQxEhL8CYt7zS0edlwEIJKRlbLqvZRsuLH6nE6Xf1W2jT7kQM0Regr0
j0HI2uR7mblgSRE/x1MHqkNFKUH2BkHg3yA5QPUFK7s9qJKcG6Kbi3miMoigWNYB62RN507eHByA
JuF07Qo7mMk5+SL8d9rI3nFDF7XREWk/IW0WnIX2+I/AjwaeSLd0u6RB5IbVZsFJD6ZOf1NOmeiu
95N51EgaZFak1qIe7HS6bIBYBbFj4VEooGFXvYc95pN3kz2ogzHPC9tp2rSKON/4zHCe3g20hron
d1gERyJtOoOJ7IpdEHyfI9BRGEDdB8QLvm1VWD+dj4VxM7ADDJHpp0txCSdOwC6w1QoaUQ/idbKz
NBzaX/2YFhGxyjwenOSlsqAwt7s8BCrbwal2sJQcNzX5mNvH6HxgL43iwZWL74DpwG6qMNNlh4PV
KGjD796g5kuVwuhvtupipnVEzSfjEzRnm2toZSjGszt3RmAYTOQgTC675fZ/1uwEF1NguU1D3qF9
eqwHbtS3+Cyd2G7FQXAAzS+vYuXz/kUEGm9KMx0UJOvbfzb6i8GmuMrx0bLS5UkOwWI5Zm1KhtF9
/swxUULjH2rdAO5w9SrNBF38kDnrVojMglzp4jsLgIoh+/zZeYh0Wej5twPadwcXNUBSAs4NHdhK
MrhPa0ZBNHH5vS602Ob6bVO+SvItUDEiCv5PvF8Vr/ZPf+89WmRHkfa4xwtLwHCqdYbAdtvSKKUC
iFqpH2sIbRia+nuXEwd/0b3RU1QDoegid980hloKIU+OagdTbqFj6VLbKIzsaKIUs2FLdpTsjVQR
+hl/EwSQAvomn8GixrKoJjd10PUEVlFgtC4aKsd32yimlpkTke42YznVY7VDNQqPBP1m3v8wE+Im
Y05ty6Tcosl5dLbNk1OF+vVN/WLvHmcv1uIy0J+3OFqJdNZXfTUfH9auYL9xLGLJfBlPCL5/hqp4
P2cZ0z4MDMVSZKtGJlPfs462X8v5kBjrJNnAffSBhxEN47fhHlFCP9TKKQU6klBI7gQgvzVaQO9d
P+snZ3DxDDuEU0Qg4vbqL2kpucazdxMT6d4GuWaAB2YRhMcaKgQ/5pQvU3/994GIbollUw3qVRR1
9j9ISHuF4gnkla7M5jT6E/35lZFgHN1qlZX9iPag2NIcouITz4SbbMReJoTI9guGkTBFYV908EJ0
vT/mH75pvy1IjNw+/10RvFub8LPAwxn4aTcp/qWcEJV6dcM+k4RVOVFaDeCJ7dVouo89iBVCeJlv
tqseCr9qdNmlEpe+IFsL3WsfYhP5Xu481dKrD2u4mTZQuPm7lvC74SAhpuedxw+KikHPDSZ0TXWU
SF4mh/rmt1zl7qkl79TvCpBuHqBK80/FI1fKTvrCvXsoseynNKYipuvAjSxTZXfuOKwCcn4Kf65a
vTRhcLF09BvdZCeJd5E25TSk0n8jLsugIAaAnDexmtzvMctvT8NId/b5FT6qUJKxeybwzo0RquLX
1Kikw/n1Z77g0lMh0FTDpje8qEfiqmcfc0hKcmJmnO1sHgIgsR/ehAeslCUiijZ8tvnI8tnMxDRh
tV5KxqVN/mwHVVChbCnoWdNEgmberFwQIMIw/K1nYBOObmbgsewvDZTaasc6aQNlzMB62tV0rgnj
2vBZcdtDEehsDSpp1PHsRoDSRmG8rjl3qPU4xU5nVn0zm6qSNXADOETv7Gi9Y2xfvLjQaehxs5Y9
tojuh3tK9JH5tfi7fq/c6lCUxShPVeo70fUqfWC8Ys4WReTm3BJjTyZP1AonvWCGlPvwYcAEFlhB
PfIG6DuxeOqRb2jCvJ9Jw6BVRRq0RVisevtbjugtaZXd+Wa/dPl9QiKWIeOtORC1BDYExgLEntN3
Q1yd5sZBR58+DzWYwBR5qlSmHKczey7vOJHk18ams+KRYM6QEjmJInPoXlCtv/Srg6eTekqT5TDX
0wFt+FkVRSmk9X5Z9XsjcCmohvJ3HNwg2NZBgzJ2H3+5n6UWSWaA39TZhs1nwwUipajGS1NzsOp+
r4X/WdejL3TyjQEerxfN/9w/Fz+Vj6HdOgSTnHoLVMKCpxMqt8FvlhKBKQpNwOF7F+aZ2R3F1+3R
CqkoXyxzBMYdaF996EaG84HlZhQpbfcZlRo99EnenxtqhecuGYblm3F4dhePZaq+opakzyQbXz3h
wDY9SLW6tI5xJ4HHesZdwaQ9b/0QCiXfXm8TazUT8KXp+V/bL0XyvqWcbBR9mHS2/xYA9ViXy2y2
SWaHLe301hbM6X3L5p3qdxv+70yG70UfCNK35X5YJkr24ifd6csisf9UiPQwa2h/hkEuY/U8CP9v
K6ZZ+H4Bh6TAcijaxYNQ1YesYNxOPZVyS61I2dAX0LH1Yxo/oRi0d8WRVKxSSA1092awFkc9RjVu
q51be7CFK3/01Tdh9vW+a5Dj5UyI1w9W4zupdCMxwGXgGZItldzqQzukH2k71J7N3CsvicAbaaRC
RInp68p5XwPAHEyCYCA2YAkdL9om/wIYkrhZWlHjxt3Gt5bHxvDSw11FAMZQ6a2cujtZATGV3dCe
It7T5NmZa4yOlh2GnKXYN+G/rAnABuQFh178SSPPOTfGWdezY8yECspR0efW56z0Pel2jGHeg85Z
MCM2x6dSFWWw40xcVRm4hM4ZXWQ1Jf85dj4gsZwRgBgRXSfY9a22AjSHtbEyeut71bmj49Neo/RA
qJhigaQAzk+FkElKVoRRMYpi6Rr1TcaEqIknsu0DerIT3uvtskwFaMQlMGQivQzEon3yEgiwVRP1
V+KL3fIJa/GmUlq8kKi5LiYAs4TO5rpRCtSENaf4tbBpfwVIM7Sgd+IrJgcNLtUXNFtvcTorxrFA
Re9wZaYdUz9c+i1akKxelk9B6jUkbLrp6pGzRFeFH7S7NEUPcDSJA/2m5J3+D6xA6E09N0PP+6w+
L0UKsIZeGl5WF8RQ4UoPCUvZ1cyb595jk9IoXmRXUk/3pZQQbXHS6s15OPe48/2Pi7md+NVpQLZ4
w9qhohKmizgU0RvYg1qowAr/TMgbNEstsjQ6VszwkquBEtlz8qe2YA+ASeWkmuljqeJZgA5wA7bL
nMPqu5J/mnL/dP23Ru0h/Bonb2opdX1YcMdRzfz+btfEHUpRc3eHKkaKYbEY3Fyz+yB34J5bFRMl
G71i8AAyRfjpvZ9UwM6SjI8LhY8Xi1V8SPS887L/acDdEgvCvTw4fXjv9zoYIt9D2Z9k8T/4VBSC
KR9MXfevpoRTiw3h621COxLBSImZ2KjkZEGsHtZfvHHilXnxxZnNInEPS6jQx5xZcGmkQI6eCl2c
iFpfVu0Ibjc17DunUfqZbPw4jHlBHQ8TylGyFOJKtc9n3SDqx+0XEoE4TFUDGdzDAL1a9dzkzMFg
vAI8q8HFzOxena6BCLmqXoM5viQq13ovUP1Wr6Dz0G48LruCg+kvBEa0DUQhSej9jhN1sRaf3pW/
oWDPqB3TY+RquJd40llDV67kLp/OSNdkqeXzSl9ayw3M4XlveW5yF2TeWWoYM2B/RosPR8+6CKSW
fca5ji+J8COajG6E1oCVOEgFNan2le7KcQ8hH/gmeBYUyoUclfNE38zOTOWpaSCWlXhclSo39sGj
oW3RmUNKD5evoVNhvvvUz/cHIrEeSsT+Yt4LxAoEG5r0WJvTCVYQOuoSwwy9RzWj1V8IyRAgID3g
Akb3IgRBujeRvs9s5UoTGhc7kcpbklzY52fg9lFwLXh29aQO3xbJUdql5TH1Gd0X2KyFJ7kQwlt8
qEspKeUj9mG0Yb2YOZUigbuWEYXCnskJlxHup1myo8RZ/t5R21GSDj5PeTTzblT9f9u3aYkAHLxM
zZ23uQt8FmpPBPJyxwKLZRJBzBYKN6HNCDMYRtPBYfbqLyZXq+AY6ntI07L+U1jtaD1+w7gWwhyg
3HLT8MIQGON7U8A6D3hyh/gT0nWyMXMmnxOMx5RrFVWweULJqF4u0LKDTQEG2lobecj49/+zoR48
8shoZkIGuISg5pXT22+oOYYQs0X1QZiJI08pMNCTmxQijYGgqiuLuKofTsC2Z3Ynf05giS8x1t6I
sH74fdDvvTZ9F5D5gUCzxlmCoetl5C31P/pjl44gm0/zr0TYAf4yo62/hV46YoGHUobBoN+h+BUe
Eoo9KB/CjW5RyU374IDSlorkpTy+GNdIEChyTKp71VSlddZ3kFtvFeW8IpQOyoCJaruKj1ii/Vfp
nUxSApfIRbbtVf6bOe+JopYbs0BmB8bzdvqxHiiN/5Qn/vxx7t/hFJV+TxsjX7zdMZnDL+2BgdlR
gFnL+UOK/UOy/ByIqlK/X1e+MS4iI7cXbYlnh+LVgLy3bdCJ+NmS5xTjKOt8+yS9wZJjDppm1jov
Jq++ypb7aHcgNcW+4HcQiibWpi3+ii9v1uDyYjkTHsXkTlq1MmbG9C2+2CWo7gRXklx5mGOleR1d
fcamcEWZ4hkHFceQs2yZkwNGKb9/axPoA+hXLobqS7lH6NSTJ/YUuP5qHujQzrkX64rrZsivd+89
hzb4kcOO+/AOOVaf1pwMSnjTzpWMvFp8Fk8ou1CJKyAy3d3Ti9r4UQD9cVIZzBLNNrx+MwmmPWrp
xmJh/x6UpubGiuZxC1VW270MOGI5fT7ZGPECT8byl92ilGSlyJbZGEP7/UxrXEf7sBN+8ZamdYRT
Q/vYp+m4wKKSv4TZ/l3b0qlc03LM/6sj0AE4u6ri1SX/1MufJ01WrPf1+nx3OhsT1M1xw//C2Hyl
qYAI+Z15OzC529003VZ2tEenodLz30lxOT9x9WWKz+5WEaZA112EyvKPj4dKnA4CR/30oO5Df7xE
kv1AQQWK+Q+zZP9XG2+GFA78PWnJW0pAmIhNRSwvELEXz+143mI4Y2HjcCulO8iWc/iLyTZKLVd5
fOG7JXCvHc9nMdRjKwFfu7lSDcRJ+Ymic4xQt5vkyPfUg4MjDWPbRAtkMC0WaMwNWtBKPM88I5jD
WK6+yJ/E2LmM7zh0e8m+IIMhlZNwWYZzXR4LSGb1m+pC31M0hcZPdvJIXlEoRw6irkmHZ2zqAaI0
NEFc/6HG5XHCXrHOnFtTFvL98FomVSU+irSCjcg3AKVztAqnt3MGxk75UUnlE13MCAykA0erlSN1
/P53jn5w2BX/cBV/tDTwiZyVEE5qzLL9Kr945ATn7GT6ZVZMQTh3H2Wc7WPWwtwt5LF/E1z38tzM
JNKeWbBupYXjmk+Z1tJG/2jXeZ7OqZhSXcW3TrUEbJ1QRdATLrbMwDSvs/sjTWwQuOJf+6hdpDrn
AlbYTxXmmpmgTzlz0rxLV+0vbAQGEqrAsXLudpR5iT3ypOHrY8uKxiRkGTjftbWlmxHgAveDNUV7
fUc2iqOEmTgAuZAsY5xal/nVh3ZpB29vtxijydybMJICevjcyJ2rUdOJse/4QPXkPsjaukdogAFl
ZT0uj/tkhu7yGe0wHbMJrW+PvqTGIT8HR5Q8dYKEgMeS/LsrPPd0qKWLWE2ojU5K+9UNJ+otfQgu
c+KuhOVw9AkdoKNYMuG7Q7lIPlYs+knRLX2d6snSGyugjOIB9M496/UR50aNMgAsi5o2TmKx900g
CWeZSQcXwK9A7TV7xourOT/COsk37PQyQUKuJrFZ5r4jUdr4HqaqVYo7EJY04NCjKljhvmbpCEIQ
EcCPnrCTG9osS8suonbI1TpBdzi1vTzFV9tdD9OaAakEls43Sl+XgMdTY4LasmIeaIojTW55dgfi
tpICfoyh2lyWYN4JN8+Z3iiuOZPg978w9dXy9n36WwWZ03nz+Dw93J5VTtxYVY+Yi31Iu9Pe0fPB
eGYgS0LVGC3eg2P+QvjVEVb5xgGimGZ1LJurLvn5J7X/WGahRJvRuznIGYUbAh6o8MLf2AvLcGL7
98RtD4BFGGwzwnmil+HF1XX1VbCzbrzn+2+buYjDYefs2J4tZ6A1jS7LQTV/6zXBUIpegJcvcGOR
LL7Zp8fedNIXZ3aLSIMYXwR1r0nSMMNYq/2rJH5MmakolO+CHiKLMPWUzhJWfjrjo84X1Ooj/t2O
il6ma3/nAWtbhp4Ne8R2sjb5euB+v4ZCdYEYTe0nYQ4rcodyJQYbzqEwzNSdVodM8B2ynyIkloBr
gIogboTZ9QXJ6PRWUXZlNAlsebzzk8G09i+ll999QRnwo3qih8Q9Srh3EjqprlHACmXyfCfvyi4B
yPWZ3s5LbW+d4VFRcb2lG630vwXAFMTJCe77+sJpIhah9gGnbbD4sPuhFMt1W58Y7GhHYg9MbHYV
nLbyMLRtClvULoiRo8DW+UeDoR73Ftu3dvrg8+oXIxyul5NgOvqRuzP+stPKnKWPb9bEzlGf1i24
M3fwxIbcONO9+a43XAC4L/SQg6aDhiiuAkSBeD3K2h01VMhUcf8BLOdnOax3IG/2wCm4cfx/tOyT
39cBfEiEn28yFKSVpRsjG3CUR1OCkNxFxvt4AkXGq4ZS6F3PPL7cDi5bnHhizfLgsAlfJnZ6yyBp
kW+KH/b4jDP9xWkTHrHwD+RsqSaBjwEoKzBA4Io2pByyEp2m8uBoME5Xt8vHhz1Fl7iklM7aWBLo
K3bOISXtc6L8GIKlMAsEN//R0pGkEOwBB8H+k8MRISU9wpFkUGiDXkJAVtPhPdIONktVvZgf+9FN
4oHLl27gk7ZNakXlUPcMUdtCOKNfbkL76WTSrN0TpBsMpTaiIf2/kNGNUUlv4ag/czyQIgQf2wHm
kHV7KJDWwV6R3R9Oa/wvqTT6yEBzv3N//Wx9ZS05CHj7ZiAKNGm34luT3Xe4kEC8YRcMSkHZZFHE
3ZXCpEC3GXFTjHwkEJjC2Hom9X/KLAHa1rcK79Iaw3UJlcY7B+n1PL14wpJnET5dNGQwytM49YiT
+SmXYGOZOxZ1U6qYqfM++yFap4R3dAb1fFmZW+Sd9y+Il1f+UPet0AY7Wkcs72AjzDeT7hSKZz/J
P5barcZv+TacvEPkAN2sw3Uu8coUwPSkU4/0ncNfHtEmh7fdIEUcgkmVIodeHXWYV0CjGbGQ9xsA
8ZyRRNCrF68E1pjpOc9NLOhASFv+iyJidclca8jec6Q0azz44pXFdzr9U0ikHer1Cg3DnTaSn0bs
n/pzWr3VaG+kWKL1sV/z/zOP6rSDnEqmmA08w5BCaw+zhYmScMBqpPZPFCQ8z86VaXNXCOZRX8gq
joqL8ARk0X5PXx7iI+62NcuLKVYC8nFcFLS0EEMZPhV2V9WeLWnQm+61R9eZuOCrrC+NBhvQwF9L
EoOoS403Vz0emwI9ptYVpUaDmwJ83BGTpdboS3MfQF8G3H83OXvNZ6YeWbxeKcqYLYtGhWKmuq4U
Hqn0Ck+SAXuksy3HG85KZZ2uzvQT7xy6W0ABQlBZwv4C5eYtUpCKvEiYTdtsbSFpShCbLq+D779h
DOEljCio12lS6AybQGy1GUP19l3hSG0R6Jl0G8ogBxZpznJ/dkNMC2ZinA3ihcFc6oc23SLsgIoI
GIcB9JoTE5zWZ/v/M0dBIw9NczQs34/TtOqbDzIYBnqDlgZZL8JVg5UHw89T5mzk8BMnv6uBtXzB
kjDxhY4RBRs9v9kWkQvxMncgRphRElYDQ6QT3xS42otcklq4azw+aMW2EV0V3qiUQzZ/e0RwwMDY
rIG4a+g7cDNk3IOneeu2UDTeCqxXvJ1ndDR4Fct0z4iX6EM7Yp7f0BSGBuB9+fnPtVmXOSCR83JG
IO0S90f6PxhfKsmQKOMnQgadNDZifdR36igW4utOhacHEwRC+IZZFKa9jkw7A98Km1ZJPy8U9WnL
PLO/bZhHdA/v1B2WixJXK0tAomXbt53gs6QArO2zwbuKae3DITAgVJ7M2qvkYri3OhLoF3CdKLNl
6vJXY0Boun3uQ4d1rjt78Ru9OGSWg2ItJ4w1J/KiB6RQHOtTWF6Ka49TP2mip7RGv2en/1kjpaLz
UwvnOUNlyBOFFLLLzxnmCmAe9ZYiatRiX9iOwQiZsJhtvlKsBAR2Cd7XW0YUHLhkklhuHPePlopb
gNDJXMX1fehqTGaS+RVxuNSGSqOfrpAsCx37c7EfqkQfH14uG+li7liPNJx0225NpWYU6OBmE/HS
IbhgXorY+2pTWFoAF3nAv/DIkzDd1CwTCwFZp2Sd61h6ZYX//SfkXASB6AnXTRW/jFubj2mA4PMT
ixNMcaDdA786tpm6MszE3ya/YI+wILXg+jk20kLOReNN6GTklnh88a6b2dL7nCxkK2z2/OWDWsmH
YNJ+ln/veg9am4ArsqlFymiMV/DtpVnLu9+MFXhdws/lMgrPOfxCJnYdGd9Z36fqMNG4QMlhG6WN
S4QcQzpCa6QvfSx2nYZ6ffC59L8Me/66RiEfEOFxjj4uvl6l9C3qWDV+hEACO3vlJdWmWRjNmvOK
HC9Bqte22ESpG3ZOfVaEP+yQaqO+6cCu7JH4kHvcfJ0e2ijR9Uu4Kj2gUtXaCeeqMrg16dfp7WxX
axMWe4E0Nvrp9AerihwMdmqNhFJlfufntKuuMcWf7m9pUgbPAYgATgaGKY7TeUgP2DjAFtTwfBPw
AiMjTlN70jcRJVA58WQbvzmcKi+i+ytBwpSyPNVq1KMuiBXlNXr86qB6cR5cQPHTZTt2ekB2XHHJ
bw/C5C6PNhWv8HDCuaJtjE4ZRLmCDFeDjbgxGmuOCtqlGu5W5KkQZQ6IsaSikos2mChGI0nPFTjA
xF0Cpj2orThf0vEmC9ER7SjmEkmuMuK1PPFV9ffmTzUNPh4dNDYvTzLnqWV01u816i3Xcc4l7oAx
z8Jxir4VhuCZ/ydw1C4joryiQOkL0R78AFBQ8mv+o3rd52bAAm/bHXtOFFeivX5V5DbhkmRUnVxQ
jNsRY8Pp/e3al9p5r7+35DFZgrc4gLZTmhR+FbPhNlOEnhjrZxdwVNN9VSJWIioG5+y7FY4NBp0C
D/yUcXKkZhr6t1QmkTdFwaOpey/F96XGEY9tUCxMsGwTRfjhC6zeRNRVoNggeH1BbLuW3WcQEdeE
fGxzwVM2e8hzEvFzTu0Cw1kyoQwjjkn5ZJVkN/3PlkGG/+VIafD8EWOJI5LRaH0JeXks/3nToisg
z/7bsktKXIWGE+ThMnIwgnRgNsmK7h/RS4j93/liJKuyKm69HOu281jiDLLLWZtfximWsfAK/L2n
vWfcaMIrdztlJupjphVcYRp9v/u4TyjCJmVbHYsbRWP1ZluFHdjDNJc8c1MFOW9wZerM9N/R/Ugg
X4QDYpKIP5XbjqXFD4XlssyUoVBEdUZoMMjzHhs7SO/U9pkc4VSVSx9PM7nzP1vG1SULg2wsC8dH
kRuGzUI22uq6muU6j6trx6rWVxhLFqZ1KZrj0nU/ShFb01rMYLV51AS7jk4+3M2PJZfDLPKfN19P
LkRUWxVv5QGaFNg29HjJT6749H93l7wwXoHPS3zrhgG/fcR85cHpcf3ik+ncjB4s2FMgUckEM118
jW2nt5OMZw8TH78YYCnhjK8hjDsqPf7KSSe0PTdJMK1Q4JYnEd8NCR07DrtfJTIhwAVbhLk3xO1v
A0VyW+M2F6dXAoN2k7+Q0qWX9fqSpR9IGuhxr1/xJSD98eDpD9j+bjn8U4h8ZD10XuCO73Cpc+3a
7RlVJdcsuD7C8RHBiWmsG0OdblsU2rE/a8A1qcX3kudeFk0+Pdo3xxsqfIaYR0tAhyDofEjtOk+Z
czYjPQaphhNkPyf3vglKB4Kl8WaSaQlhhGpIGPt1VUBvyGdRsdAsDTwuiIlwVfpvKo5nB1n1Xh8T
qaWykjMPskykqj6kVW4NBgBXq+g87uJ758MFvAon7mNuApuuASoEMV6Wjq1sbXOu1BIO0mrtT0JS
aWGL4AHJs7j+klAdx/V44/kpCMCumRZT2jyq3A1gkppTZAf200YHMGMtM3bSgondDTr/wqHvqtaL
su+4GdIJultY+N4ZzxWVHX6p0QdvfKTEtlynrvdrU3YtrV8OImgE6xgW73bkjUpMK4uy/S5bCceE
w7lGGZyH2FqVNw2qibuX/gD+c+FlchpK4JJMCX9k2d8oMz2oprLU4ML+EqjJJrRWyZ8ZiILCSx+k
0cqrA7WoZrv5KJsU5YQLFcEFrUZJY+AnX0bHbo5HLO5oYcLFw9eY0GMVm0xoSaMY2e+0zmUZDKwI
Cg2ddtZPsbCowhnt2cZ7qL5u0ZRzXYUrJsbO8WYKPbNGgp+M4x8cak9lA1Q68Q1Z+naOhlHcNq/o
wgpW+qWKCi3BZer9otyU+6SXNRQNqunMGL64A2sAVRLAVqoAa0EjBpv9HsdL1X86LBY3G88IqAWn
Drot3PC1nDkJaqYoEcLiy2l8tImIvqtBIP0kSafBc1I68t52XcAPDIfSjzCFaaDz84n9j1dx0DHj
aMBKB0MFXz6e0Z0fxuI4E7VOXjuCFwtQQOD9nuW9sADd+ZuyPMJWNO87ZWhOWxlrA6LNu0afivjs
mmUEd9gttbme/djnKDWkN6CRcTfvgQj8FtAf9Nbqe8y0jnQPq7bqn6Ye7mcTHx4akrL2WnzvvevU
PzhkWLAAQYnR6DgyTXEO+8ipJE5Ry+XZq6fHxrWyv1mNhdHrjlBl7JKgB5fILfv4SqgFwOcTRT4v
/O+XnmFg/txAjh4o581V3xj9fFfJ0lCzzwSvKGIFx2QXbm3SkwqOsPh3i/tDGj/+7+Mao+ez5ibf
C+PO7WnZtscRh+j7xQEo93W1SfqXziDuGvKbPDaI2n2tamf4vNIwPWUboq7h8dhUOab60Z5FC1GN
qi9oFrzHAiOJLX8E1Mq/L2WETw4trUNzgX1COGA0VOg9ZC60686ic4xKhEMgm+zVLpVKrrrCigFr
R8lef1LHNLN0M7ZjS+PB0Xr5VPVuh5Sn8pTfDFR8B9RcNo0/kGBEAHWs7VMfeNLrWPhi2Dv7IoI+
NaywXdSMDUThZHmS7FzdfQbyUUAlS8Ur9bVVhoDhjMt5mM9xv1rZEPVtqigIA3axLXnhMbpeniCT
RGCxOMl5S4SIVI5M+FPL8meW48INcB9AlWzI5dp+I2OhFv+xH3pmoQu16stGMYlJTOCtiqXL9kZM
J86riq7p3IZm7e1tqmDGnuLglA2G7jTcR1fx/CjDHyypKaJjCQZVRQLDW7wsNm+9kc71uN0n5v3b
dvSNnl2OVD5JOeQfbofJ2b1LdQQ5J4SGT54otPdEFnV7Plj10zlwvL0gb/7Y3DpSVd6kozJF9ggQ
8ioRcm8DiuER+eenMKC9rIjqhKNki5G2xuB/BvtbBcAeqBDibYBGQwnRdmKvc0Ejj1vAzGraV9WM
hlbE8HWqy8e3lIoKHBioY+kGhJZVSuE/8EQBR0ym/UwJo9djPdLcwd1QrTRdmMoKacs6WCR68ATL
G6cSPqR2aTrVGlGb7Z3hBKsi1HViuKqAlgyWtQ0r2x7NM7s0A/1LDj5JRW6iowY6kAi5dnKZcJ2G
WXtsIgLG6b3/26Mxp8p4sd+OAacVXmCzt7ObYzK4+qIXbQEVRqRpe/nmfiq3YGU077ZngNKHdeeo
RWd9lnLkUKB+cKxkIH0eiwg55yNIY2wzjGL4+HUSPYidhmHZVZAWGV2+Hj8nbcZhmSlJZ/g1Gtok
s9wo3lWIKppEzPJFe3ADdPKXeJlRMlwdwL0h7DaIHDw2GLxM4/3/fQGGdo2q5lqie6njFADkmJyM
q7lo1Dvky0yHX5Uk4WFVGgd06BZ7+lelWxRmv95YY+J3TCjV7xqjkh4fmx0NOpXN7b+UIkMmjYn5
SHSSZzgJ5bScT+fhjln1rd4Wm7qQA+FZ5lyjD692JRh50t56PSmVFgvvV0mwNOKtpNzAYlwEKhJM
EkKIEvTSAOIR7liu6URIrrPGwih2reqPqfpexJQI02rRTUyVLz7SlBpzk9iKbpXUlySViZu4CP9i
yBC9LuODZq4kSZQNFsTJDX4sOI7R6g8p2mT8NPWOWnex9DtpKOJupv/iLkAB5FNhBKziYkk3r4Wr
ZCx6VbRVX4VANPGS/Q1yboKpwEpjOpvjm/jHyfRKY7wLPRLxy8d7rzk6ahVWe+RAu5uVvTDQkvIt
6u99JfokAnzTzNMNhvMqaIqcwd0zwrwr14H8aSCPAu3YSM1csX84/QBXQto2GolN5JNaiJWCJ+DF
HIP4/OHu7ty8PYtb+lEl1BcSqcEZ0gEy5JOylpVTkqGfJfpRd5GYhApgIlzA9o/MDnODQ+2I3xhJ
LU/CaCeMhG7W6PZvDP/McZQR8UC2gRrpCBCoQrbBDBjZnyiT2ONx3z/gR5VJ096VTrX/foJxCCZ8
3mvxPPjwRCM4cJ8iRXI/u6KZjI5QTM9jYEPahYZTIxBNqOxe0b/a7VdVMByh/m8IO51bRK2Z49o0
XJfUtUV3Rqqp6TaYP960KiqadAcXK/dVqbp9QNuRrva+NPqBah9FearOSKLSB3j4etDnmwkNC2lO
BgYB51x97eiRxAQ4TzSSxeksMNhyI1ZSKIGzTO6WqZTJVj1XUj9jrFgef0aeWxrRHD8rBmajmF2N
yxl5krJiBSdip4Qj2L1g/bHQKRKVCn2jps7TUpOM8zJweUWXMFd6a4utHUmlYw4MR3i+P44uotku
zQ1XahueZqFV7gjedEpz5DinVM5NXTSyVSLjfX8+hp5KDXAcfM5RhjKdbn2O8miE5mQluFv3QMct
DRSidw83TZT8DSwZ59cApFruSRThMDBYkTu0UyEuChDsn4UYU08kbroIRAXhdTrPAQWqW/p7J6Ke
hRhwup26iCYEoE4OEz+UIxFmkz4VK42NHVyN788RLUQC4sx6fRFZReY6ttQzUKBSi+jUTN07jGfO
e0xH8f59HFGE+Z011ynRxmxxIy7rhOGBSNLL9yvmvckzestm9HPs3Vg+J8wuXEG+nHt3+BtBKjLp
xF+Zdo/a2l2z5NNgY8rowsEsW9tA6E/qqGpz7tCIdAbSdeGNrBIQAZfTbqsU/7PmgcKHkpM4LyGr
5iS2qp59Ub+9SBunas1dplSfKhvahDrfGEzr98D1TomyQAePWa4Fya7IvFYw8rxKnilttUMcfb+O
JFvnRTGBdaYIxpf5KkQPvA09xNDSuBrHHYYUEHwZcbXOeXJrIKZlejdpnl8XZkMDGIRrI8rQX1P7
bf3Ff0sUW9eYmCyfnnb4Tto9bZCNL5yrFuvbHe9YV17itLR4MRNyXW214d43+LCeQyx1bvOR4u2u
ihUBKsw6XY553DEAaQDC+sVbzK0pJPR/2TsBuOEvGLOa1ZOybx/UIHWfOpFJcQkW2ix1O0d6SCIx
OREgMMG1hvxrjVaV+PjZYaC227xC8HBVqo9Hfegd3wu+AqZKTbzVIx/Mwd9bjYKvl7uP4wSIsKRo
o1SU+v6sq3L4lCfXGh4AP4yKd0Q7thLCa/LInCWoVyfT7TJfWdcdvERmyAg7OLARkRYQ6bspqKXW
6kAWi2Zr5Ze708BQWZKd6SziOODor42I48A+XVQmwgHWLqeRQc11GBLAdyi9QyyHeZ655D5Qk7O/
fG6g9IGS1rLZeKQHPk2RMmb3bF0LUl701UL/Ne3h4XUHO2hIwBF2WWpdrigPwtaTLEaJhCdO1df9
eioWzyB+u4S3YBOLu+kza5ByKDAn5Q2x0c72RVCjXtVoSEMl7bMb9xDaa0oehNCDv36wEgakY6LO
gHQ8pGJ8m39MW5QBCwieuB0ucZkYNGDhlQ3M5nAl+JfVzq1iUCOKYRCAFD5ptbZjASvHOjEwfC8v
21JOjD5jige55gwzfmIWNnTUjoVp+C16fjt9amMMQJLuyMk0lGLh3MzZY05b9UGWnpq3ah/L2kiK
1sKV42OXju3vBhpjpOHjf7apGAYKqUIC3p8axlhoOKpzTcj3hOptEOKl8P/LM9ukp/tA4kccUTN8
vEbZf04+rmlCo0MDQghSWwq+qyt2PgOafFA+Tg3zsP1Kd4f7OWO2IBMv6OOrd3G+eY1a33vFhoPD
jJ5RzqF/5hJY3R5vzVe50335rZDPQuooqsM+hv+h3qvkKBvfeHABaUMu3S3LgQ2+XUSI5VnD8OY9
WJ86YDBS+HWYR6DKHmkbMjgMlSJAy4hu9xOWEenapeS3fpdzClxfBKHCnN1TvnKH83W0jUrE98Rd
QAAliLrxT7MTCTKGvZ7ISUW9CW7KgT8SysmZIcWH556mWZVq+AjV2rfWCm46LumJH20Cz0RbKM4U
yASsw3F7xDyNBS+ukXA9bl0tvB4/5BqCZoCmQKrDgcQrZjDcR+kYwsz5u0zzasose2l/QkHNp5eX
KaSbeibIUSVTelv1kPLAUJbg2RCNTYfzAYJEX451VfNeYoJRUI5Vz8JSml+RxUMZJM5XRLoUO4cQ
5uQD0ohf9GNgY2UBuToypjU0AlnMNAYbrUk7zmufr27UMsIUvFAUh+ImVFGruloplavOwF37FUxG
d11S1dAEmpiW3njT63KspVGUYmf09PoYDdbecShtm8hY4WG/4BxcaSzGpmz2w6NfOKHsob8PJsXX
/KXj2+b/aChFBpAOUvM7GCJ309MeccFIfh+IKwNvW09ZFCHQS2QRXcCgxHwVgiD+wzdqqqivwBLM
PcfLkcDI7FHnnIxQ8ZNM20Lkwom6BiKHwaL/smG6agZ8nVzF6ZcAt67S0Uz7slFrSg4jTE8lzz4U
8DGVtWz5K9Hybc8j2Q1v0va+u1S5MeORSYDbDEY1sd9Et1AM1rLEOyGGbXXzDGaDnXi4XhhSFBl1
iUdNlhDOX+Li6YC49gPrd474QOPzouRg6E050WyL6UBA30B09tOmjFJKjr4wjgnLNDXi7Eg29/Wr
qsGphIEa6jRea/R20UJTKqe1Cw/j9k6DfE0cIX6ryJUT9Z/az6DqK8H2qjlZdkOVyxwo9wG3l8Vw
XyaInndVYgFWxlyBLASI+zQWJDs/iK9iOPSy66Ma+x+k5faYS6nG0Xi22+k+YaRFHrvqcugMu8ND
Qa4up3XM6PMiscPiWxKdd/XGsiNx/PQJDdZJqAXwgs9xVHknEYlnR5HdrCfSEoXiPcYWAHlz1LPR
1gM+eJLxt4LXYg6eGlD9uYMRWamYP4njyAq0VFd9fNbHOYdyjbDHUqdSU2C4AUtOi8lnYt31J6AP
W8qwuKSpmEh4B+At2S7JVtjTT+mTNvUSjKJB9iZ2OrgJXf/uSFxcVmKVitXc5u68h/F8lF6btjXR
RotBq2cdaTReFNt6u6DYHw0HLdwEtcHu8LbfPgrDVhcTXj4Hcb+zKp7f6FFevZiZkfk9Rz0Sm59n
92lADaLa0GyaRuT3QSYyYrTpJp1uKlPTRjCkL5s34jtxMRYdDfBozy0kdHjsxWNhQBoevU3prw2A
jFbViNh6NmVtUR0KVUK+B1BLM8ppHE/1GI7YWQeMTJu78ulMJSLv7np1kBT6sKc66tdrbuDhCLnS
m3Ye4H6RQHtJ9w3DVNuQrLkAo2AJr0o7jH/IGZnL6/+ZhpPweaMOWd22hf3/0GLmxDCeZLWsucnB
oTQfqN0UJzi6iP/konEZu7I+xe8b7vKtK81y3+WiLtQhLT7NtfVqOL0UuqbSn7VaOwqqqKDAemcG
53m4ZumrwWg8qnE45UtXS/R5hfS5lF/wwObt2xAmRtQyp/GuB7RZLGd5DQDFO9njj6862RKUHjpt
Qen3N99FDBWOMed99HkKZBJ6OH+Bxmhy7k3AlnoFSaitp/661Q1nLqSwFmu+b5FpMtnH/Pgqaqkl
QT5t1wBmDaUB6Lenre5c4ENrKz2rs8ykBvPvXjSzgbFDATByr89990LEvU6fVeHYX+GHgBM/fVWh
71iQTRuzwgyKOMEpDl1H+OlmdVkNGWltiVStRb3+P6B+Fb5gatse9ahyZfmgpidjNMoiw8KSeUS6
RMzDd3GqhQcHineEU4U1uX9lYvb7UkFqnyiUVFo5d5214GqPpfZPty6+gIdy6LuckFD7/2mM/S0S
K/G9Jgh3tnJrUdaBpSEH9y+R1+aLK0GgRftni8CxSgkSQTtiJhjWM7fNRi1lAZgtzL0fw9FozFcx
RekIbxd9DDqowG4MnGEA3DEdqYJKx1lU+bi/mESHnuYihNq0iUdNguh1Tq64kjdOd9QpU3Qjq9Yt
k4dgQ38jqK5SAhy0n9TwVxB7LwV9GK9153nlS6E+CYNbXZsOWshHzbixzY6LMDsq7C8JUP77ldfV
9RbGt36k2VWssiywF3s3PPVRVAU5sBlDdjS6hPIilEetA76Mjpn27y1THeIKraEbiYg/RE/vVhCM
z0OmFI/RYzkNtxkS5D0p8vRFuGkJjOc2wum+E+ced0BGnEnvDGu0uWMySYvKlNdyLoSMhcpo96pa
Rpdt0puDiLMuG8YLoMd4crMdrLp5+gvCSVe8DxZpD7ooZPnuFrhz8eUK59KpmaY4vsk1Nr/mDIBW
fYdsW3T6eVt7tVVciIixx7vKTuZI1COlqvg3UmwTALlxH+ZTb9XAjCskJrsK95rDvceHB3U9QhHN
Qfx+EtP25LXWP/5IJJ+YSqDgUmpwRFWoH8DTcXAldfI1bN81HUNEKChjVDvJmAmKt3smeanrVJ42
GDgR6NCxfSF4Fw6s7fD4PQtfJwpzPZQ+LTwqFOiLBKsPTlyVWhoOvH8XaalF0k4doHBdjqKq+UaK
cOpPv5pI11Q392Zgg/zsgueLA7BlHJyZJ9RZ97Aw2RjnApDOlfgLiU99u3WxnCDneLRhOBGLtE8m
zwV4fLeVRngjpGl/iYLB0eN5kIfuwgMZeDGuhQxF6WC0YDRFwF+ATdw4Ad1mhDN6oQbLpDBU5rae
l2KnchxzLkKhtcHet/zoZcjhyh3USiy7NxPPh3ZWRgFB8raW4JAc0ckZ+3LfEmuYc2Y7WxdvoC2b
hLbq5JiPzAHa3i/w3A80WT/p1VEws6Loklz2SR8Qcll3qmbTI/h4iLoRBKNPRNm8kEHI2hO7PwIN
vIQ1EOyOYBdIGA0/NczqI866MxMN1rkE0FeU0pob/RNFcGZWIs4cndcGcdvyA7ik3cktV7d2lSUb
NCsixJcAYEYDWpN+G1+GYfWfY9gho9K4Oq8fiKZOmdTZLXbQkWp3BNCMism5JqEWQ8D1z00qWfIT
QRleDUVfIqkvIhyqIJcq9Ln4F9vk81ayK/sePfsK6DDQJyQWWSFTQG+EpWTzpqpvxEDKdn/hmsSY
+/pm0wqUqATYXNFbwkcMpBnT9m28dcLRb5nulOgz7rEywrHqyKe18Gi9hsuxjXrF0Z5C9gV6Vigy
0+jspjNtoGlC4xZQjWaDbZtBz+EKw2jlAcr9Y9HrNBsVKupWPkumJGhTDk78mMRqeL1XxAsSSzsm
ndECeDv2rf3hDfQMVWy2OLJqHUtjK/wLlbuIa/yKhnsw5h5MojyFBYIg+ve5pP48olt6+Bt1WqOO
D/Ak0JDo/czDZmRUQqk2zzixWU6BrPVD1YiYsKAgrxBb6M9c/SFBNo0sykQ6lZZHcwnaxBGzRaKQ
13CMsu8QPfC14TLO8314yzLNcpZVuS5HPyKEJcTvCAuHrXmLezRXdytKpR3ul+33l4tdVxQ+Zyy2
YPKBbSQ74+kZ4FPq3s+ZX8WGQDiSL1W5VCtbgTHMoUuJyvq3VPRLW76dAlT/F4L6qKuPMdupid4w
8azXrTqAe3JIXO+OLcfrgigf6GiI72hMoFvQoQ4yLL8TzY3Hc/l7N0vdXhTX9+qxeI7wLEHAtLGp
ewJS1J1KSaXizGV7Yxyu2jsIKm+I3Ycb1FG2bZTjcLFmAZm7+XHbUt7EKBujeQ9uRERczVYrXv7P
OALcJVRv1kj0NRRow9wpWJCOlnopjZWtg8jnddHrcrATEnyLFXGFKT9Zk1CZVDkQYImYIC3yQh0M
Rx+WifElKQlgCBhOpDqvhnGUvkkRboS523gAOFoZAlBmhmpuOr6+PHQASjj2nUPfCDPuhXeBvQXe
07p1CkcfGl6MVeL5i568pGkeDnPh9LsrARYmeNCk6XuEz7ZDMm9pDO6IbuQYP1qXT0KUwds+rNsk
M8VzhzagIV/roywhmuY71vT2m5S59pP+FpsTWvTMJ53pbSdpCVZAf3weewTrU4w6GAqK37KtESaq
exTJl+rjncG2kkrYYG7em2dbK0sOyCdDS76XY7l3M2pPgbc+zLHbpiAufr18hJ8pL7zCoNhQutZ2
nDewgx23fZ3b4udHZ1PWolM/RAogk9a1pDKqQjegKtQ6cJAQCBQCnFLupPWNFvKYglRNFFkVVdHf
isW75eu5D+nhr1vgIqDTZPG/lur4aUU3mcWCo5U0W9ZHGZYj0AUSxhU8RVG+i+UsnkNzr7vozPSQ
QgDSO6rCYvNGtsB1z3ndLtCbvM/PAC1rLSzbOrAuvrF54OD/lYkUyfQfEXwgWlZs5Q7D9GJb8a8c
tsrPoSKBx6GzGKrxPsIu2ZbqUglG8e8owboBzQOt4KxQtgcfUHqyCEUS7qlXLbVX41PRjtLsI2X4
doGhMc8elm6SeMyivgNW0nlqyNsc8UIZK+NEFjYylvgYDjsLXYABk6p+EWwN+QKUckWElYtLlmBw
g5IQypksbapra/F8RvGd1OzauDKGC7PwaT23YnAUvgwelg8MVcPYh7u2sg1d9Tc4tHGKnjz0kYdG
7KKG2yUtBc8iMNZxKelkspl80lfauAoY7cq3Z+yQVpELdO7ydlYqOV7UgZwemrvlBgmNn4Uh/Lps
06maYszE3iV4kqARdGmyuQvx05DTm69RSrH15x/Y1F3GsQYnMktAvPuel/E/sDFQsyzpvXEVykKn
Kw7n8JalcG7uToiSfUNx0cG4mGlz0UfBKTuZMq5z5OPXdKW0+p4Wkm3ZqA6WCcIxXNKWwlDh5x70
+5qN3VgN3Nl9aL0kpMk4cpZHgGwYQMmZFvUUEodr+VBoRWGm9tvUoOp8aVs66dbWtz6XqZ8h+zCa
Ie78iE0QQFrbUDqQ5VwPTIKFVqIzU7vI8f2oFj8//Ge6I8Uq69KLwlWRWwNHqZPC0cNwgviNEca1
U5VY7vS/B8Alyjr6BCMG6YNgSr5fKf7MLotxRic8PQuXCZ3zvoQJzlCHOHxZF7Qy7HrlyxN7zOuA
bTqkeNu4+xvCzUwiSCl15F1quGOJCmV2b3dmEN5Mi0mlsoqBk4IDBR7nC0OcHDnzvxWdtcsO/cN+
dc+zhoAgA8d4MdTuQNlCqLJagSHv4WT7uCwqn7tQRgpCUVasnDlkpTMQ0rjpa7o25nNbYwYOudaD
/T91HFXe7BvZq8yUWe83gE/LDZW2S01hO/CdIcyJ8jQPm28gYdu28JRmElJ7mZ5aQlE4j8MKLHJA
85Hi188cryUQVYZDjczTcGFjiFd7u6zUshLXcVUMagarjquGT/sS+XePNDc65OtFYO2dedLdi/cR
0RWOtlPncC0Q5bOXCdpkEsBRZC/9fGXgGkb2rb6tlGQ5HRR2jYD3ykEBLyEkql4jdYrjTunYB2dF
kR6SvCwr+DWlQbfNT4XJrCi+lBcQfIxNBLJHDwzkLZdIhoDpTUY8woKSDJXM62LJxincauWBO5rv
qXi3lfXbObYUKktUI2AUZa6BaatdyqWlahDlC2ax8kmXonhHxiZz190//FJAKTqHgov+qnnXlmN1
hKNnyKYT9HDTld4EZp5JTS5626XCYn4YcoVJ4d+bRmXbGA6hJoTR3oc4eb55ROCaeBT8/rgPu1A7
x1bqfzJGT4pzCL2j7CYGpmfI72dzSCc+X752UUSFwNTs2I2MhSZ76YBR+ObybqiDF4jXuSiEdgMf
3tnn7iRNXNNupXhDWMZU+fbUR/eb/F1PzH5PXG1joLDH3TFotPUvWH64lSSRvgx0DZYXFF16ryUy
ODGtBYo0L4zolAQhviZSdFGU5pOf9Ke+5vcqc8ui7llDHKHp4eTzbTbxWynlguyU3j1xAEY4TaAe
7oE61AdEA/+NYJpo1GU3dGYeheBDMJFNzHCqETrSTgpQ6v8jvroIWHZHwt7lFGjfhAlrkJ8MJ0RR
md4G9xcu6c5l/X+Y/bwWwIcNtJNJGNI0wiZPR+JgFdzG9ERE3CyIBxRpKTEUy1L687gM9H6Ir6sf
izURs32FIPLXv+AQt8t2Sn9jTKtk4pYWfNGnQE2v/+dVkrTMOSzGWNZNR0HoggelbOIlV4XdEp8l
7dgDxhThqqOpU0STJ5aOlDGDbdPbP040Eo5KIMQ7NY72ikXkFPChVqQDqT4nLLtEq03I5pyP/tqH
gA/0XhkKSwbGEfnc5gUexVUwyFelZlqpb3VN/xUxh+1VQJ6JcU883qdqCs1WOD+V3Vi0NHMHG8Vh
G/gPkmXJoPptGHS7Z5b/RbInPVjCwCrp2FUHJvBC4EXloFVymp5To/3S7YmNdfLCZMmxwHfNgmNS
IDV7uba0QU5iOIKC404DhYIQp3Tr/v7VGG3QAfKCvUmECZWtYUSaxQli1Dy9aZkFnbMkMlAhvJvW
H/qXDamOZFSwYjmTzWRoC62AXhvat8ufNVwYDSq2WmZxACwWnf/j4aQYZQFCYoMCXCyctnXGsfQz
h1SC7g8GW3XHF3kvMIMv2gFxrpM3rwKUblj4hHsUIAVZ3cqj9V8wVRZ/F59tg4trfu69Jd7zk4NK
CMIv8H2WqygUdZ4tKwUY6Zq7t2tP0wydyg3kU7gTSAiJlKxlgYmyheRQlslzvvlJhBITAuKY25Qo
AzQPMOdAdq/lmQoFJq6LQAelF0u8XPff8RWxew/Htvc6+gHumCBdx+E+jN1Uws5W7WrnDUFH+NtN
pcJdXFB/nzSwQk2Af7HsxtntzyTM0jp9PYNGRG8uzeIuac2HoAw/AHWHf5yzum3OAkN3ZQZi7Fq7
FpGSsFPUYwi0h01c5s3/3bpeHacFIM6f6byjcANp+034RbkW3mdjZi2d8EnzznhxELXqXABH1sM2
K5BGHOO7vV2wpoi8j4qrUC5FSNC2pn7q5vP5vBeXvIFYJSMmoFiHMH65R3bwmriZWMu+ryXftUiC
rtKkQ4mPQHXU5mweTfo9W3J0UCnLPINTXGiDIV9szdaTden1t//vKIieuXZGsMor2UnTacRv4Ld5
1GXs/RWdBfW6uKgdhfALy1ZQO6NCCB0M2I2pGyqOExuivJLAYCRHbtB617B3gysEefzSfvXPW7e6
V9Z6kc5PTEJMz4To4bcmciMvYI6gthi8OLSUmfgg/lZYPCznx9+zKxwheUrdNNSRUo27sqYt+mqe
y5CanMJwwWZx+SWlkT9FMVbnkcHxUmJOWZQrcTdF0DKL/1qLHCUSdD+6Qcsvp5fS8axGjZX+14l4
M83y0sED3QArI4HOITRVG+xgVNNrJ/DF3MWLDKpjZeH1ziqTS+LfLQ5hAjFR9c0Kse2oDIEdQsJ/
f7w5myuzK2fDGodUnEYMacFDoZrqstQfEousblYl/gfF+vSp9LXv1NccBlWjVxx/P/yT5U0a5DQt
lsbF/OIIqMIKSsoDoIbiMxf96rbVlXNXDzqyC9DLD4XnZ0PhIOvwkDwh7f+f/mVU14+Fg+MKMX3V
+Q5qTeKGBG1NJhbXbO6jxsXO/r9jNamzwq6MZwhY0qj1RBY9O9sbz/30F3Ftz72XujI1nYtlChl4
edSgW2wOhThOWWMl7vMQi9LzvwNv3PlYY5++hK83Iw33fs8F2sBnL4a94uucPr2FJtIAlQhShIPq
oh1ysX1OMTT/P7UbdzmZDmAj/UT+TKpYPEScU95+M/CJaixe5C5xdi5ZFMiN9bnqcNjiMwy4PyEM
fEbJSJsem4idcJU8wcTIXuDtwQUX/T/ggiOgZU5lHnT3mxDh7p2IXzc6kjaKzuw4tAWzNT7A3EkC
HgGim/ca8Pu8RsfcVjCmaHWq3iSl83VWktYeY7QjTb2/y/LJnf7mWZ5ZUf4v+dZSsLYjRjutDGdd
4kE3W45s2oPIUB3WJUy/adLal9FwBRPTNNXE8A2Fwns9a3klAqs8QmO5HmvLB0mIOzfjd0tQ3Omn
bvK/vrt5ZKgFVGZ8iHeISvve+wSLzOB756jWgPNu+NuNPwTEcKuvh7XrwNlhezz6PmmKWjmRRDOS
cHxaZ3Mx6VO9kKNxaCdTI+1jiqjvF4pu7LFKgi06PZfbwemzGM94eAiRGaDlMoZyIsi7zRf9AqHz
qNePQfDaiTf+s72KyDgD53tBa8utXj3XHCE6eGdUCChevDA91Uy2QB4d1Qco/OaVlU0631ux7JJu
uonj62szU2mLaQVDveyoClA7DrAX+pN6mFZWkyRMiYm7NTXL1b3IhT42Ol30o6SWdPS8KlPURRj7
NF/ICZnMnOpq5A/lezsyN3VRyavkANzWEl4Lm7JyQBQu4OePa5x455PxZ61LwEb0J7u1enm/cn3G
u6LBC/1owu9sBDUBjGjWC5c9geWgsUXMYUyWiGEshxfpp3khqAKtcnw1+PDqiQohK5Ion1BIRXDk
BFsV6aW5O1qT7uXGYOSU6yQu1QrBVHAfvBqHzrBAvnfMGfRiYoZE/27ChLKdaqP64FrvFXOYwslp
udLqOTGhga7FdAYZGv8uk0m9SgR8VVZPP/OA1GoLNGNyM60iqxy5izSfcUL9P2gKKxvT6/VmFtZO
e70nbVO3Y/gR41mgPJbZVm0yOFQKVR+1wh/KG1Ib/FdggGNR/la+kYw5mVw14xeBZ3mShmtZMtDz
LxZOd1jbU5V0lnqUCQuVrva77p0aDK4HaetS5VxfM4DTBqsJOLEDF6HB3PtofB/u9vk41bm/24AQ
3z1sJ56ZUCaagEPWnn/oXrJ7UVma+UpX33VSpCpWRhNV59a5tGfMgGAEgrnpaHuS6UVWw/L7iPfX
/blmVUKZHoEFGgIyL7top+rKRngnN4GtqHUwKZd4z68ZWfWATMZuPvkTkVDrjB6yIrudIm1mjwIL
o5yw6fM0UIrJ2l8TCGNYroClfih6uBIijpwcW6FAjktGlQlhK3AE3wEumCv9kf1sBaVaiYVaGxiR
cwZnXEb8DzaF7Sw4LgNE/VFH2Y4etckYny0pFvijZryPZFUkidGYXDwTnUBRJYN2FfqMQi9dhem1
G2rQh4BvxYMzKPa4IuxRUyHVUgh6MafaLNI44ug8nZHH2SN3a8zlNASfPoXIzs6e4Y10lV+AmRtM
jT36r+CJk8cfMHbRFTl9/lPvZL4M+ds2wLH7/X42iSrjEQdyXsL7Eg3prV8uABdt1caEDCDUFCbu
yHRqH6CBI/TWWQJAqQcwIZPfwNSdFfzicuKvsT04wVswyboZq4oc4Qh+uIY84b/Tv9ovrsLO45aD
pVfZcxBSlIAxhdm7u+hgZaDaJyj1AmFHBk3ZtuZ1xj7+CalB6W2UY+uZ7rLWGD2gLKqnOcTZShhu
6gs2PmZnthx7L1WMvu4WM2LBjvBrqUZsoFf+WTEsWsLzqF4tru+U02Mbdb6voX/9LB2/PtXgvLRB
jZvC52uVzuyPIZfR+ay8hiARTUD/dUl+u68iW8XnCwvtWxbrOAbhyqBsr8D6leWiJebDh78RBp5/
HIHrHYROIDiHYEmh8eZ3tghiWU88zzUpDolBzgdBS0qduxUyos/rzZWV91jK4L2SgiI5sKRKEqVr
Gtgf1c0pLX9fzEieDKRIPRgcL7cHT0xuKPUT9Jf4a52iX32Z1+KamJdAf9/DWTWYPaf16i3P55IG
EvJc9OFM4tSjHGq23w26BFdfCEVPXqVJsovMNfNHqK+wHbfYhZLAuEwZFCDrsiYSOGxMIxgG5CUQ
grsUYR5QMFWnEoc4AFwbvIwL/oC7mQkNU5n2OU2IqjuqSYan90LytLIHL5aTRq8v/1tmlWDP/WvR
Z3dLtxcTiFhrIZoxaSpxksbg01gbd9e0ci8CQJJCX/x/4Z4xIsvYH7HwkltoAm0cDf94SbtLdTji
JsrxcRzL/lZNb8y9SlwS1xnTh49OIng2tkELqVP3zdy56ldwNISwx1KRYI7TkuKESThe1qBnRq2S
XoyXUAd7YwnD9pQbQ4FJ8Vje+m4HqSsxL/HyG5qrU/CMHudvRskSr4hA3+sLTB6SFlK9Pm5EGlmb
NqAtFgTn2iVGQLU4G7N5/aMF7PwMl4h+GtoW8xPW0TUPvvLlWsQRsCmF74DP9XoXlhk9rF7uV185
rOcwdGB7GfB8P22jMDkoxvMr6XYohowHHoxy/hVeHx7407jQRblc0hk612D9FvnEKHz9e1zOIjvq
WFV970r9OZgnW9PaXMEs71xoeqfO782DeATfQlU1QvKA+Nh5Ew4Y7VefRPV8/MsuggTnOsIXOOpC
wzGNivv9Vs0KmmM+a7Jv1iTm+aEzGJr7rjyVo/yHsSni/7rENXMmgTJZfW146oH1d90WOXwltgzY
4A2+o+26r2g/4099T2VdN1UvEx5hoOvUNxPL7YeM/o2ADi51jDF3juplreq9XTcTGtwfMfFKidKJ
K9en/dwTceBxZsuADsDveZlwcJHwQjHwYCojRlAFgK+FMlk4aA1/cPzgGdLObiwDmoeQ5Pb1/v0B
sO6DjnxV4jl5q0eEJl+pWjYHSFYnG6bOm/GuiGYO5u7Iu5AHfk2rktmMaNautoH5lOl2r6BaRsm9
e9OHMqi8hMBNT1/GXh/tYRkHol+ac9eT17qFoW08LfsR0D2dZe9ZlKwbewE5P4F3cjI4czgO2+Gq
z3aLQOZo5NBxcr2gKZaXDF8wTfGhaJnD9Iaa0gUpctSpnvUmgUUd9yvj4eE8z+QQ1/4PJdjTo7aC
hr6GV5LGguo1fNgBmWG/3cdfq4OcnXUqBm5d7nI9kT/PQNKc+JhYtTAZSq+1RgWmr+s8ho4oZvEU
2biov+3PT4LsNguuK758LbskmYOnaKGnuhioAFKdQQIHRoJ4mys7J3pFaBj3pAI/co9kDy18o1vC
D+t3RNdQsmCBF5MkKMELv0MT4Im38eAOYw4rXzbE3evrINkzCv9zuSaoI3xiG8kjEWhHaQ3PkjP5
w/jVT0yfyEnF9VlLOtm0Sqd/aqByLh+QnuocoQf6ri+KJ4mXaLGB4f8gwBVV4NanstX5nS5xAqfA
cVIFEaRJq5hyRjQNQLNvgTtpopACJD62q3hGHh14w7MvlmIGfAmfuLdd1v9+h+y4rJKVEF0ZVxyM
xzifMbmAmLTLJGzW3ix/rAz6x0go4qCvkfQw9WhwnIJfxdqYPeWYd3QBYLIirJJVwRZ1SFbWNXBE
iqXqVxppa+0huDB7IbAipO1rGHXhFhmO+Xhn2Rg1WE97kuPz+0EiuYYL0TwIxkiqbDJLT8qQ4mU7
bCGv7eOYswrs3Sm6VWiTS8PD8TzTpR9fKa6SCreUrMx/3Ic+QLQtCfiLm6kczsZq0/BITU+bBMOu
LzzSnckmDSyOYGFFOYh+u5uWrIsgcR+VauDDLu82YfgephbtJ6kJ6QTEeTMyBlEewmn6r/M5rDKM
FdIpfugxwdtqea2884KyBzwQtKyPDxYgvjgFyJ/WM2fKNXIixKMLgC6WJ778km8CGVd9Gk72upNU
/Lu4qKScPSHeSq5uVr4N5dwnNpjo1U3lJmBkYmzlMoQgm2PiCZNAROqLBfJIRyaVOrTykqSsM9bB
wKYA+SdUNnkYSdzIzv2h3DGo5lfux0dOdR5kQjNWzIMrIU+ia0Cxk1wO/XYEH+rVj+RGrsgVU8ck
/6uroRHKjkL9d4+IwLc5GGzN2MQ3fIIH/NYuoKrEnxbA/67orCpvmInCOxZ+1owx8x9jY9Qx1L+6
fJu6/zOV43ByJCQ3/n5gYNrrn+5oI1ZiAcmcylPU3d+uhgWdcSyv80afo1ElB2czRyLgOwQYDGnV
CpdJVtwrNd19zntBHJPcDKn6IWx5ueHn/fJOrBkx0osol1cgPfQmMzYf8qRa8dSoKccY9h5J/FYm
/6n+ISWuJTU6Eko2Gsi6rKRyPUvgjgbTmD4my46KVz+rlEBFZ9tq/IskbnbFvr+ifGlm1N7bMibK
JzW7DmerWnoNINHNaQ6GRQsACDB/gaWvw9eAoo2M93RJyRysMzPNiDfXJtTznGpt5Ho/xfBPvc10
f4T/4/ZFJjDfJ83lm1NXCvyz0lWIZutyqjCkRKdUxnniN+IjydoG9rIgETk/N4r/cGFk+Z1iNCVP
u5O+bc0c6fDDCRmP2GoKadX/q6sL5boVCIgJusJvtfNEr1IB2vzL3/FmZnr8K/TVOrwoZKcXJIEh
JHqPOqPvYRtvYpVcMxrmPpRYnRjUDaZI0Hf+O9kiYRENQhveyzOVjB8Iygx+aVfAyeWWyFVO95/o
Pyn4Z2OC7DRuTIP3N8G4p17o+Ngc9wQsR42NDfydEczZiQNuFD5KdCj+Ele1bGSqW17sfmflmupN
d3XAHHtfvVpY0ujg1EcNFSAEv6ZcFr4DGxrWjIt3jACnwsD76byO9j9A9haxR6GSrMT6E2cBLgU/
Yd5U6/T8uvfCD984Ou6JhxXv+xUe89Km9VIOZHrPTI2x9VGh2FXpAUi+awbeuepMhgLF1+7g2ClI
jD7js8XkoD0Za9106dSiacbE0Nwe1eK3xwjsnw6uRe2XTHR3D2HF8nMSMqMaaQN5+ldOoDTbyqK8
3MfIugagpiCE8BHSjM4dSh7oABnlvE0ZXS/fTNr9SZOkKH84mpJ0xzj/AzOw3KO0BThuHlJ87fg/
UitdrS94sVgGnsFdPB1gezNyl2Qz6GYLptf6ijVHD9yYs5MTkZjhj9d1b5NJO//Jcp8foPjRny+k
itWfN88ib4Ahlf5d3NKtwxBfxInIKEes6SMyeRyUPf27tKu9sr4bjC9m67UX3KBQrmljDUqaqFjr
WwSAfbW2dkk29pWV3HzklphxR1+HUMUznFf0c0iGsaQ2zwsqaGzQojfOIZFsZHlD61YFxZtmBtkh
RG2fzTe8eha317heDEoQCKcsYMOUhPcFf5h0obb9DRYiPyzjbjWnpCA5ZIZLbh26L9xH/LIE0XRQ
E73RVjEjHa/fbeaYBonhXB585gMvoclSII9SLOsKxxL4IOpk6SLywRK5qNL0E6eWLSI9FN2o1YmH
LlK1AFiIyHF54CDpMM7WNMCE2T5Z01Uwk3f5lM36KjMn0ZN81Txbme9+K1ovfC4QjifwBMouWkLd
20eKKe5yLRbwv2ToQW/UwKt5J4c5Yg+KimX/7iU79yXGql/2lE3thu11xPg2gYG8XZEP1iUMYK/c
1LhG7IseT9xhafef3N1PRK3Uw+a8yxcT7t+n2uRMrDC+KHhI4GhmLl98qCyaV9zmcihAZTNvR36p
7NLTxYT9jT61qKLA98lvrR1clv55rvkBihAA5Xm8DGPidx4n+9PtQjZtNdjuFZ1QPi0FkbUCZXF7
wG7VkKVSxWCkvWs+f8Ycf0ksZHbpIjD7BaYSVoSj/Wi4qBPIVFyglLEZsbT+v3uDuJAIZaBn3U4w
j4i4yBzNRRUUJKwe4OmAs28qK66fH1amYucps0Y1yDelJnAdpqFIZz3P1HqVr9LI5qO5bT8Ct84r
nBuQEzMK1keYMcsa13/OfC+Di1y6/XYGHlQjakC9yisVTICq1cUGcvRFRIAxXbswSuygztuPJljS
uXErgdus+YWfj2po9Kp4ugpwm2FR1NkfoAQSXxgIQl3SposH/sxvyV3SfAB0wsNQMxfqvqEenKK4
9FBpvVcvcHN4fjftyamF3k1375K7EO6nlEZ0/a7ZLSETLwQBJ5TNyZ6uT1aO8XsLyZYPP/j4/F24
TWHcMArDQQBoB+9LU/f88RcE3+FyBxGbYBsWBVUgAC59lQ7DfxDPwlFD0fQotI2GRGolFeUGgWn2
djWfbKRPcRSHQZ2Xvajq/XeYOEtX44uklzzHXr/OwsF38ARypdf+Xg5w8kDbwT5hOFaTJQfrAnQp
L8RlA9Gqb1T1pWDRVbVtZJGNTYQDT3WSp30wIoBTnlm/oqL4U4VMD7YGzi4NZPCXBfrheBDJSrFI
LYtg257HzJUL2XenO+wMVVunABcjGBg3URPp5uNXFxTCDLO60rkvM0zt95Z5ATaArIJJdf/9m+0y
2reXF5GiDdx0ve2aJ/UHNrg+L2KKloiKHOXaES/qE6x2FiiKdfiFyEIJZ1qpusJmXVMZdkFAvCAi
DWaAFkBMdB6AXrgiQXyFkkSS8tzbBlq+FOh0ripCC/8CkQCqsIKU8n3EJ6y0m/ZPN1ryaPRnzW/0
JCfP1OumKIagexowhKUHGu2zAV1ICivETRdxcOOxJqui2Dbw/1homxRxcvWpiDRy6XZBOLBZofgs
VYMz4wCeQhKqGMKSn+18dsMqS5X6RwBiZi9Cz8yybtKWkgdZRAK+KnGlacgs0Dtrl6S+OsUpLWYY
5j79tqHwWhSJy8YAC1BQ13ZCz1D3US9nM8NMWzJHW2XHDrEleIYshG5gXrE/6CX9HxvV+EViWl7Z
5AJj0NUVlLpShrMbHUiw7MCUqS2euROyrMwZVW8ol9QkEwvK5AeY/SZ2ISpi/ANPDE6kl9fmiO+t
d6+cdEVMyaXxEJXkulHGsypOiA8DljEqb57Pk+lGun0E9E3dtlecjB6zVb14daHCUAmpcaqysR1l
opRfSWuGkMRBhpOl7PEtF6lTm/Op8E1DEjNU89UHgz0pBmHP+3LFdpxnnaf+NoU8GXNHPTHJUMkr
ZCE03UMfNaQ8lct768yXcC9wTdFDZ+LmvS8NrsvwXiQ6dWvAZ/ZrWFtiU+lpRvmBIubGLyzAugXl
THk+iEjWuwv7sXDZUhpd0rooJoIM2/oUxWrS3x0xJU4TDTuymXGnIGxn/H8Hg4GXXj/74lBYytAV
ag2L/5ea6/199gRxrTgwsQn8vnwJU/5AQ77AEQ1NYondRZ8/I2anFxykwCvQS+nCL0OKytHZtR6X
imIyA0BJPvOG5QwmoomZV58KKZ7bq3LBRU25y7LCuEALlcFIYMj5YqBJtBHVUblAexddc1Nsqexc
bOoZdxu1TIrtA26SCoShdXQ1t1MVgNRT91myK/WjHXxy0PfDWsk1pg3aHWYjh+qYtXUhxc/DYO5B
R+gmfKQPRaje2OVgyFVuY8QTa2bgaCUN0QycxJBrhMY868OrgGz7Y0o0nXd7c0Jc3/H4bNMvs5vU
Pnw8ZUvs4vHfG9wf6y0tsRMJsaM4Tyh7gBePExXPX9OgCaj76A0aSXojjx4bbkQY1VCQBpcy1wHQ
MEVeu6a4TIYIznajrqOi3A+ulBSS/83+OBFqT7q/9ykQ1kHrQ9+tyDSUOaKQr2QCZvsbUfXTG59A
oyJW7YQZvGjMii5rO5IxlIeyCNucmYTSUIkFajXPIiI7KlxxZEkSYnQRYVk7yeHAHQPO1eBMwnrd
vCxl/sDAgxg6ndC5LuAAdGQJY38rwnrgsRLuAuXwGT/GtdriION3McI4Ipj1iATQmQZgkyBcZSU/
6FnuUbDwbzrrEMCts2nuPxcayGn3C52t0JmnCSKEurUdJdBpHdZqMYgvIBUOmqqhVACycT/xGADz
t6UwEVQJzxMF8DDZd2ywci+1q2kexyOrONwXKYYG1G2nfXw34GhlmdvpC9iUFEdqtYOiC83BrJVz
arCsFvrGwrCjTZ79+TW4pbOT6ttvVTkGXDH9rRaoFnEakIABfNYLhbvXXi3zMgmk9j6JJGHg5LvC
jkXglQjKXq0D/4CmOA6FnOU0Qg0lGCdg6q+2yuWvJKI/iI+lD2+HIj1DNXsMDocoTm9Qso/2UdFZ
z1OYz7yELaWuTm1lRkgn3ZNxcJ9jGzI8+30ZnzFKXTJ5oIwI64acxAFYkCASxIKOAh+G2AtkEC0Z
um4tCcOKnEIs7kyDiFQn+UQBQ57Z0W0trHEK8tbKhCq3mPMLd5TxzzVLa9n8IkqnNbCfD9nv7GXf
MSorlLAx7io+Mp6NIy28DRgiYV+XabvemWFsDnbfMAz4sRH5c3SlcE+yFCCbfJOKq13gsvzmlUgX
rGbJ03pCAIZV+uM2kp9BCZk3Y8tA1/TTwFYK6sKLmCtR5HpqAZ3WhGqwumckmHtZNqAUxNBdXKaH
AKU12DJ1fDPqflyLJTFeYuN5G6uqYuYzgXVYZcddZHiPN2mK5svS6/nPYTGqUo7oS0kIhcH4hINi
SZoU1//Q4cNOtQsHzgq7o+gWwINubXu7MHkiIZtDuz+uTrP5xVFiFuf5H0rajShySEkEPoeqQ4F6
qsLI8QKjJvmwAzO5qU/je4eEks/XOyuTYmiffSXLR/8u+3LqwkQGKDtPcbrqfuEyaGHgrfIu8zS6
8wnIaF6JGaMh4R3+o2YNePCKYMDLywI+qDI6UVrcKhFbAaalhRokQb26ObKNoDtXYl8BvNnT5TwL
RbpJNFpju1S6oxYXj9oeMPKPenXqEtbnxDiIU+g10kjMcmNkPvz2iqObqfL7eJG8+Tyg9Umo7Qo5
3rTLgvrw9n11S9SxLAOM769s6TUaZsNRbiGBvLS3Spd48nGlsIwss+kxdOC8cd+GNl5MjNfQy3YN
pwmMHtdnGJsUDAIVZn933xF3P83PFZDc0wHZKQELlCYZjB+jLlRNlOoAh5JJNbsWTy0hSUhXW4Mt
zlnI1K7Drh1hJaCb0bM7hgP09bxK72wYpyJU0RxSV5QVIeWwNGajIHspog0qTffc5ZQN5hg/V5q0
XsW6tO2QTPRTAVSsaEFdZjmllfxjBIIBRHo1yyGa7CiBdaZLTZaV22+U/l1N0UgUHruUr/QwSerz
oVp9ISRaj74sRBVP/w25tCndr/zSoWxYWGzDmjRFlPmfOtjHKaADih1HpfFkzR/hfJkHjiwosIiN
tKE4Gucd5imUX7HV/hE+LySsrw2Ob1p8DwdivY7xzCA/VoBzYHdICgKIBoE66BDsWWZ97FsT03B5
OIW0WPKNFjZ7A12RRZ+lGmkEqmBfhDM7ldK/tToZ2WM3LsPB+AQo4l+QMfjNQnt2VeY55lth2t7V
Sw448rAgFJ3pgQb+pYP2U4rPmgSX0OalJRwyepkcE3zFLZHiqoHLi/8oxyb2M/7RdKJ6QuzRz3Kv
7SptZOEQ97a8aq/tlpyXif5MU2h9UvndmAeVkbcrzYUdQ0gl0BMtVE7ImrOO4UNqd8rVGwF/Vqcg
Jsxpfp4yQyNy74HONHi5uy7AetgOJqocgB4NLGTeoCMxc1P1KMxCQmoNKYfUQGx51H5NCqLmFGgm
YyQvoCc2xNP4BbDn9Z5F8wy2gzte2uwr3eKa4GI9+iD1lmfsGIUrX0q4b2Pz9Wp7go1k/nDW0qDX
xxTC4xIoiYAz/cX8IPHppmkJ3waj7mMidFlhL6cmK0AOIDfOFaVodcG9YA2iqYPkZNUDrkdvW7Ar
2pcY3RZDGFcFFzy04yWzMLhP/JEkdYI5gVZi9mC1uBaLmi2GBn0jeJYVrsAB4LkdMCVqjOHzjaw5
GKcpoNG23L87imS3Mk//G6mmI5KwMtjQPvO1VWgfyWEkWy5qBLXVK93q1EQ+0HAT30SEOyV1LQJe
QnU6r2kmimC+sh3FiP1yVH7pPml8ws59Yn/tjbm74G3tq/7+j+X4wmUr0UH8rGCY4dPQ9FAGrqzS
dBvOAVQjZXCSThNN7nl9I6/u4WNltP1oXKfhtB7v/o6pYMXfbUTbqvHe0bIpdRMh86qqq+0eQCZg
fKM4mqcJSzI+VYzOJxjkQ7CePKp1aKjBhC+n4O1PDlz+LfKz21InUIvCCzdlzSPU/n44kfnb1tT7
Ye1Qz+hZvHS9pFdM52WCfaJJB1lSlj8q4HVXf/UnYhxKEzO/Hi9hGFQn6vJI6jOGkhCd/Amz1KbS
wRZlB7CuY3SXXesVi//2FMoUF1esKC/6LoWcT8TAOZ2qubYV2vYGzMlWaT3Sq/ZDg6NXkPW1cb0C
4pd6J4iG788pyQsOpf+2mlZ/reDdEkqmAt3izsS7yit1URI4SOhXSDm2pd6/CuOv5mLnYf1hrNGO
MaJ54kntb9T1tRJ6MbJMEa502+b0EjRT7EidJ3ipBZq4q2Ah4dfW+pE2xKn0GB7droMaA1V0qCmN
PPx1xoHD1uU3puFHaQdMDxYrKuUIxGDH/LWKBzDjpDly6tKMZkLL1ajfFuGBbFX6fzQit600RXEM
YNFcxJCyQ2Iv71Dme8P0W7S6EHEWzBfw+apx6eD+Hsk7Nj7r47PzA6UStciUL3EISQd3DhDvTNgP
uVZ4xDDSVC6rGDSsTwKVn/etViUrkEXTbJ4fvpJ9TNKORS/frBywaYTTavZMLpBuoej5mRSU0f4o
Yp8SsR0uSN5J4+Istgf6T2jLiDvbDtWDIEq06V8r2RKdwec8ZuKUh1AzrtaSHlw7XocUD+Fntxki
Yp7fdNKBLweoV/OBN1ZENI/lSYxCT/CQ+DLbsffqmzkL8npnV1sspeUWa732oQ3reN7PH2rabK0l
1b07oz0K7Lb0U5IG7AcIz2NzH1HkVA9NoMl6NWF2yf1yDQ16WHBqKwPEa9qKPvsep6xZ/5oV1Rh0
FvZ26gfhKZZk9A2ssz8719uo6h5/hZx5m8X200dCHezFfiJc188phkC4VksKYNxKUTKuXmKcf86X
iDemsi5fXDHYWQ3R4h+PkEHWveQcR5opEFlslBocBEnOa4YzNb/sDgH2WJZMeJsynYS7IYX0XVQx
QnJY4gKBipFSdPhZ2vdVRBV1EhY8tkwG2LH8W+vfxr4wR8LMYnOyNjsQJ+jioHkLMyTQ31LE4NLB
J5xByi4zNOiEGaZPF+W+pxBttaCbJS9gFoCnNFScMV0vppybkkgta4cCBjb/1ok/OCfL5MDdjMZY
jlUicOaEcvl9SwN7AUbAw1xEAlyASvyP6x3HwKPCE0a19S1jwPo6XrJ1arAHqeFET1dajMIWlNpX
tnWJpiVFAsHKrICpMxZBZp4fhnHW6ynRPpRe09L0VpCYj61rsjRP7fu5RkWKxfSc8h6TeKWyjdAV
szcPLRfBikIlXiUhDq/KHDIGcSiOJeSE3tQaXl/mmVqS3kHeLiOFdMoa1DdNjgeQowPIJyhTVVQ6
UNMAeLmpGsGR5/pCR/8CIU1PXPhP6zNDO4E6XFqaoBIrSIgUZ8IyngNThy5+2fMzsEZ4VY9h1b/M
u2ttQz2bCwi9A6MvqoZVjZNNVFzNsu4RqdBjFvzHfXqQWGEHc0HYotfsmecFw3UDEvFfmVtN8zsG
UEyvqBjc2VqVN2hC9YHiusfTDzvMKWb0DSq+pmKeeOc5giaxhROevMOeltgURCjQRa6XyDB7kSoK
CNNxU31/Q6f9VTpTj7EzLab95JaOLk9Oi8szLKbLv85fTQXCmhudoLaRLWybapwChssxOVOmA0as
PsZI+pXlBueg6N24AxaNML35e2YqUsgMTG7Pm2wvYDGSIRuoP5yb76ru8/uMIA4K3PTIltYmwW+s
wedvhRyLQs00zwWw+2Lmq80+N5G4P2IEOrjbRBO4GbQwjdLx0wkkaRZv/ALJsyVi094K//Pa5qBm
riAjpiuG/Xsh00PIChyLbqM5aQCkzgzpxTcGET3qHYELFyrhORNf8SIQPVzBjPY8cuDvt8n98NEL
7H/IrXneV8W7upNL5Q8B5FNNaB1sLOPOgE1k+XeXJl+GFmYy8zkvWkS0lCR9jlqKzB9gLUzMyaRa
0eaqshZeXC73a6Qnr7gBHte6YObl0HZ4a9sPjMjXkIk1cINe5gRiRIyIpj4caOmYF+4XlZow5jqD
0AaXnfTr+q+99oUv7ZaPoZ1c55BmVNj7/nUBu38Yh4Rkk/Yy6GyTJZtnjS18RUfKVnPub8+HlJ6B
4/TNn9qGQis2O+38VVrpFrofVnNuPChKGLu81UD5lCVMIDG9X10z+J2t+nGrA1XXph45lyUaLHhZ
Kj3ONQv15PCCyNZJ4UoCMPcaz1sNZKNSAY07u4P+mUYwDBBbYyRy6NioP9prHg96cQF4bKjKaLcB
CziXAkIQYk7PoST7ecm3yX3uIq1L9KESJVN//VX/UYO8J9AMNWpDgIEOplwx3iSkQTBaXh4yCBkZ
NeBn+kOL6ovjd4cB63Sr143nnC0vT2Z2ewVuBEYye5A2u/elHTsza3OUxByzeJZwfuRicjFYixPs
tQgALJxYDqP124H3ZqHqqzvmtd7knnPUWenBDxY+UZIJFduE1shb4WtJQUwX5d+lcruM50Vetf2T
K5sXa8DE58lRcUIuAkmBef426hAs560mjudunfLaqa1tNNgJjCL9LPlKKeJaaHB+zS+Y5xharRYP
zR/CvwqkqdKnXBRHnbV502mYe4JLeFz40P7yUWh0+wTGWDjKGPO6hMh18BSAAB1vXA02GNHKz8G+
8s9HOVIC+y8/+0FO29vfvg7Hz1ZSHRqhgYjHvtxr11TDTMU8l4EQrZA8rdBflcr5zglKoZJKktTz
cXDU4FHGLGapysqJpKu5uMaKeHtIIUcW//sj6/uov3XKLW2GofUhjb+zN971LGi6aC/5hPQIXNAK
EYhBVN8Y1mYy6vI4WO757g+9I+H30OMb4slIrGBBFmEOBc+ZdhHIc/tGghEwC/Em5c1PD2Jez6xk
dPCuP5KOEXV03D1o7LvxxsX2iSCV+bJtQRiccYEoDzryU1VxlzpiyztoX7RebmFfleyZBoUSJfmA
OwfsoufVIZlPuFiN09fGLQIdG9pWvU/yAw2gAb0wYHZM3qFqBWJDsE3nX5NXFqr5woKLMlxAVADx
t2g9VCthsDb9sNifLISHOPrdKTyO64IL1rrbRFTeVtQZEvoqh24Zyo1ca8ZQqWCy5MJKmMYF3DON
rXRDIXEPd3XLNOd9HsqsShuJhraZrr/YHcUTHc3MvrGkKinsqU0lUa9gG3WNIULjFvmeBCqXiXoz
ADtkNvO5/FXSpWLCQgqQy0rzd2acIImSKOrGth/glnOldrZOUZNbUxSgDC3kQiBIWHAuyxdnvjus
nJX928SERbvy2BHjT+fbNr7mXJHLYTpWnQwM5K0tdpjXCwgu7HeFpLWQiVL/gF/RnHi7/MqmbIww
HCKcUy7E1Bgrap6o11mSaHvpHVy4BJssGueWFsH8RbjlJ5nzx3mY64wYLOzr5xscNpGdt0kzgVrm
4TD21jDXOv6d0RQ4u/rPE57DeQ4UZtNyMJTP5trxwOXZCRB9/OkxmVgXkYsAGpXH+T9yvLyI9BQE
dbCO3dp8n2Gz6NHQHJcJGNvhjcj8vZo47EVoVDbe+KNFuSGJC8WE44/FXZCPA8euBcBG9uvS8cCC
RJ/2fc+I1wkUl0G4H55SmldsggFSl6YFn+jQjR6GgYh6upIeAOQWEejiL0Uxv5ZaRATzRB3EcUNE
0A7IrfodXZ/NcdT6ku9d11QF0FMwFhofGeX8l8c1QOFJGnf0mALkFLGMqLrWwfc5A+QlXYzi5OfL
yalRsaGYT47tFDOovPdEDrcBjTBAO3ZIMnktKZ5SmCeWiVOowmR0Jcw+f+F8QxGZLvDBOt05/XIm
hS6k698MAYMR5syjNkxvQ5mgVW2Z431ACeMeJQExZXXfaLdWxr5pQzFnsGKUQokmlpf9QMXYvSjJ
WO6JjxVG+kf8zmiTZhsXyqS8wwhsAInVtSQLadVkp5z6vfMH5ulltHv6POgnP7MNxi2GKdjoFmso
kaq9fvg299NycYg6v7B4jRRToBR5Ai6Ije6f3J0F1MANO/U3HInFQg5hy3m/p2Twcd2tLFG4sS09
k1CWZ4ObOAmd750rZ5viKqC6fch+/Zuo4mkuTGpZCHYRaR+vBsuy5atDaVlAVSfzR8njKsGCs09O
f2Ue/gYqXVDYaAHHhhQMBa6MkzTzdkhb0KiUe1bg8KFlDZGT+mYQK+m67KeDBjs7OtnZn/ox5ncE
nWl5qs1fhe8XuxOz417gPTAEXXplwSQGqZaaEsZdCdiPx1Zawi5LPVZqURGt1TSBmSRyc+bUDT3n
3jV2DSalT/6w7/277aWvdmIFzLaxVoTbr7CgP/gMWFqycuHb+6SJctEtKjX83TdrfbsFZW4uTvXe
lrZMrtJFhiVLclyk4wc62kZYGqMyii3ox5X3Xr0RiMfRNM4RURTz/hlwNjR+XypXB5LHzhlaU9ka
QycTvl81zwIA3Y+jv+7iNctex4YiSwZ6QEoRj12mMluOUF348JXjxMS9nYOJhQ3hYUyI9pCHw6d5
YPNIlsyai7oGr9a5oAt9SiFvnaef5CLUXfwGJAUjkwt8aXZnjH1eSQwYP8wv6sxW24ZlLk/Uy7k7
0h46QXoeflNeQMjk4tFYUNH8AL/35k+FicfPknyApNc32MYSMC/by48RmOWjrdBS6ZR34nxcck17
C/djnUxPFWzuZ2zUa3ykvSpJ8n/GpPLw5R+lN+oZoNxKue0uj0XTKexzOSj0q4pw6/Aup2RxClW7
v9KG94gGEGmxAwDuPNGDhMnkns6xXyWSkpPrJUPpDqawG6GNfv7LxthX9UQNrJReWj1gpQqRn/pt
Mpr1EghPdu8D/h+9JXOxWTt3YXUUZSX+3lwU8WX4b00ACrkCG+ECof0IbLxOl9VFeZUBpPVf9jqp
gvYp3nhNum8rW1KDzGRrdGzxKs3o2934zB1EG3nTNJnyfV/jlB2oyYwS7cC+e582KxWO4UgCAn2R
b2pP9nR9v+B2YFFW5B2D1iCc2gJVwG74VuJRgXrcbkfzrsNPH7IpcxDSZmef/Ju13chcg+7/UUET
6uXJkcvFbWKDySKVf49m0+G4A8AF8XyECRDNFfwy6lvgD1bNqkLOq/8YcrSdWKQ08PED1YP3v+DG
dpcXuv4oAASVo4VavXEL8Xf6hepb0rLw719T3U8shA3t9NweQA/uxfAKOM2YtPrM4bp3fcViHVaF
Q/TMw4UBzfU08yYEl45QJtdFvSWp9rgNq2idpeWff4IRn69LcyDVbQc9uqEyQ7QL4r47JjAe1aeV
iZLE/MK0BoR0N+U7CP8DIXDXyOkIa1oAedfppuQG37zkAawCo30janFI1UQHUmKwdxgK+fNjXJcQ
9hAc29k1SB8cVdFTHJ3LEcmSBCZhfhhrv1969yM4Zjm0SIxu+PQPM0LMrxYj5c+pLxRWMWn0qbLM
nHtN+B1aYHEar8Xxq5FSWZSpJmREjhSHAcDXestvYJueHux78bKPVZ+Rg1Z2rwheNhacvmCgUoIr
ZzfyT+C9+f4UGwdR8mPds+ta+sBHCzTSSyEs8K7WBy0IEHCarDqxk66gh+FlqCm5HtHmWddOVT1T
55HOPagT6F3U9G56duuGX5APlk7dYvtuQ+6nkyrTgIvaa/6Aye36DOhqGtN15BjkMfa9Dienj2wC
D0EEqBS46difL8noGNNOq3c5RlhW8LfP6betMUf41bboSGudF2BnfWhZy19ZSDfSCTVJIaLXU0U/
oALGXoeBslvk4SqERuY+4+A+nvLtyD2J46KGim1vYtys0xXcy9F2VQ8X9vsGpUWrO70+mf8U4NqW
IuUig9o17thptvYlxxcWPU+ZZZXfRO392MY33rSRebhGQAxIwVM33RCyP86qPb/IyhTQ4lSS4De5
LZrebsR/r3Pj+z/6h4GGAhMYqBKMAiQshlxoP7fDvA3HbbjOG0IVL8x4lvdiAwNq0G7OGV30MBkz
7Qm6YL8L4AUUbFkt++R65GYNNhJyyY7YS7Hf0L1q69WLLbzwGYL8x2Tuwvhop2lxMLfvNLz/umch
7auPH+8d5h7uLIJQfT0N4znS7nk5Lrm7qPb+tb4XYdYwWIt0KasdcQOIk53lvpLKiVoxtDUkEL1C
dFnxZQUIZCtq7n3MwnNrzD+mYiUzD9qVaZekuW7CNvxbcHW9t4CLYXepCWeEQaCgyyB+r6hT84RS
UZ19SC5Ngrtv8I2OKmasN8KdvrpQisonPP+tlJdklnXNyJ6dnp4BrGj4v0ceQf9tIdQr9Nm90l8G
TQqGQ0X3F4+BPs7jFDx2qQhWqkE3cdfhoPg5G4AdOcZLJ4SfpII2q4a8TL++KuiITVtzFbadxvzB
29zl04t85zIkUDISPLQA8zbtgX+waDHgvNTEDEMakoogT/7/t7JUTGwJ/qy1UM002SbR0SjwGWls
3X8eqE82UTgkPH9FTa935uBLNvVld0VyjplTHOT6kiC6XYZqv5g6+MJnCkB03Tf/DYWv0uexX1q4
La0uIyiZOU6UBvx+Qy/chbJuGJV9cLfxvAus3CJv0eVHCQ9uJ6JDfGbcuhMw2AF1ibd1xxE0/I5y
7kXVWETLQr71EUf1T0QvTVufPL/0qKhK2YWbKrTJ2s0pJz6mrTQeqzopQeHMsJaGJGkf61epIvE1
/puwS/jfLNuKHTsLjiCo4TgKk+CoCenH9re+J17cA8g8kw+ULf62a+6NhquoLc33Jd/xssL3vL1o
PUjIUm0KUqQeB8JMjl4iQkPJLxqs2zFwDpHgzknDLxlWvBxYskQFiGAVwu5K8EtOGcE7a/juiRjN
RZamnWb0FJ+oEvNtxegPA3PSY0Ulk08xz9IvvuDgdlS1jUKsYR1WMW83ybWlHnM0oeb4tPELJ8zj
DjWHEyz3wcTI5eNa3jUWtXJzREY+nV0xInZGoz7eoKdd2i7UCjlmYJv10SVCfw447/M1h5KmFrlU
CpMWDkBVR9/W6FHO3JFpB1zn2PZy83TbNq5kJSqEWfDjfd2FwSjK5u9VxF/0+eo9CxtN8nK7IPmo
bm0ND57PzkBJzPtzOEYh8DGID5Aqyomuv8Wx/eTHHC2pDSVLqm0O1CJ1MVr8WiqyoDvefAnyW+4h
83DKRwivib4R0v4Dr17A90zZo1TZAX4EQtqF2DUnLjlpGLk3hEq5QCWrbdeaGHhkEZGMNYEayqU3
xILTDhULL3bPWI1xhshP9dbMVmz/0ICdbCNkWCaNFv6Io+9oPFujCu4YgoPfNkgEkIlSHW4hl60J
P0GlZooMGPgd45xa8Ci/p0M+A7/FPDIWwSrvoUBIb6hIk/CtNlhDVYn9HFVEA1CupgnqFKuNy7Ii
7+FbqYpC+Gehx1CFE668MwaueF3mctbGNmJsFBmbqYuJ1BNASwuHixbUUMftIX9rQN83sc5PYGTQ
RyqJaKeprltwF9UeykqGd37kvUk7SeCIePNzkeF0zWotZ6mvdRPe9PBK7YBW7lBT2H1JXWJd2dhW
qS9KmFWCJykzOq8BMs/BCWKi9xQ5qtk3GOyzMordPvPsGL9QkJYnghaFoLB3r89qZoK4KvL1br1F
Bg4RJpAJsBQahGDGeT7ACC0G7Q10XzOkd1fVrX4vKakqwdg3a2Ss5l18bnzNraE4wyTok9rBYYge
RZXAOkmcayJRcjJsqyzwe+4jE75jenkulhA6lCsgTkOwHeUzhGqsFr5HfIayh3CmrbXEERvrRfbl
QEJehyZu0NWK1rb4e1OD36t0xTk/mSr6zfrsUOfExFV6zLCUOuFWe4vfd/NYXOkJas1Ip+1tXFW0
wGjQdRN0gNtrS4IM59f0x7KNPz73mKOq+9J96VyFXMbV1/YCOEfIc8UYgTmzQRCL2eJUELZVfMWm
nba9eVmXNzUWuHnLezW8p6itcIbdp0qmK/T2xm9cAMI3s/acA56Bhd2hfKMyU9GIizAt6fw0V0w7
K9zjD5CR0U8eXgTKAw9/uJl23TuaE44304b4tCrtYXCzqSZ2T6pc5atuRHOKY/qSIZOG1H1CDUjA
9ehe0EAUhfE1QEv2gPAho/qaJD8Gs1eXQpd8r+2UM5xrXnXMkjfpzBOLP7qimCzbPfD2e/+2Gxc8
iN/6oN3ujyBlvSrLoNKXQAROWp1PZuRkO21ioRZTbr8KNyh0ax2mrpldTSk01sAtZTph2ASmHNKP
TV5UzoOJkkfl+O3dmNhWi49XAdoGZgpekDx194irjjPre6hCwBfZQp6kN5yFr9DcKyXn8wSeC6ub
fFdKWg9RBtMigbL2S3KqIbPp1AF06QK2K4IM/EXCRLLRrApKN7PS74hxgNjcm7FiF9U4MkqfjcSJ
aJn8cnbGgJAm0+UuVMqamD4MRB6zdLVWb2PQ3yx2NpjEf/VZJR7VF/imoISB7sCS1rwAeh+Uk+bK
jQ00QL/1t4n68cAILNCnQV20b057NKqWC8oxNDH3Ga4S1jldiyWtfBWlBvnJdlIJPITc1AbuvI/V
UkHvwL+CG0edPZAQM/iAHbrr0IaqFWYeO/f4cURTAJHXGwWzuEt9PIQenfw5E8IhBTihZ3Wgojjp
dhDLwObA6g5krhmaQMuXgjq3mqKllGR6yWWhHEgz0HQy3UNJbtgBirVgTwkpL44R46t/xOdu49dF
UIRYjT6E7sySUKh/ZHfJHzy1N2JysISNFRENqJrAlDPlU1mSJwj7NmCHoh5yL0Dt5M5IMpKjfIA9
6jXOVqt/MOHYA2iwbv/LslPILP5lU5Akd8aP6x/4WYDg1SKtxJO1MdNnLarKQLcFbREfzxxK8sEZ
YiQChA2nxjf3Bkr7uQiNvoSkxs+5ViGcjxmIEYvV7Fui6uPBtjYaQHBH0XDiM10HvKK75sqbOJW0
9P9o8Rr/9cI3Go6KD8bYmQ6xys+ZRrK4DPV64gIng+4DU2/ze5Tdvw/f0h6pxcRXVvbN3+kieoH4
7OB74L5osWSgxpvlumMgnUwaLfM6GH85Qo59dBz0ppJhRdlHqWD7yoIqx2dN8DDpy/3Lgp9jD1Lx
7oNvR4WFVA3EhnczOcNLMWJ9fbs7IvD/+1zPhtNOM8VpOrX6FjEk7WhD/Ap5kl8cFQs1E5hjfsO/
y0essDhtiYx//7WRY7INuxI7OBaHdvehmTbpsKeYPSHyTqmvmURltWNu2pGLh11SZhdye2t1f9Jf
Z9OJBUdJd5o7aCToW2vFt8duLHnqn2xEl3MPU9w4zwQruasVRSce8EB82B5AsBmyawvr9kJD3ZJW
LBRrV/Li1j32CkRbf5BYbkzLrA+IKnrZhQ5jrYcG5/HSTgv4kLUjwOlRTI3PmdMYcriTnbpvqt7C
yU5gUEmDPDeUQwI5CKbfW6LN8ZY6qb4CFvuGVeeL2ElXjusjgjOGi9EnUbBD5hTwYj/swVHHJD26
BSEY/46E1ijahHujKQbKZLTMoXRtecLeNkwS2L1wo+lObZjrHP1mi+Nzz5CVmWejWlblPyHe977C
45Ay6yUS4tT2ylDI7TSswry/qT6/9E2kdEYFm6coj9xgoK3Du9K3Pw2irbqhwv8BgvZnd+cbuaIJ
tfXH741zR+fk8VTM3YE7oZFBO4HBuYbc/e2g2JQb1InJ2pm+ZzYXzo9Z6baugS6qSkBn5PGmpYXQ
2v7bf2hne1nUmUsso1HwZlArN48RXoznMEd8bLxks6im74rg9MYc15FXoDunm6HPDWzvW7pajS2X
xU5k5wfn7Ic3K3zkJhcarsDN3BXrQkdS/G6tQTYHpLSsAIkmM23gH0aWGg7YRPPlwim3/I0cX2/L
kN2JyOQMdH94MpJB5AGwRkM1U/Wv8T0wWH7vnTjjHy5lcaE465e7AmTVGq1kT2O4e/H03GsNAh7H
gtZpJeZgRt55GR7mioKe/kUi3P6IDtTmqcxDJ9uZSRG4ePnOhvXJsRRQOoy1LftZ9/rhhW04Zi03
20thCSQCd4tVtTT+Z5c+cizdme/WoimaLaEPE8z8zUtMh9LzcyRHlUG631j+NfYlsVGb0YLNOzD5
97RWLk5KtX4J2oiM18LswqqR+vg03SfKQvXdNwVNWj1oKg5skcYXZKbO/F7QScfZW6d4N6AC/O6+
nCYe9E6rOXSKXwHOmcXibiRgr5bmhFQiYwQ3yxHS61G41vaBVV//YFnsR8RCJRFmZH3A1tJPY+dz
hNACDPOXVZvapxIz9ltSNep1MopwU4gAFL4MqfkuGT077Haneso7sBfvscR85cAbHQ8PhBClozua
84SesHn88d/nga4EFCWWs8aIWP4mQgM1PPa/wN5cjBN5V9/SiKv24icTQRp3SObnYdEZ80XXB8N1
CYs8SVPlFPmm9SbOVnVy6exLYTm7V3JcCI10Lr6zibpTXaVRVW04IxfM3te/RXEB+lH/jpIexK+k
PARSrbt7ZD2BV2sARJne1TMyMRKq0hi4qjzL6Al11Y3NTJtACwKZUQT8unSeALuxykDSZZCiag3q
NWEJhcHJn8dT2CC4s+Mt6nhYhsPLvxSypFFD69av9vgM9Cx0Oquw6QVZBV+CGkXW3FRWa9SS0B6n
S1pAHHWDeYVpHy2kTKc+4HiMfLQtNyvWnMbrDIZDOGiKEWu+wXD0b4zGUtVps9nwtzswK/yzEP5L
MInXvhR6xsf/SN/zV8FD8MRKgN/W+Nsx7mRo/CYvXQHcWiBHf2YxqQGTq/xvlfres+Xhg/DaTkLU
GUuBu+o+AFCeiysMF6O/xdM7daU4/G2pLCEnJ7Wy7B+On24VJV2S5AhBUHyfUx+IQBtKwZjKj+Je
ENpRd9btsri6LF8UoDUcdnHcoDQ/CQprTQ11Ul8qMv3XRmCKkfqaqMuj10A4bH1ZxlqIYDdQHilj
RTjEmzAAZzeQzVsHDUAqY5Up3udE/1LvNeMcTW44f52scN65eyCB5DPBq9hC8OTPk9eNyhLM+hw0
sakkRsxd1giflvOguXmkJNCfNZ665EFFQ+sUWDt2ci/TYN5lRJ5/R833TA9itdG4dttw5CvI2ksb
cJ0+Q+RjWQ0swq/ab0Zj5d0oZ9DgQ0RhLkZHLfaurCplmRXbY+YS9pU3tnkGMVIRGZivmBDMv2d5
KgS/59xMnC/U7c1NMdBD/35/587yp4GUYjtwHlwZmTQKC1eTxGOkXpijjvTDC4BE0T/8SOgPGA5e
qTdLzREdhCQdAOCFITl1mzzomy0jLu684Tki/jq5oM5C1dOQCbR9dAI0gal6LkLMcjb8QBrpoHcv
EZ9oRLh9qwz7O94cSbsNYX8aWn3rI/bI0Ux633CBWBSRnXiML0QGX47rvVbAB+pGhQtbaN4cOusw
l8Feh3LBn9IABj4GWw8CWWLxl9T9DBuNMOzWMVUHrHYs5Aa/qBBZhjwvIIvyiKwnnLZpwcsMhst2
zqdVat5Rjtj1fpg6g2ZTDMQrK1w3GM4WszIedZCncK0NOEwL6du8uous5/RZ3mGhzA/x72b89PII
DTZYci071c6SxOr5knSG4nPincZZL3UD81Tfe/EbFOr/0f8YEre90R2O02IySYtRmbuScsTHZfUq
bQD1TYdhvYGzugra8+W1T9D4SV09ZaUAx5BMcl1aF475A43GctY/PmC1tunPPjqpYh4nc27G5Jh4
tGkV4k5q/yxU/U3IsqWO/QWatEFl3Sr8pNKHZWPIXqvmRah4+lt2C+gPSIQ1jEwsPWbnmj/bhc7H
U1lJoihWG0D/SzAb6HnAG+GncaVZEy+EByOMrWOG0HIUa0CE/uQTOY570ciqtl21cARnctNUdBSW
MMExQcbMx7jgC6GIZCBeoBJBkun6GphAU4JKFBK7T3iePXZf9XdFCFs4Wih+sE74YOjzvL52ggiS
FOV08ap6p8n0z/WMfT3gYwVrkxY+Tp3jRp6ODyNJ+OU6G0z58i6K5jxGDaWkZ/AYHPE0dtc/ZbTr
ukBhPgiNj9tvrwM4p+1XWbaj/xcvkklfcjfI6+G4smaW5Ah/ADv52+Qsbv5ILUgSiyfy8sL1qnVm
W9ug1nrFUBMxrISxSyS/mq4MtiG0ZOBS0ngKen3xEp0rP6yVd3t1yU92FLAfghvSwHiElkFMRejn
YsB5/nUhXAWgaGu9hPaZrDnKUR3ENtiVcUzpOfWCX/Wa6Rc6xCW56zwEMPxbxJKVz0ybV4DpcUbL
urm+46XVnwITAtdElH9SRiaozTzFj5UKvIG05Bjn/xhblGZV/B3opV54mBbaX6aUfC/rrmJDt/SC
Q3R0UydFHPDQ6N5hjnlnfa9kc27gqEUNjqglIU8xNkpCaN16HoSxytfDM6Oj8PgMv1JbNwIFjnQT
f+ELM2PNClZcMTQcS4MyLEK+WIjCkNB+rmGuzGqVdAHgNjVxqUDw/LT06HKBm4lzRd/2gSWYhdYz
8pJmBpR3OX1eHKK3bMxBqawPB3PqTD7ziHcHtvgSpk3UuXjEANNqNA73ZzErIYOxorFqTb7xOYcS
71UsK9GZDrJHi3GmBWz5HcuxVKTwdbHe8d6vF/M2rBSG/ZsAEf0LgUY4EwCd6NuSOqyIRm0wusPW
acIkitL0fXSWFX0UulT4wh4Rr/+VBsc5jGL+8xSOrSzPoUkYAzgqo994UXmuM3FBguh/vLXnXze0
/nIv3Kp50jCiy+XMVPfaj6Bo4IJ5kqGyspL91kBDojZ503Ny2XANWrc74kElF2qNAQh20/Czc1DH
LTbKBUq7jKU7tLUcTE1jv7Qfmq7Z2LGFdRD+i33cD6JxLnvkhxYvdnm51ydEROfLMW8ygRE1rBXO
aMpGTEuzdTHr1o0tw5QmV8bV7lh/XbXPGHShVw3SA1Qc2skucyI5LAhKClQSx0L80qVmDkTZLTKl
8Gitybg83SWrRjida5oWqoaw+GR35FHCFd3gCUzLboI9v3kUxxG1ZL2lzExzZmMrCVb57bBrUJZl
xlCszZKnhyNwX3Y4NIX6MBxqIfDLgBCMxF06qjxyCtuoECUT/5RE02CPg2xcscksn/2iie/NzOP+
pGW87P/oe00bp7uHaHxn+n5cAtlmRHkfW4YpTLpivsUngpMcJ/jwzZ+mqfAFD5Vj2aU+YbMnbJGD
IdUxX7aUkO2+Gj6q2j3e3zMMTMLPj3i0CWPLWYMzLQGTfjvzE9POVriZQ8PxUe+RD0WihgK3vN/p
daubMr09/KLWm/nluW14X8X8tjAVfuuPdZGaE5eobtt6utRRVFRyR0FUza/ZEpWpF+St8Gz9lon0
2VCFgyx1pTWxz3lnXBcAueAhYy/uS6e9Lo4s6HHjJiNYUd7fjxGBF3l+vwpidFVtn2/S1rxgmSS6
IujClIhTIfypOPKe8STVhF8Z4DqQLrhrBRInWdVv5U5QPuH+KBDkgJQs8CGqAZ7GXcO72KvvFRl1
vvbPnM22RKeWdmQU42EdAwgXyfwmy4LE/xX5V1kgQO0NcnuKAOYZr1mbaPBoZx/KFkITXWRB3Uxj
pvV0xpxkQOEg+o8farz6cOw6i7NwMYt45WTKneRZ6RoL6eiHw9ReiePwQYzB0PJTivkP9+Y+whzY
SZst+S67Yy0QdIpNM9QBWxWqE52cnWWfTgqhx4EQfr3uV0YYWEepEYjbk3u5AaH2qifCZXqk7A3h
4lLKdmRNVctlY6HnTUkplAavcXaia64NDJCtmYNaNIiYklq8WoSLqUWHPhCzl3eMyEoe00BvRvSP
4MKOv4t/4VcHJjMib7lEFGd5AZufABkNeD05a+qvd/Dtpu7KUDoq91MotqB8yBO9QG1Niudkb/Z2
LCLwv0WhcSEasVO+Z33OIZpqRzkxGeRJhJewxdGWCBqPpgr7TKsH7eVAa3U9U4KODhtp6NhEyBff
3BFDJFSmayUyGwV0QDpW9eP+2E2eiV3N3sO7RqfBJbnvkbElxzopwagq30gP0Ei1W+2PLdc1dZmj
Y5IM8mxx7Ny7pJuo2izoURUE14dQJ/UIdferj/dPYQ/6qXDdecmyPz0Xn2l7XsPcEnYjTau7qTfl
SmYEgE2vNPMMeymMrm0IJGBB9bbiB0qO3mu+qxuvqcVfVXpnQORKgTZJqKnQd2j8FfmI4xp2EoJn
rBqqohksyKIJKreQtnK5g0MMUgZ07PQUFec/fYggI4jzXsZzBCBWnWGXQSaR5NpS0PaJ2bldwzu3
L0NshZFqkliZDeyrPXQSkmHfdZzllqfWyLyNG/PWotYAn8DE1td47ZUHPcdBQgqusDKzqCO18VFC
ggaGaSTT626jHmuFF+kqFNnQqCH3Js9js+LP4X4Lj6z8HYrtA3hcBKOUJybCOK3OYTU/S5StMQXx
WE/cFCge1lO9OQ32xU4jpUHhsFkkYr0jM/XTyDfAUtOqZ9YiTiO+8kXniwhKOuEPMbp7DtXst4IU
vuFkfnnMkS0nCN0Yasji04lItCpC/O+/ITA/7rc+NLmse4+gmF/fFZzmqyHtzwlPRPErgvKo5bjg
AN+PLaWHeYSbMdJ5QJoHVI0Vkqwx0Rirg4oCVEb4iCurV2gN+rAti/UyaRdwYCft3mYWnGaG8p/T
X7AmM03cw741qKSudJuTdj0FcMhk8B1e43J+J/C0sYMBbmlxWFdeH1LULA0y+8kFur88czaBC5NB
EzM0v9PJmprXvks5IQrDNtl7jmIJgJjLVjoKzAdu/RUGH2vEdMfUhI0s+nR7+F2EgOb7XEGTAFz7
LvQgRkpcD7upHC+wYNlvB/2NBwRJ/Mn89UOWejBQlIscCV+7vucHqHgKcFHvmm7vV0GifTAa7Zsw
XysRz4cabcMTEa1l5yWhoqYwJl6pXH9Fudf2P3k2uEar5pxmUewwKjXt7RGZnE+gFn6Ikp3Jdko5
lFrD0Kon6CUWtgg6KToluF7UNtrdhThmwjAA1fA4ygvf7Z2ozZRM/6IsFyDqHTf9swozc2Ih9bVh
HkiGhXqRtTmMeyIIbvhPvXTcROM+Z6eu40rNG9OoaMsZdMpjz7sTKLW8QiKVtPebV9qKjAVNJ2rU
fIokbD9kFo8xyoS53/GqKAcagj2WnHjHeY57s5sB8NPwGZsTXJNe4KpVxLE16fj+WQWq4JDMdZOA
1RR1sg71gAz28HJdfOCMr287RU8ZiaFobneSJAnVGdZWyuSdg4RCHGgca2wF+ihIykJxX0G5cAe6
QJ/xJrjWHy16A4B6og3OPFaWXNjDwRy+OzuzaKv5TCZCd8BoFhldCGkcTFFeOed7n1roigM/PTDR
3b8LSKMERMEs4XQoS2ca0pHAvt2QDwbcJ5DmMNkNRXStYIB8J78tm3RBA+A1ec47cHTKb0IEpY5W
U/Y2MUxcdtoSmMrgayjdqqSj8K85A7fk+ZycqWh0VJGtb6IY6fLaX6a5guTH0Wneb9fz3f4qXd8N
byrwV4osdSIxRETI3+QFu+7uqGNkfVT8lhwX6WVEbIpgwbzKkfpRZI3KPLiLILccua9Ih7JICoAd
yU6ftIuTLrVOXjpHBF+2yxmS8cJ813SLCAuOzjIn3Ljejo5vzpevmwlUt4l4PxkWMBhm+QP0d1Eh
Wa5AkDZ8HDhNGEEOHrUMxXDYVlW3Fh2Td4VYwGgO5Ymhobuc06S1jRBpqfAfSrBu+/ziMc9L8Vyb
brW3uIZVi8moNKc5/laAJNbHW1YEykCAIShR3fq+8rr6kH74mVnRR+x0QxCPLC/CVvV/wleYr7rB
kXcq91npkjZvDd5ijwDteXqMn0kRUFRbi9GdmJ59qDe3oFC2jGma0z9nKhFLSie/OVNCogUqu/tP
IHckstVx2V0GD/VVKB6NJ29KXOxZYsuMw61SQyiwVDGwCHpW5DNz7OXz//vGqgdhiml71i7kepCb
5f/OXZeLsxzb8z3JDj+3R/5c9aSrEKlVz8kE1htUGbMJvSLmX4kzTGqSbQQuXt7G6c/w0JXnyeN3
sTkwysqfi5akOeW+4PaySYym054uPJH4qJS6xgMUrfxuSCWv9PVH9as51Kw0JN3rs59pxegFIDxf
LcirBzhmKx+adzKFkk5/2dY7fHe2xnZJnqt4NK5/gUdDTVGmpoxSMA674ov8ivg5oetefUtjZ1Wf
DtqFBtb42HHpbgyWUSM72sAZdvbtrrqoayd6J6wKWJ2gYNkuc1lkoROH+DsQTLnjzbMQ3gXLKTIp
09S/iRNclfJQ7g1UWA/1gIEMizZPtxkqpXCTPA1GgJkVsw4108c1yfsxMWEogU7Ln3tRt0ItZJD1
Zs/f/o0f4d2rwINX+WJAFItmi4xjfK6upuQ/gmVCIriKln+8CBxWiwWVXZddhw+uIWnF0P144C9U
xrNJZIgWyq7vDjrGsmNsiU5+n+FW5bXLPw5Jusjymt9T07Yg+62oAkC7BOOdPxgRpSqNUvVaMYzP
p8qQnPK9P7AhQuHEcnIWzrTTuph1wrQD7g3nTXOO2VqHBbTiYaxrbEeiKt8Ataq/yGNxj5JEfsjM
QFwg3o1pNGn5GxYvx0JeWFsyma1gZFDoB8worPdnAKb51a/qN2hmo1jribx4VV2f8rVcsHTlub/u
h1gpflK4zvU6vF1oLdn+udM/SAbXE1FSvSVz3fFp/CHWSF7KYFxLyG62ZAOva/2m7248/xeHmUDb
S33SPO4Tn+DXAOlzEUGM1i4cc74SeKZPIu7s4zf3UizfWRJ21Ck3kD4gPDkD7je5SKwVDepxwFNZ
HGZ2mpJE571Sm7648uiDLkZk8j8gL7YnL9VvyJqpaKWm2nxwjWPOw5g6baMzjokqSyUkCcSAmdCu
2tusBoLvTfMES1lpx3ag5bGx+kXjknd/kinjwL0dxRlyJLGeLe33v465vLPaS2N1ydom34AQxf25
+GnUju6NXzHleO+uW8r+0jY4kvA9bZ1GTX+I+UbBvzZpqHc+hSrCYDScSVOyP6VF8jRkpsPhwAlB
uCaRRo2lz7j9birXZ0FiaECdrl7jeRP4qG5oPjI//ifZBrcGGVxmLSRDeNuG890lEeHG/war/p3R
tkEA5OebeyWNpvt/Ryv2Dssy/E5n+bWl990AlWckpDTg8dLNbVeEtKS6lyCG/X4dDguusT6ji9dO
JipF4JYfLA1IMeaScDYNc2cUqqYD7h551ySNC5/44XFBchuhkAg4XNGhh3fzFroNn8LBGtNLWGI7
34DVscavfkTHr8XD3NYX93BxElncOgYmxp15XPpijps3MMMJA30bZ1AyHutjcOYZq8z1Zgkpb+ZZ
cBdiVBqzCvOYL9bviZs0lChwNLSKG6PbDXO1s7/KjRtIsPNXNxRXLb4Zb6cU0j1ehbuvdpcGGQ69
kspUfT9Wj/4kD7T1LwmchSNEmK0jxG9B9mJiyboW8c9m8vQ603JQfwrWcgzeUkyTPh5l30aazzBx
6ez67DSM0rk2V4ZOwJTwUPIsUL9rRsXBOCCs3HsAPuhDg4j6RAsemdPraKiBxQJtslGDgkzuW5ss
wseXtsD8d699yynr7d60TpcznYyWbCf13jdW8sosi6imB2g1+pDWAkxW4sm/HIfYoA7zzAuwt7bN
I4bnmznntazUOvQPGjt4AYVmw0UwD489SBdYaits2zO1Z/t2sJSXJwVwNtfYy5/fSX7CvGPkB+rg
6NmxPgjB9H3nxHr3rcfLjd19lQyt+WCNiRU5lDuuUCl7UDeNBsnRTA/DNYMJBAfjwfkCV4mo6c5q
67KWIcXwzZhVlKfXxtRH126OHu1DWciMF2XJ0Yt3IUWUTZKSMlRIKmavbGn6CW+DkbvfOsBOksWw
jsfT3akE5reBHzZrjM65VnxPfL0Aald/E0tMkXWTM9jq75aacYkfwlZaXwEjcC5vPH/UzjH8y26D
/m/yKehO8uqRrh5THzgeknji632jc/LPJVD71vGEBMEUDzeekMK4f7k1+ipPcwGfrqewfex2330v
EF/HMJkXLNZsXKT1Gn/CSNZnKodSAicBJsPCVIKtSKLoT7RYEC2Ed/7TLKO4YKNJPi6C+tS+qsTh
bk/Il5eXFTuArDdAV1JGnjzdNBcUKnf0luzUHbPPXbYp5uHzBgMonUvzXwmCZtCYwGk1z2IRUz2X
CTqeaFQijwXsbF22SZhMkwh1RzT2eciGus+bnvItxrtcT/gXfu+AFr159gCoSHbpI9PatidP6fFT
24AW4yU0zbX2FoL8f6YxdRuLZDYK6mLll41RZF0ZfiutXJuTFr85HGL4ENPYNS3rbBHf8/ytfp4V
FC6+vy4eBgsUvsVMo9gCP12Bd9QN8OESs4brVdA17nSwqdTWj8+Zwh8gactXECfzRuCS1ESm93d1
XQ1P2tVlnRb2YfFfmGCOexqkKiifWYoJmKMeeQChamKdmmSZ8ttt1oPZ2hq5vYBZpJj80DBy4Aug
ABHxBqyaIgEvtLTrA9oVFdExQQSl/S1j2q6xG6kWkiVO50b3Ooj4eBGTcU2BXTXsHIeeYysydjb+
ZNyOlW8mPUzD74yxIid2QMx0s8tHeYc1xPC4/9p44DUX6yb1AA8BV3dOdvYMn6hbm3f3oawpDu4A
0LeiIJeth6IIRklFSMzGXFb6wIvMjxyriC5lFL0sdGZ/lVwV343fxcWQSKc2Z1/pKoYNG5ja7i0Z
z429urp/oXKOnjtljnyY/xUiYKituJmJ7k503iMvLaHxYuYc6azyIzraMNRVlmsCiNcGmjYZyB83
VG6EmzyXszKjt8iB6wgs/zVHKo21vZXO/WhhM6Aq8Ht81XWhH98KSjjYHwR8gQzm+fkvri5mS0EI
t4UTRZgcgm+m2f7FJx4QGCorcmnDeNlSPJ/zrOxdEqy+qncEQQpQq8j/8lO48ajU1+HU1BH6ZcWW
ZC2Q1lajcSAjTYw19fZci1XsWYC8nkdyxGIwdamI2Nl7JytD0P0gU+ngriiT7voAxyomcXtIXV8G
woqyFcK/W6XkDW40L95e+3q6fUPaXPtkz5Gq4obve/Eoajj+tMPKaepMP95wQy1tBMEk86VnDTFI
Cgsr3IkfB1VWQisS+YL+tnFAQQexl9TDmE5tZ3PeQ93Ecq5fMVhtTcwPEd6fNmHrGQzlHBnvjtTC
V5rGkJpYw/CFGQ5gqjMMNe7JqyHAbOLFIEnpQ2vJT6EkG+FwhDCMXkH6s/reQTpQoprHR12yy9sJ
iAziScw0ZX4wXUC/yhe5P5VL/AsbYYhrSTRmEz5m3Jljt7YiXAX/DHgQ89OEeVuyV8IcupKomAIZ
ts4PNjV0/5I2L+A5x4yNqcxD830I/kMRyOH+NMCrNd7P+3sD3Of0US4mx8Oz/4AAl+M/JtqaH/mP
7O8SlGU0NEm5VZRDnD+IFYKg5N9AkVOpfzNN1kOajg3nHvoJnfaaVlFlAKCo0g3P7HBNt+1JgKuU
LAv+WDtSar1dkhLnHADOpa5uWCd9VxMyEdhVa2gCuny8vOYkFF+ZZrb/CdJ1ZKy9knLcL2BneY10
J3w3Uzrz1DTbodRufIVdc0dvzrRjxRTMdML9fpra5oGPllLVBKHp11ArEFM19BY81IZMSVydwG06
LuUwPur8nGOQbn4icy53ej4UUvTdoQJVuG2UKCti7U9Qrgz0ma2UabEnGmIXoQXbft2KEk7JY5Hi
OPyFChaxpGzXhoNJr5/Kbrx4EuiiVqr+3Z9IR497HG4NFCe+2KSWB21TeE5MCjoXg7rw2GzRnXIk
YdRbBRdHAP9gi0UiFtoCNPHIaWwtsJFGPhyTvUzvywPsXLHrLPdK+UXZXDUCr7AF6TH5f2P3KxV/
JmvSNmDUEEg+/tBKBuUgvVK1YvVvC/zfizYo9STysLniqu6t3PjYUGAQIEOBVuRWp8stwbicLD1a
+LEDI2dAC1QUMg8rn+5dAWptz9APvTjiNNKOmF20XVJrG3TV7705/9e0UzAN6oMCZbJTpumxGOXy
XRbNsmyQku4tci9qvThnvE0d6Q0Wkh8+AsNe4ZmrF/bzRCf0t1BnXUz3z8DdWDbBLyNjU5TOGJze
yWnMcvUeOtPV9yGWNinIMC2kMZIXY9Uv6zOaZnRK3dcxpblLAcSwBs641sWLG0/PVzM3AX7MZJwk
zliZ86ROOBa1Oo70ZbKr4x8BMYA9ZKqjRB+0jmwfjJTU7pOFXSEOgM0E5t0AlaIHmHoQ0FS2gbEL
2+bcai7dqiTbDZwO7AIG03PJjZcX+y5yGvrHUshmgc+oer7y3/8L4xUKuy3Ff0HgqhAQBRzarak1
97LMQrxMstQZ/2iklTnzDdqZy5IXOSyP7uNgPcTS6U/1Y0NP4fDUf7gyayq9madFYjaV2QQoiM9u
8uSGNDrzvjEjk3GAawScQuAIxFYIHztsoznHLYl1T64SAbUrF4QJ2lAK0Q6CFcqXnBp19gZyVzz1
lUkKwYIRY52DlkZ2uBdMkDxTF7wfjJ2o69WmAyee1K1ciDTzcCBSJyvxmVtow2rtzkJp7fLAFiMN
Owv2rLhY7/jsymsl3fvh8wbMvHE4+GN7sWpUdToEUs6yylGtagZU3WWDUpOx5MoPVVNb/vDhn5bc
mnzCtbsoS2+d9UKzqTMtN+vW4oRVk/fzNrJL0R4B8JXhVRLOZUfjky+ZwVUdp8lK1LFZdh+JI+mg
wb289RAAnuZNVS10EKpSsVvcU6vEDERCX0cTeowTQ0NmJWC+G/AuwhoUEsccZqXXwZTtj3Jngp4G
Wb8vMRMWHszgSirT60NS/Z7i91nCVoLfWwXmkt3Rs31QkaqVBJXWb1q9OOX355TuczNS1PaA4GoK
Kv4RoRO7OHQOwI7QUzeiGm8h3Zl2zrgpdqZ/XN9kbFxgn14m2OpGvazVkICQMT5nDsrrUa58jR/f
knQaQDsSshoCSi6ng4oPZHPsnixIN27y/NUqwux4dWAD6EmZuBxx5cE7/tNQu+RUCURL9Q1p3P59
zpUpkfe+o3CbS5wzkwJ9hi8wth92KkDU5OvrTRf94ckpWyDtujgwcqT/I/5OtSU8DP6YMWZrcSKm
bXS6mXwB7bqn9B9/7FEpCYKpCTWSSBYjZW4EL6FCr4LZq/xRUJdv4C9ovG85TD9lhZSaVBexfSrf
7Nyn4PT2WovdxFuaio/67FeAhlOQPyqdR6mA/aF9BUgXgUwHIq5m1e8aCjs73x/0omVMBNSgVzRQ
QdSceduSINaK1t/gQ3hOs6RAXvY6RV+7gd1Qu0fqXrjisZFtdAtwitPvBTXcNAdFX67/rK95z6m4
dHYXKTCYj97qoKJNeUYODtgo+IaFFf1JORWWJhwGt5VvYhKJ5YRHvk6I8+Av9OiGS77bO3K5P1Ko
P5HpA0eILUTGaOgSRumm3X/tqcZh0pso7rIKd6oHxrs1j9kMH60iKU8ncLuM3RceIZrg2ADBunlr
4h2PnGkXBqlVscM1SsM8EYu9xUXx7q6eqmzX5VHjS2/ANsYV1AEcB/3SjTLSWY7942LiIDbxsML/
SoN9oyUYavN4UuJaJBTkqaWVBzs6EYiXv0bR72katWVie/CTOcIq7jb542WQ+mf5u6vAtaFrJQK4
CUTrfZdAOxs8AMYC2Y8E5it0lQVjpVL2rG5l7WO2TdRb/MCNIWvNChlgleFKqFc7ShQ4B9+eQ/Rf
P3++1HHgUWFo4eqyNDFnSb6pH6LB/d/+Ef3SgR73peESHX6ai8KR1uypwID+TRFgclrT+10kU2QS
w8qbPZXjbhvhrnLRAuWkOyOfN45PeJQ5uWxjKVsQQjlhEn/prJHWr7Jio3OvSIWKvV/v+KVr299f
yhCn3cdvrfd8v8njrM60A2PNIwCff4fTmCievDcMBq8TfxXl8DyeZTgny4m5ra70d1doLpy4Arsb
OgxYY0+VJTRdQhwWisaq7UaIPPgjgYCfaGjxU0yQGWznmCNmtaGp/FOPEz2YrqSuZsoA8h+D7EMd
W1NPi79XeCdQnG9Co1p6xmJLC2IZHR2nV12yIEzPpDPesxIowIMJhs8sqJECtvkj8xWfsHsqC4ic
BqoaEPCTN49JLAkW8W8Xa0xrfATMsZ3aucXEQY1OwRzUbUNi/Z6MfTHyOXbQn7aUSE/Djp92t44h
28HmFTFzCJNf1dRfDjlaVdcmMwlGdoUZXmQb8sD5vn67SCCthnwdhQlGZUaX29DCgGY0TucTniTE
P9FWylcKYOWwFeuGjqppWmB3weDBe2TRumZYYn1yLnErHylc6Kg/3Xcg+4GVQERDa7rUT1WkouFy
tV18bKMOC6rAXe6uB5VU3B7tnvIiMOv1Qqqu8QR4TGX6VqLYu1zwvxzrN6hSvL7h+uD9JzVQf92r
g2VJLrYYMv1sL1tAmQjNmQR/Ra642wtbz1c8VANjWQYjhJRBnUHi++a+v6Hd1Ei6NZCFT5sJAcrV
q6fIOhxEIRkq2XbFSuJqcxkXe1o2jSEzIYRgA+QmkPa0zZOeu/iG3Lk+ADJF8DQ+5Zwie2RVXCDG
FFZJB3saBWkj0ZVfP9U2tXGJbjSuPMsJ3aCGpWw2Hq1PnSnzLytlKAQ0qvRPaXO53iSxL1vHHy1P
yShlsNlHSv9oaOOYYzMsN0HXFMi0CgSb/2zziRiQPqRidYqO+BfAp/jZRktZ/zsviOJt7VQ+GUFD
H5+NXeW9jTEXyK24syktHF0x6L0tBSgFWwYxdPFAEDZWvp2HH+ak6IlZ5v7R0MVFOzbDYVL+l09M
3qEEVEa3eFx9L49FrIDabHf2DlfudYyJ0k2mHxbckAJbN7MLKzb+pPAMjymeYNKUr6Ib42iXw7Oy
rIV4ucpJmanyXI/YFzryJAgBMOxoLBqi9eGY+GWQ2Ke9GJVlqbp4iD1WGUqBYZUBXFupECXxqpvG
P/hZVAwIp7NCh+8xw0M4YZ5r7N3adLLcgikS+PdBr5EsRcA0KttFdBufxDMcLcB4hxmmftM9ObkL
KWnRanGXFR4udFQlKqXxX+WTvFojthB3I6MaonKhGmTMUh2e1VN4hOh/fW9pIPGwj5vCORAN/lCF
3aR8vA0hZqUslTMvoEI/x/YBP4ulldtNib5bzvo7D+DwVo7X2kyM1Uy6DdmJonGLilBkdSqjO5/i
2CnxV8KAMMiAW4ycStsSFYPC4BUhtVDQ79vcSFQOHo913KrcUMx8car6xc4BsXJ8nJBak79TcB5u
syszN2YpcwO30juFjPz3HMH7yVuwNfhoGYiNwuWxqDjiK6NGR6mpJE9cxVPa3IUH4yJUCeGmeik0
/wNYuLAim/8Wh44zQwZVOhCNzACWPwxc1l3AhpPjKxe6wUkN2UkOM4O83Z3Dd7JRSI+MpJcvSgrQ
zvb1cJ1h0amBM3XfJfrCfRwbu5d+whcOS8wTfSZh/zpd5kB9trXHrIqgb524Zks61OASEdH79JUx
QiemW4XGNuMdm2KyXqyMlUfNX/7+qTwGnj/jafXfPJ1L6Shj5C4dq7AwGciemTvWg+eCybwi8SJI
y19tjtjm7f/8049S7W2V+ZiGpGJnnH3qs2Xxr3dG9BlM49Go56DK/jEtaoQEXob7fbxGlgrTR1I/
HUBJpS1wMXZCgrMum3RRCYnOLhwzMNZexe582iBg5mDhu3/4CmZl5R3sJbX3+3+aiFK3e1Y5ZHIQ
bh0Ovbhjq+A1kL6M/r11PvQZDWqNn5F0HZQvAaJaX2CGAXc/t1+AW36OEGtS8jfZozC3pZLc7Yj5
ImeVlFaX8vkl4X1IAZTdVzzs+7uYRg6Rr0vexZurR8r8iGi6ORADxK3m255g6zIg3+jCVK6D8HwY
Sh7ApmMTlSfINZTzARZMkAcKm5kIP5XTfbw1bVkW/054Q29vhJ+0fIgpAX17XBAHi0s9acfPMuNR
gxAPDlqYuGHyTR+lylimvgcJKsB+gLYrnVLiJkcUefOVXPkrpPXIl4EDRbVyKF3Cwmw9i5D63rKP
hLI7WCVIEj/E9CTdhWCHad7KnDMZ2yM7cSCVNzh6xwmP20bhCuNmXhW2uQCAAPZBZZR6N9OGM2aq
E+PPDBnt4TOJh0ReXCcTLg3LePLdIOS5EULOqQDPPebx58VujaqqAwDjlkEPq8FL7PaCllr+lCZX
TBvPOqA7bdsKsJbQLlBkqss6xDTOG9RjfbTTAuGdLoDyWyXnxi6S885w9Y8v97T5ZzAOKiywGe3k
PKNXfKMect1UD12mgl98qmzDgGlq28OtwCAnOE3uyjmwmLibklCq/WbyvE7lI9FoXSjXNVi4Qnx9
FsPLSrWm8c57Ad7xxRAh9lyVPv9UXzOfnVR9PcXFqPSKtCU6Xvd15zPSgmfY8rY2GXL+20ErhVv/
CQrTFysaArd3fbEegpgDX3sStrw3trV58eh+Zrk0ZyQDdrn4/sYpHywl6nBs3x9mulhxXWTx0RvQ
Gxwy6CkKkbRC/ATHNW9ovelF9XZ7jrOAgEt+ZpVF/b14qF/GHc7lKAgIxSyDT0aLfabzpy2sdS3Q
gl+2AYsM1zIloRyO/w2mLRMeqwy3Q6IF4WpVCmYmIpNv4MB1poDdkxR1t4zFUTIg5xEqlGV5afKN
dLaFXOdUdjeIuZxe5QgOHyYapAOHWcm2pDK+7BkN5HoEp5s1jy2rhCX0tu5jQCV+h2Nz/NI7Fj2D
qq0Nce7/f8ToxfvPirQYSg7x1YbUAtPUMYGaKW1tZDrcV92cW/yhY26MlH9nuSvZGf4xFZtix3Y3
LnBOsAArLmiNzEk+gNy7/Pn07q0aOrRxGWkWQ3YtTtvnG4xRR/fRqK3a3vdy07PxWDcRZSS0QUnE
We4FvCyF1+9Z1y6IVbxmaBqR39Yp8whpN5FXo74JxY+cBaZfFuMN3LgKEu8sIQ9Wmk0WDxPmOolM
DMIr/lvZRq7Gc+NSJqW4dL91wygpFgfigUdNTtfiLZH55OHlegN6mrrF6A1ZtwvynURjaIucufal
1FcTILxklYHFKZWjv+pXBply1TPPsg6vTk/HM6MAOJC4UNp1Ch/EfzADfOXAe+wySOKSRiIrZl0h
ocNFhH3AXkGUXB9MT/EeuWzj1FALR91xZfa/psE4ffOfIxlsPlb1l9t79bJkQ25ZN12MuJdZnMQ3
H3k9/TaPMGTu5XUCi/T2dei5FJu6OV2IeEFu/GuzDpOOsbUAsBKDrc1u6Wxtp/lLOSuYuIE6uC2/
0xPHFWXZZFrTsVlusox6oOjZhmci/WEqAXZosHCvepoUT4Qr4erIB6NHH1sSjd8dOyl+WlPzqSsc
eT21pD1AW6yFb1ANFS17FKoihQM6KxOLjoomssFfRgevhl8w6Iu6IhXhz0hqc+Retc+v8RNEyDnI
4euUTtAIH4gaOTtIevgWb03DWuFXkLIKOHKcjEwYHIc8nPLaCvzyj+L5wbrjeW5hF+rnMPwm1v23
lrwo35Y+fRrhMbtj4KrMOw6y24t6QxD8iNBbRS1+2zxSdnjNdV133i9Cv6gGl0NSCTtvK99FT74o
VPDWoAavJpedLLWtv9TvCpkWwB+Gs8r++YiSh5QF53fyvsTs3EF8VV1WHhJydy9b0fpP3+gMO9jH
KQs0q0je6FbBNZlN8x4TSHFVpwQXUqFO12pD382tAYuVEreq4BBC68sH7zqOjyPeKm31jhxckAmQ
sFnoGRn6kn6uKrXatDXXrpEXkUdCGVHMnFS7MddwsT5g06kTEEEWUDWEwH4mCq/2w9SyiZzxVD6Y
DIfyFZ/pyaNNqHd2L01rJ248W1sUxMUhcxO5GAaQ4utDxix5Wycayi0CIvAWVGJCq/lyC9DMgOvX
zdvGvRkr1Xcifn8jlIGyODA5Uv2iqdkxCQ/NGuj9gsoCIHBwYCML3P/lOqzLSgK1DVGeLqVyXKNz
ZFDkmnrFJV7Pe/ETV2vw2jzU+MobvpFUyC8yu9NxAZzX0NBsHCoE/yedgRE8uEifhKcNs4U2b7nM
NC06Fisn5MrkAwbtDbHlrwkebyYGkFht1ogSiM+OMyGEQtEL5Bci7yFQB/O2+oWFqbwE5/CXixrm
cLtfSvzLb0+1REVVxxNxYhIIRhUCqzLmoq27efdUvfRwBUHWwukhw5KHFTe29hOmiL0+SOuIFAIS
lt5sc4hIR+vyYn8XQI3pPknF6ZClYli/aqD5FGlaEj3sF+jCINS5GmyFtyEF/92BGNm30vrz4flZ
hkJUfoEjYPdlsBnMddMdv/Zb6WbxT7/eiDmiHdXHFs51nq7mEjt+mIQ+kT7rrCB5mNaO0wPlL0mY
23O2p1Xn8vnkxOe+e3pNLuwvz65/8URSJ/G8gDyapaYcRpt4YxqitbDgGK7zF31zOMR70koMKynn
ehfdx8Tn8fb0LU3Ms/c8QMFig72TXO7eVc2q5EYcnD77g+RwJdFL7mLFEFcWyPfIrCA/u4QZEklA
atYE0Bq5mlsn4zEI1yJ9/WyC1MtHghhjZnTXZr4JlDCmEYGbKpTFUmzA3r+BXZLrnpeC1JlT7/45
AQefoMpp38HVxhg1jSuShARoMjq3IM1BWmhee9qkErlblBe1U/NS5cyaPpFauTJyRGlIQg8C55dM
lIRyWn8svApL9myS47yQZZbW6LWkN8jIPuqVd1pXrQdDKVsy3j0fjSoZ1QhtxT007PuoXIJ0QLLa
zm6gCe7IlFF1cvjN0D8qbx2eMC/iIrhVueF2EpVybfi3PclW1u4tmtilaMHmQv2N+pSSO3s81OFO
kaHjom2eZhrrcvqEIQUaX3Wn/kiCp9V7dCOUnEiSDLg7gxG0vm0Sbo+1U0PF4yqbVfy16K6oI+c5
sA0Q0b2NkiSgFRqlr/81Yyttb/KEbccwAne/udbqLjQx6ewCGc7bp9xBpsaJOP2/wPfALNve22tQ
j/lsm97/C8s88Qjzs/xRaRhtuVVO9XmitishbzEVVHsyDfJV1jBuiqckQEP6nfkFA7V2DxBJFKGr
EvaQTA05jw2pNHBc0tY9JiGxl9XINVhZ1HEb10H9g84p94zgI20UNxX6QM6eoFW6CYQ8rCcqD0J9
9Y/XkBvN9RmxM2sEY6gsc19A0G3cYYhQYojR1f44/HVSxMErRrLMvM6j7r4lvzszK+VzlFcez4RO
BO0xbP1faeOje5NIGaKFaWOc9d81B6vyLfat/8ilBpobn/EhGDbQYVyhXU1sf6Gg3qdr5wX8nwpg
gvkYkk+XzWOa19DeEGdBVVTodKE5ULj/mQuuYrF5942c8KzyXg/t/4d336BYUwUPRe/kGhhaILPl
igiQbJnsDSUCOCWy45hkkt3/CzbGDPJEJGCohnrZ45fGoNQAX79uYk9r1qP4XNWFt1SHbw9AJoVW
JJB01qEeTz/cIotuIMglcD/HJRxju5+OZ8RYzB0rACn0VNAu1gWfz3Nb8QtE4ClKUeZwaxKdP7d0
BIa8np3c7VOpwka24MpX/heZl2O1gIEp8T0XjWwJncYOeIrXuoCpbU1xFodpxzLk8OnBiyv91FUb
xTUGIZsukejZMiPlYu0MUyJT8So35t/9btNQJPKZ8vGd8Jaqw8u6Pc3jXiBcacO0Ecf5aJ2vIlOG
hpSdsGu9fcPraPNuBR9HTavJVx5IH/KEV3zDT9LjOZIiI4W+JZGpvqmD7DPfPpyd3JAtB3sIlYHY
IucStCeuWMx1dSvg+3vEdsIX6QplF/aw55RULZqh1d5JUd6Rs1q2doIqe6p96CDV37HIgt6+DzVP
IzKqTf4N15ya+E5rxaSk4dnTFFXnovW4pvu68RcRtaMug6IMVEvS9rCF+26EyJEVhna2Z4cZzaZv
ei/erWmEdOB3Xd7yvQmcab4QBNeCv8zwpHiqJ+AhhAXIyTsuyoZ7s1ChWOkw/sTH2BouRNhyMRJj
bUxPkUpst/bX4rSXHWzI03NiQtX/IU3TjVlCCVehAkzb1MwiLRok0dT6ULM/F+ZzYGsgi2UEAyAl
BeUXnMmsdV6URBeAYJ350GedS0Y6rHBK4Bf+svGfLpmqPNd3FILm03aUIkywgJ0md889X3WsxkNO
OGudZnapdHC7SOh91sCKisLjvv1SH3gv/YTWoPHC2pvJ2msqFkS8LtSh+D6zdLXy+b6NqfdwIiHm
DDUQrmdv9TkOSzEZXeFI3T46PyVFG4gQriHb8T9Rq9dp63WvELvxQGPfnzugvaW9NftUwYwaru+O
mjzZKzdXsPJXYOPIC3QuioOyqy+ZtIb7xqmFrJ9YOnwwavae3eqRrGKxcpUkRXu0BGBnVSmiQ7ve
9d6uLHwtFVDC3EGiffV4NEF+6eFPvpOIElaVNu+Do+r/KzUBvq+8HKwEly6Dmz8ztinLHZl3AEJt
2kUf9oVb9diMkMsbTQlL2lco4whVeNkLj0JPr6I8dc1/ILmpOKe7T9mFYexw01Mh/5eIK3uIGsGq
USOhr69e092VHaGVHId3L+Flc2jHVo8pLGXnXq1CqCYX+b3CiPKzBMyRKtYgdtfJJfrqvIFnAzGs
YCSnaSc2W3a/WUNINXd9eL/jr9fZMmh3ne7SHRNaB+gktvtfUYGloRK2mRw7R38YjiJCcaE8slvv
Du/kP5dYj3ZKqil07gAGnQvP9gUYB2VV/7FMgHr240IQPcj4IcJX4PZ7ymFki+5DmpYgERv+gV01
VeDlIyGTdc/mwWr2N9YjqpZm4EWbyH/4mLLCLB/uudWLRTWXs7sr4DSYLsctT3lXx92fcRgGkd/C
bIuB4Yhe0Za4HLCjarjZYYMgzW6jFitE8TtaE4K0vU0oCqEJiqcM2vtGqD8P11AN632Y5OMGkjDc
6idvReXsS5yeBdTe5VF8P1M5YbADq/LwqHimnUl+9muIYr+VOdGOCSNKowBhutiLbpU2nYSCGyjF
GpeHVM3Zz6U/bWE8DzyvtkSU8mowcQHPYliwQ/U3NsxWmoiILDioD1Vf6GyhS7L2Xg6o/fCV+yF2
GCkwafyvBkQXxB70yxhTOOzqIPO2A2vyEfp3ZUSMCGN+RhRxwm9rsDwrXCYWch04bZGIBc+WT5XQ
uAWPtfwzK9abqMJ5HeFidm0mgDoaNLJjKi8tj0nUaoZM0NqtT/BnKYQIr0/wbbYWhAeiQxcfHPe+
3vt0C+2uHhImvG2wff9COysDu5EjO0urXfG+OSLbwvDDCEHucJk6X4oKG4fDcIRH0XoWR33dD/Lb
slRCSwRXywu8HIpG3rgt55KQgQwJis4sWOPkxIq8G2wrwHb34mFuZx0rvXL/uL/JLYkVPA8huphK
u2gZxVqDmybIxP27dylO76yLeed1ljvXrFh/pqDggMiz1knEX4/7Emhvafb32WHNR+7eVu9s8q7v
62IV/1ktkpUxZ0ycUaTTD7xN/rypeKuJAhqU25zR0YV6wLlAlV4pyHGc9DaEuerWqCdsSO8PDVxu
k5J6Egt8ysEr+JzWr5XXFoH4iLr8ArB6zCwA96coDGvGMEsfn8aEhx55SQDNGxcj6EwOB19ip/B7
rQIBDKa0bJTw0ip4crh+XkCMTNi3vPl0FjGcyDC0BF+41w0n8dAjfvIDIUz8f8BtaI8qyeO95Mr0
qqGEj6n9C181miF5A046VTXA2Kc5t8EWe3QQCPzucGAAO/cPN3FzegpKGJK3Q5J6b7/xWUXTZc2U
NpqsLSCEMz0J4vlmgGQ/4myv6TQqJFxxXcDDH16S+GHR1HqV+V/HcgSlzgnEGeD0ZfdEWZ6Q8P/e
EwDzWKJlmufZA7tTidb+eKCISDK9PMyZQC67blQq+nRrIOcHRClgSwhDDGyFzv6j4iQ2RSXRud2k
3n+WN2YnIkGv5NAYtHxdQvd85GKL2bgCN9vtrc59JkI6RXzRimvc/ipZ8+/0w/R5WRtSlyPzZjVf
ks1dKngyfGL64ESXKGqkxf2Wkjl/p5z4LG3/DQkM/QD1nv/jGSkmXIPo+taeODP8FOZyojoW9m9U
kNT+9ouMnZVR6PVPeBXEuY3Nut6O5vsfdSoEVk85kqdpi7swmIA2zeCaiTooLyKrUFdq236b+3FS
21qzFDcRo1OzR6i0xhOKdrgJhG2D652KEK5/Acn4+JfmGoT/VNTo1BCegJGRzyVmKfKD/t7dpQI9
gQQP0KFFQKeJbzqW8Qs7CXo07UpD7TTxdD+LDQpfZnU004qe+JNUQelLG2v3LuBw7SCEN2i3iohx
m30Huu2a1gwv1Pk6EXjGn40N0Gp1gZLWmrgqJ+QjqAuF0BK+BZmZ014g3B6mF7s2Yjz+V87QbshH
Ri6D24D+ojnzR8K+X/TFRl8NyYgQPAHdlwVu+OHjKypsMO6vLxj8djagVeY/4+Oeh4UU6OIOOhU9
lAK41l9QLqDcnimyITSxPY8aRovyYvq+fmk2fB5TnUTdV1kDJ12gTMEhr7S0z3+GnfgpePnL5Y7R
zdOJ8wOZxNJdxGw+vM1ufGAgg3sY3CMRrzfpqIDDpoTGCNrqIMXTuWApRlEvIjP6j64fT7yp0d3d
02SZuhsF8l/ImP7hbJxMXXa6BULR5BCh8V4Mx3rmxKc7TYHuyzt8Cgc70bcr70lYsMhKQi0dGqFq
OTvqyIHU3yXbKws4VmvVcyWXWYtJyV8EWifsjMpadhrGmEVYtr3EZ1Wpkw9F69+VVPvq1rJgVt6P
8m6cvH9JUTmv6uxk0PtfiSLFbyT2ob1HtogMLHVt+fojJYtS0hZxAE2g2dSrOa6M3Fr7Zh0zHZLE
z6XU0UkOhqhT7wJ013Sy2ocJkpOc2zJgbqpz6b8lA2is7Zq3n8fPwTrYWwYnu0PTyS5+OB9pbeYq
J6WAg6bs0lsHpOFhXq2NyVkHF1gdON6fQpRNjfJ/K1Y1+ZtAYkxk9nZ8OLu1uqVQSHw/wz0Fv+Ol
5sev9LzWDmiMHjS6lH9cNYNcsmtQ/KszfVSyfUAxTIaPaovKIdl7O2OZ5AbZg/cclJj0noL8NrCZ
l2AqWw7nRxX7kzn50Ub9HEBxgxTs5V08upgBMAT1fNpaMyUY6jxTuupp8V/bhhV9LpibvkW7BVjd
RW7nTmIBlAf8Y07LdodO4WRM9NuvZfPr+PEoCNSWMQL6za62gx9Wk172uWTLTQwT1cmgVFr5m4dA
IR3PD/wgQg2MYZzL4uMO9E97PfMmO7C8y+Jm1oZuJDSmHv+Lmy8+2PA1psqyaw8gomiPIcqIlVb3
4ys7mcOC+UCUARhXB+9wvTtDphAabgN14BetqE7m5QzGcw5ou+dodwsj3kCnbDIJzgr/esQhsFSK
WxPe4T8vUeRSSTGPzUyflyr4s5cQWE31WqswQFLKO/QFr1idzV6i3Fv72RvuT49IsHYEP4s9bXW+
MnHzHZ1f/Kqs7e7pjUuqt0iMaeSxnDM5nbr6zrq1JvJP2f3CgTtTgHagct02BbxwXp4azTu4PSeF
Aki4k05ua4U1JYLcLG+RWOWHhBCVL98OSRuxfFQzai7Wh9jRSNdSlacu4puQkRn85yHed4Ktx4C1
+JrGataU5lNmBfeKLyGoxHLGYd1E60muWp9hHbZaiSG4v7nNEiHiCF/Jm6ksmkwEnN0lfq/DdCz3
L5I5ch79rMAWt0YIdZIrkbWvR6fBGGwke/HCymdjQG64tsGtK7TPSBUmA2sd+38qycJxFah0fedh
DqtbZrkC52ZXgdoS/8gOMnNPllQei84s9USxTPcXbj5m5vf5CpqP9OJ0eBG6iUXHJL+mIjm73Giu
mnIv5HARL8IThR4oApMQYDFC94ivZJywMIt0M0sHB8ettJgaSGpLdxlfEgmi4JHwjilIG7C1YRS1
Y9KaU+OW4nKZqIdvnlVQrO1VB+O4xjhTl36y+7ea68ppeeyLGyijoowcgkpWGgSfYQBmDORBIE2W
ckDRMfzGGyuHxZny2oCRE3RtSQGjqmLkpi7rOwMOzennswEy24Peydy2w2Ea/3S7+BbNKGFlVhrk
Q69tYrCy2iRvIxRhsN7M/udH6LHRh1ojtML3zA08ck1wmtRrhyNNNhFDseiqdozuAgnzNET51+23
/1LJCH75MPKaI1Dr3VcfMp6xfSrbOZ91hjqVdQt+93KRKeboIhp8NObKAW3xkkRchzQnwJber4V2
UBd//Y8FaxjlbNHcpgh3Q1NIHPAss4/5M53NrlL/BA1eWsn+yYYhciN2owmtPGyVKZvvyqxYE5A9
Fb1hEO1kHgweAF3dWTS2iJMC7n3v5tV7E+wluG6GgBYIgCWKOJgfpoN3BACvMtUeQ73cXP44vzgl
TbCAXJDbwiThtqgR9nGO6qfOhId+fG4yGAHVRn1xElZyqmlZ2z7njYWepeKrkp7SWuGFx8qwnA6u
jBbNxAduc+QDqfkGd+qIiaLljjFoKhyaszVPNvk4NiD9O2xd4hKn3gSg+vVdTtUWaKMQioIK7Jf9
qlWZO++OjuKogBr8AC4Qn2HXpzPcL2/xrPUI0pFhWwX/RdILNDIXzVdgkR2O6isIVByf6yXUXm5A
ch+cyVHMyUReltcT0VUTBSFJ3ntNWTWfVLSjCJxb98bXRncIFkl1EGmiC/G93BDMZZWbnzI9gIj+
cw8epqEMp/WOceg56S0TOqIsNfIQwrkau95942skwqOX6CnPtVz3r8kZhyqBGELL6dOOWIqVmi5T
k5Q4S7mDng3ypv3+rMrT4ii0wKy1dMD4qk35gGtipgMk/4LGKliszVaJCfMShQY2tJvNZrqEnQBm
PRg0pWNPFSaWVThMPw8pC3sCjqR2phPc2YXB1EgCMyOH7Nw8F6Z0ehJlvZ7CNsOH8s/zfajtSvAI
d1CS54V2GFO2xR+y+AC72TkI8cGOwJH2luiUieG2OIv6Ne2yXEI7Hx0IbxlxhoSVTEprGzD2w9lk
KDdCxZX/3YDQkx2lEVrldxUein4Xx+52uZMcWfYFSB+K/vMdtTTMnmf8TUhbjWLIoQ4zaHgY3qmS
UOkzTXOys704yISJRgZfzHr1TrGolGyn0NKVSpt6eKWZoaxgg4r4TUKqiXf2uhYmhRxgXDMCTn6P
lgKBA4KF53AIGkVdSgmQYjS826s5Hdya9DA1mt9GlASxUtx27BifEC/wHUf9fxPo+3K1sW9XWzIL
iqjipLWwnOdkvzb/n65YsvrneWgTD30c/7Y9SX7GY5MNVVquUSy6HqfuOJCKtcxggKCtRSB1AaHW
pQiRIZ/xFJ2G0K46uE4E0OaBXvI16aXkIiu5l9L1DNt8EzfzUWYVtH+vMybswhNxgtoeJsQ+ue2K
WuxeDqv85tVhvtl7xN0fEckU8aMVRoPVSR95qMPOlIXE/xKB9G8nr1ZJHt/ArabyKiLUEi0Bq4Ws
yaesvt9879fE0+YUwoTLmmanNh730sR7biDWbldCSBX5j+HJA0finALqz+Pr3MHEUgYl95sxySX1
cjMm10RU8H+YeaoI8Hxn2TVAnoPGRvspVVnBmCOtURbELtTVbVFCknZlFTahCgBrw3UJv21CQm8r
tNrqgXGBKeZsgo/HQLPQks7Ir6DaVYsxpY3PCoQkLwlHD04exFqIzmq1Wn9lnAk19hCMn3Y6/N/T
CtasaQ9p8goHUvcT2PJ6+JcajYFP6ZBDwO6ddPoMWU+A56W9rfZtvxZgG3cKyXaj3z+/O9aMkgtF
RS4Gmr3tbUzzL80u52vet7NCHNNmqrMdw7/ez+O7vBIV2EpfkFLRrukz5XhO0w1PVkDCyDrO4Hgm
/RaS3s0UFfS4HWSqpa7m9ettkj1z81DP21ECvjqTO9dxy/KVhM70bOX2Tolow3d630Bbn2cb5Imc
mrASi/bYTiMPtrqrk44jCNc3bZAYW+2OeXGfM4xJLb5yDn6zbqCGBNJVrkql9HTS5mvRh9tjA80s
pH/XP1jk+bRshbQbUyDuQ8l0bctbQo1+dKKjz2j9Q55f46qwrH3LLTbAdbH8tApRLofkvCaomzPl
C+o2ymhDvXqFT2fEtVjHQQwU6tGDKCVWx5RqJkhBSLzAof1Sn51qLXC1qZB/VfIe32Cr9j8pLS4a
snY6faqHKPn5F5asYVEZaoRNMPIA90+EMQDsKUCjncwOni1JuPZrloj8wikRI8PpVwGS1BgLXwVl
Xwf+nmxDaP5/Ra+X6vZZhpAopwfXCiUiyDB0+JTYLINv/B6wtCN4fbExkY1TDclPT8gONRfHK+nE
wQjhEVq/Z3RMK9BknVrXmud5hhFWEcEBDWz+hjWC4DuV+lv/h91tcAtcZ+WE5J54fCpUBq1qTFyV
tYumXyPAM40VXtrg19TbWxDWCX7B6/cpXbg1g4bmSGq2Ig8GSyNTJoXs0CNs2qW2nRC8Xj20OgU+
utZAQeHKuA4LQZQ5oKP2Hd7rDLgZUTNjNTy3s5Y4/HBjx9V1h90JjYT9tabEyl2kXf/R6NWJ+B2M
cqv93QjlbOVwE07MhYFBOMrEofd3yW2784RjXC/qqSekKp9l8yMkd62kIEbTQDqTNbr9n8+Z/ryj
1V6hxym1vdivl/zIiHx/M20wZ7aX2qK0rkEQyrWfp/7tT5Yluudh+AyaCj+P/A0Ou87PkgSeUmzZ
Z507srqXyPz4am6z1ZetO6Cnb5z26Rtvaj/R53eMQhj7yEtETDc4gJjDXB6yoQU4aKQ2WIIDN4tZ
f+4mR5S2vLOKJDssAPPqnOFA+rp8i147vJzPsynsV4kjiVWd5bpXF2bUUNuXTgS/c8p7k5Hh4TKd
j64l+GBBcp/QSeKU5nIGKLNYAEga58p/E2z2oyZ68A1svXr62WuGF05fKBJj8EBdUZiTpd+GCvUO
qgvJ8JBkM5wHwWqVRavRJwG8aXSAGlNyaTlI+/b7P82xRgO5BOVjzfZCNeCemDzY+Nzo9hnZtN8c
qsx6jW+Hx0dzpQYmyVMsIYptmzIUvFfNJKs9iririZDVra6zrBwM3Tmgqdvh1dPdoJK3gshrH+OD
QUOODYiDflwf31V840YgEQDMO2DzruggA0/8XliKWIcJs6df4twsNsggfe6Jn0wLOxpftozVzctw
mgfLyRX01yJsN+/HYe7RvnhT7t5CY7SVE4ZCniFdozONBKNy8aHoU6PmjsaNltUH4P7qcCp60Y93
QYRAsSLa+Vu4QWavyQLMh9Oq9wUwx2GVNhfTX7pxUgL52WH/UZ/hIJTkvxv7NfrZtgcDRyqqJ5ej
X1nsA1mPMBGC+AGfz1oAMNDHo8zYxaOR4GoKqxdgKDKZBxwJAzEYfQTnKH7ookN6Bbr/y0fNCT76
4rq9ZhhoEGCsbvRuRbz3SO7hjBkRX8pzXibZXi8jq/hi9kaP7+DPUPr7abibBn5x9npiw+ToBtor
gWoP2s1ldEOdwG+zpHjltz69wsX0Hh+DmHEkIYaOL7wnBuQLHLXhSPnzq7ZW5LdoadGpcEmOGc74
U2F+Gr68Zk0nAOfZZfhRQYvY1tTRgQb1q7xBms152b8bOo2aCxrRwI0uohQAStSFRJVRQG03zmEi
CziTUYox8OV7r8JCDOr2M2JscBsWDFuuBlvwDLrCu1vMqLD7q6F51ecs7eoDwnyNyUO4AYDCZqSp
RQ2E10TDVE4rvKQKXS6D7FFI0N+7k893zjGs2v+nyR48uLEmb+hxnNf6MVKxG6RtTYIQoWXQod7V
hZu/ROgQjMrKYD1hsjKlgYvEk096im9e+pjLKbCgdVneBu0MTBI7icX/43JremcISkoQheKZk3nT
kXS/iCTdETcfq6gviI32KHaOpNLtWKPNSODsXRw9zQv0QjwVPXby2/IXKC6ZV4ypviwFPx4GArSG
6GILyP6MrP6xHCAeL4lDNOdwrjGyQWMCyK0qaXGSz1ZhkQGjNoVl0AvGUbugQlc73kHufCXYfzLo
10onuzvHQDJtA+3xcP6Z66MURQTHhlZVmJdxu9HFZwzeHMTqDwqJxuZBesmYIoHAfo/ET5hb9ax9
k+9dmyJi+tJiEYZJ3g6pwpypvB4FKmqrE8RnAZFzj7huja6rm9slgDk0cW7+3SRl+Zh2m41gqeVa
/q+w6P8WcL2fK/TuOlkF9jw3rAGlA2l5eJz2om5tqmv6NDw7rb6Q0twhwsZHZQzjWnxPs5dqsidB
+EwnlMJ6URdBf2zwWwQpW+S1dCZr8mcT2DuVUQ84BNTxTh4qs+OyyN0VZ8zDVgqj2sO4Y8/uKiXH
rtUUFr2m2vb7ZJRL8CG8bLxo0jsL0l156OXu7PuNvPJpdkUlGqpRGVqmj3WglyTGNfDExPzMpfoB
9Uvt2HYTCWrDQ5/xIeH13WfQ73rAumuOQ3vLh4lVXxaH8+Q93uum3RIMhQmKFfICRxtbV3PqR8xQ
3kpsRNF3eIASQWXzWwILpvZGIkOc8Ep4O/RFisllckbnQFEOXxeAogpZI6fIe+nAS1AbZ0yu0IpT
LcmqfVYkETfEVf9yXrqbmzNW9DZrBrX8oaNwU0UlpkvfQqA9Ub7xpI4nzCEJgvHzFQ70pBmBccxX
5ddRxG04i/2c9mIzibBlIxcRWbJuNKvqg7L0MT5rmh1HNS34WSGxyxU4oDz2h+B5Bh+qhXQ5frBQ
BBFoAZjGr9SYSEhP4l9riGkmU3tHGAnMA8vd6b2KY22zVKyWmB8J5N0xZFAkBorTNhlflnTpri28
kQMa9oFWQvNl1+qYtyHUSA1NfZmr2HwcCVWvz5nN8gh6/Hp72Gi65TphLmE+4MepNgK6f9yFHTF5
IACn/kTy44aL/fWY62sf2tKXXs81p44BOYDzHYtAnBPBLJyQUNLxfKbPUuhL4HKA9TIN+E6lqptj
nHiQ47QXafGzGKsBVjeH3cqkn4Mc/8FavboFGiCnt+popLhRM/yeCs1LB1yizKW+OE4Lo2L3sGPi
Bt/fViIvuUE0rL1BccsL5h0ebMPLWgwQkmA6/DS+R+oQ/rmDPGJdLQ9w3EFeZdWOVCzmOaaJ7elo
v3+U5OObGylgmC7RcHHPd/RVFOe22RUvpNp5Jt3wBUvBrwkzILINmzdnRolLs/ULCAPFCtpPzQYl
7I8jqbsSA1Ai+OTuHq5WEOi87lODifd1hw+CS93mwbcgO2nkExLY6F8kVmY8sOMvoowbiGQ0mtH8
+Pkgi+yLUf3jAHIudO0/pcDPflUkltHZEtBmVCL9NKvpmwbz5NDnbP7Xmyjhtt95nyMPCzbsAyTY
M6JWRhlhtLZ5v8XODRJjzeNRX2DKhEioh8k0MeiLGhv/uQG6yqHuY/hvsagG0eV3rp2KZ582cI5x
yrgY1CjagdWegnBIdkgUhgOPG2++RX/iqNtCsXMGxmA90jaF6rk7e6QhcoZB/fJClKhcZW5sGd1j
3qWoSPMhZcYFVvX58o0Cl7Jpxoy2eAPLPobHeeR8hFCQZexalgxUSzce5YhBaT68Q1cSRJSMuSgq
0iOFAYVyp0ETfONQqM0IwGoyPyXZCu0XmKG42TzEuHhOw8YlRPUgCdhkE3mVMc6gV7W/yZ95Af3N
NLX1yKbzoImIuPuBJP6ZB68X+VgKqGka2l2No/PUxG0fLle45voHngHpEjDNXtZ54Qm9y54bNDU7
mWsJwwGCOsnVuS+xkF6Ghh/Xs75c23AZIBW4DyPXOBIWxhx8dnbkbRbDZ7zXPnuBD6ikdYL9nU5O
Z+lZ2f2WcDmtU46kFN508p8MdzeCeOxntYSapHO9e04k5DBs0c/kv1RF8Ky48Epq7nOuVcXlmMLb
w4RZ3oN4VTigKMXqFmiP2qmZMRr+NUA6qQE1f7p1RULWG1yPwxGjEwZ+9jO4fw1IARZL/SvwTF90
bb3OBOJlX8UQjlZ/4jxZczqB+JHnKe00N3R4heyklduLhnav5+uP6zIcC3N08I2WeZlLfNfQHPJB
KLP/iZl2HihYMhn/WwDuxEQEiwJExXmWbn09nOO1EB/tZFmONVa681CKQiNLLqj/ZHx/geaiBqOY
kzhuJqFqMp7mTc9Byungw40B94JsikLsY+roPhZ0b4Gegatlon2JuV6AeUEZOLSH3mx3chJd5jwo
EFHA0ugdBI/kMsuQZaO//s1P98liH+zAuFSZoiWIweUf6k+imLAILaUiDfe/hSl8REzo3sdpkMOR
ZyaAYQpSCKhVVHINOGYR4DmOqoRZlNH8Coar47V9neR6DZHyov+loUlfLDKk0vo8duD+qjvhNvut
JgfdfWbTXsggFW5h7/j6aCcVJCDTyYyvb2VoLGs1fYdkvjJesHP4+y8XsS9Cq/LOi90Q17Ub6gg7
5uFpLuy/8LppaA6rk+TZ5jgW5zNGfM8BZ3OQ86eI8D6QB29P4XZ4W8u0KtbAGmsimEN+7RM8x7hN
lFUvTlKUE4pMbWk3pavLDKfR6CyCg9latJnBhiVJL0NQ/V79yDiGO7O9jP4am6n/DmBGd84B2Rjh
Xm8NkNzYvK39N2mxDkXu6peWszuYcE7E6cXr/By8w5DgLIjMtGT6So1UO5hLJEk+m2CxSLftOlwe
gmgt5aiE7zeFVmJNSu6Ve/eRH0F7lNOGzojxa7hkpfbz9ng7efce9lFSw/3HUus63i2NxNzLdI+V
ZnKUr1UqYRIbyaEMB4jfUXQy9lVOFvxUO4kM3JAOwAIWsq+Kt3oCmuHs5smwoYSlobFcdQbhFlLi
IRhbqdxSR0acfx5xek7R6fQat09FFXUw+uLpIxgaLkydU4qNzh9+DLeltdGtsLiByruWqQAmGRM/
3f2zL76eyWgHGA+2+XucwDDJhXJ58v6KCI5r0T2ScV64UdJ8U5Euxmc1TOpnJ2xr9FHL1ZIZaYoZ
NEZT7m5QlAR3hM4jQvyzFjJz/NGKZsI4JZghi/2YGt9pyYyT4hWsazCIPiGcsncoseYezGx9A6XY
YlksgrdrFLaAqQ32yeZCS/ASeJiLXVfLfviA+LLnFYpLD4JiPonCgmTjTba/VLokptnjv/b3zvjd
OjcaAI0IWrfZg3crCAiZ34WfvodXKs7/uqXPMgPmGZbMT8C7UUZoMOHB/OnJ51ibWIS8WasUG4nj
0mCQeC38qNDtlak7Ch7HeyfqLLvaAEBg+qITjOMDUfxMf5QX5EQBLjG56umrmsJSlJ6Pe4KnmTsN
c2MujCVAmS+OtwMvUCEz/V7nm3xfplM+y5VrupeTNua640+6M4DRz5KFX2+28bxYD+jQO7iqskFH
uljIIYgQqwldafgYyKU0hBvEQ3I5QTKrS3pA9HCWRFoaKBKGh/I4q4Flppjt3e15J4sLU2pXfPFG
QgeKZeORCa4dJGGthxGdwqROqU+VQSCfzJPTrunczrTO93nDi22uZCJ5V/pI9/M1o3LDVMf0PiLi
heWCOW5py2ZrNMixwUDc5VjjYKfyeaWHFf7l+73nOeYK9s8RDzVXr3jjCb4G3y034IFDZfcNCp/n
ZILjNLbhTZJ3HQi52uliIfiufSffSsrA/5QDfzLXbo9DugLcIM/MPfrU+p1pKe72lcuNE3VeayK3
ReCEot0mrMPLOThJW5wGP8JuS+SkHU2gIYqCRvxIeo76YOjHqvHsJS//cGY0sIxQjby1Sh/xBwo8
alDeTxYxJdmOBx1lVx7MKN8YVGFPURkJgejX+apFc++VUHSLmxC6zaAQCPZwZaPFMwX6QlvzW00n
qllj7tzfbSLxKrcOmMNQsCEIJlBoyaSMSAnCtlV2nXvnLBpTeaqf7dbsw9OcLMZxP0iJ7UDbQQNQ
Y7l9HVXYn0RehzLhb66MX9Vim5G4a8ZZV2njYwO4T6IBZtHZx01J5nnM3GKBeC+Fh8kUo8qE7RF1
UmJxpFL4GE2PwSqqdXK0E1+AD5cx8oxbjA3EsI7+vGHfzs7mvWVe3sKdkh33BPeSQW4O4YsUdPfi
7xrxZBrQ1R8nt1LSZrHd5qZpfIqErxG/DlyZM8oxbLDNG41kpw+BZtedk1og/W+gplttRPl+IcNf
hrxf5/Ez0wcpizW+/sz9InahoBTXNgaWbwwSWzcG1CAxTO0HVFRXlOO8kkhs0FlyMhKpdVTMZkD6
Jz0IrW0Ns0PXbb7MK0UCP53I90Fbd2LbuLKX+DECravAitRzkvO1JgD8er3EKfeRfxd+GLN90SrO
RINegeL8VxaYxzAXJ7c9MytBgXIgoV07HaaFfjpTTERFK3TT3eYlb5iQzv4nFDyzrrKoEvErFSUR
BgA91YIgvWw9TRkqp0HpuwOeru6HQZLSzKqKKA7Q0s+aKP0kuxREZiveOhHEvekQqpzPyYHVstQy
WYc1Xz5hHj+o69+3/KEZdQQjttGw95hwh+yKjiQkGgzhbbZyAXyXeBXaeRbzSlVj2ap4ag1LNUK8
XNXZ1cdb7gDdf4l9YauUNGkVUYGkh/qd3brTPD57s7i6Z4miQy/TWznk4CKcZmNJ2s4pOgEGBM1r
r0elxDpguHV6yteT0zseLREXl3bjAs5IydOPvqD0c0Y+9VeXFwpmHEP989W9xzzVHM2eGaTGmlqg
gMI+A2dqqiYl6BJlApYnwhes+VTeOABPMUCKywsVU26SK7TFN4iDSz63wE8oIQXVIxbGd9Q/VYDZ
smI7zaln/oo3hUSFd7rUFAdpiFmhfR4k+iA098gP8lgv9SJ/jN6GVvoCpfwn3Hk3kZ4oEXCr/qg2
dMd3HeOmzf7fu0cm2VmBciCdtC9DhN9UfPehetaBJf3LQsf+x53onGsWIf/yKHyKTryssATczeWB
zKyldB5vw8QZc2SjVk6kuKd5j0BxTSXXiCLasqqDQa0CGnQPTKxnWlGhpM24PnZwxEYTMwCaz4gu
aYdhc+Z6Se9eeefVnnFMRhQyV6kvUgWX3D2RxDnwlT5o6Auj/c6jixhrWOOHTgtJuVDTNOShNYP3
4uTicUSUWPbxi8+CAw1JgFxCkMog/rqv5rLuk1Kqj7+b/AZ1qNbykm2Rdq6iSXyXFMATgewrkgSt
VW1Jdt/CIAMgs+WmcXgZH7NZvZrobbrES4imnvHX1Z21KM0Anaa2AA0NLdHrtu7YeaKr5tQ8krVE
XnVHUmXfkQOm82PSECVljER3NcF3EJiXIPTjKIO5iuXPpL7L+haTTMvtqgO/4CRDIXSI4AIrZ/+P
Zi+ckpGTxtpc2tof5LhrSI5l0wuvrW1f83lToygni8jxu6QmcpVBic0qOcRxP6aXQYcOJME0r0QX
KEqePaVWkGzxvpTzjBvj5X30NfAXPfxIFHD6d9dgvlmLBa9vCBeDhGmJamO1I08dhjnpFMakFCfK
DLlS+8s2n0H9MjiMckLk+WTqcVpetygTeupqX/viLmrjDkSVzCR+gjXm6eJ/71dfvB94ZS49A1ro
jk/C/N2rLaWtrRUMEPfDgOjb3e+KiI6fPIXiKMXIsooGbJITIC/qvnuIPhsdOrRRx/M7RY2TXq+A
DV0hcO19ul4mItzpN2KznLlUl0vZe2iQdeqlFaYfHx03BpceIQH+2z6f9osHcj9EVfPAx23TVDeN
XWuqtOQFk+Ui1GLnuDavAeMgXsEXKWvtRaWDCtxgK8025BtYWSkp4g91YLXCVkVePwn1nM6szoQ6
bDtxdl0ux1POsHZfQQYue0yiKMvw6nkB5x+ygsrxP8WoPPlDggE9TndiQhtioMM0Ta7kno5jIKpz
mIybPsB3+0Ba9JH0OM0f+S1xeGGeWJ3bgI8+tCs3KUPFFtoTjshLBWcoZAWnMt/uJ7m/RBCSJnNf
0u4mZlAHZYXWzqYd7sZiIWc1vZxG1nbtxMXb/KfDnZNZelz5Sc3Ga4e5SSBq88e2M+lw1eHSgctn
J1Q/3yt1PtQKTt1JL+n76rC7zQ8dF/RGaASUbXGz5chGpewhjmhN7hOJJRScqiMVSdqTz3J2GOoX
gKOkc90TyJuKrMcVxroo0x+pL2feoVVScbcoZayoV8ttmLKJi42106quEE/0/v0KS3w8s66Qbm8z
qjC+pNMMnAYHlqKesTU3nHIaj2jpHKuwsWaA1jeoJIsCCecISwytE6zrtrMsKCKFqgG230/mVQZb
4x0/Hcl6Gm6vL3FMjAC2dVejKKRlhc7M4pnjh1cYyWx1htW5WuDf74i+rnAiZncVsAXQO2pVxAqw
bbxPW+OQbcwBdUGE3uTuSRwCIga3ZmTbkqY2fcQFTGDLhuWDPH0ve6nncmGcyoPNzq1/bwNEcNAW
LaZmTQ8gmKm7Dm/UQNZEcyhtynLFgpFRQRLz1MKget8ymYW67YrXHwG5wWJDz1HxKKbplkIAMxEY
jPmguhUxGP9PvCj3TnfBoa6tEwECbRCoZ4ha2somwsMSJySCVbOzKfUInvQ0vCi4m+WPgzE1Z588
Ff8cdPPYwiXm36nHLnFLbDzq0op7nReJnsWAQTxXhfOLMInbkwi9SYAKLru0BiED0nHm5jAZ5csz
j2PuC8JtREDZlMhwJyfF9PGws+pn4xeBRig9qshB8nVt2w+QablyJ7J1zbePDPANJopZYlGuOdPs
T3MBbTVqtvHV37OV6QQAgfi+Zbc30nGmwL2sS0ZI/9T49lViOOStQ+oF/OR8zAeh9fN7UE+Extfp
5jn6nrHwqAmehTWfEZguUuFPeE+8spFTmaDbKCpzDh5VpQKG3KgvMuRO0wpoBlqihnwWLchhYVci
IxrfcGltNs/dm1HtagbeDbPkWuUn5k5ocOrZGL236K/QEgWK7qQ5glHolZtFZMtPn17vAzFWAQmn
FWJ81lM4eh8THD4yNca/q3ebTV2EZlzDgO01ulbqil+npXTw88Uf2yxZ/WY35UIuJaSjL/n0E+Nw
Lgujw4fxR+OE41qdCPb7/kaMn8PqXH+0lCnLnxWZeLtYrL2IsAMKVF/ievmR/+1TpQXEJNrlQ/4o
X14U27Qm1vOYGhy6faMiZoatTCP2a5Q73N96JsQHEskxzwSleUBzc0Zd9SR1gj0mmdY0B5wRIo1o
HfAY3d+hrGfgA59XOHfTdO+UI01r/TYbWlMe/8dOP2dtkELx/Gw7gGBpX6UWysp9aK1iVJF7NVyl
djdvfcfhfKJAZiSe2fAja9U6LhmpVezGURnF0PXfbCijnsbZ5l/7D+ze9dB6c1rs++1Mxw/zP/x5
pCXjQUxORVZyTaXqf8PTSCbybg02f0ShkaX31KGqJzfkiICoUprQtRsU4WWfEFQgyqeZRDJ/eejl
AkTCppaQDb9dPRaOIRxvVGQHTHuiNRi/6RHszjHqfL4n25KGRKyu4Oqi2D9ucKBEp7ilbVZsgP/e
7yN0kQE4ANtbRFw2THCCB6+NvvADQuDj+P9ot2H3d+YC+CEFCtRto+cvqDodS/d2gQosOnIJXOLg
kS7nS//k6ZMjUv8MfhMvawFj5eewE5R9RqmzH4MVyvAT71UYxbpFBZFFpguVoEnrg00qEfxdraJx
62b31mP7eU56LIjGrRsVaKJXVHKx2PrzUdpjyz7Q44XSY7KiNxHioyNvBEp1pb9CXDjXFRl/Y45K
q8sXxjcaZOlV+fJmG+1/cz0uc/rC3FnTPg/hbvAy+XI6WKn4v7f2HRY96o14ZWEnYJJUqwEkTUwf
GsUXNKzQvdPZIKTRvJ8oRQkdBOPy/nRfaZRhIveabMgn/s7sinRk2k1/agoow3Sc8h7qv6Kumufj
Vxy0hFgvwqwoLZsqMNNJHVh+nSh4cM2ilKkIn1tT1v/SYkaAhAsTFsJshgV7+DqY0fe+TUbIqsoK
XyF/hhWRNuCcIUGcLu9h1fr46key1gMvMTSusm5wAaMFRY7bXHkFsBPnKGsWVe9Mln4PKP4bTxpn
X46hWiZeHbLmbsPhW0/Qqe4Lcs7vL5/uMLrk11Qb4ADrk2sRbCX/ISescc8FFAiRUqdsWN+JP1+L
EoKLINTvd0G77Tr/Wpu0dqpC/gH3SkNVH0gjpatE/8XWaZsMhuj1Lz4cjcVGjkptYQjlmqLYmOeM
+EsBb4N2O+Pd0UrVzkEJGsbRr+/A1Sj2hho7zG17s6yjJGQEn/o7+F8KHEfBwzL+hDk18RPTrSyf
q1GYwToRFVJsb8Rh6o9Ri58r39ilSZGRoYRa4IRr5OlA1Ed21HO8Yu1niw2znd/z3dEvPKBJl6xc
z63Fgetmc0w2t7APYRrxPjAYwaUU6dDUFxhXmV7aPO3CxDsd3FIXL9lqeWEgGA03Z5bTcy7Hqez+
Ur3Aj8hF1Z5mEaQVxnXXwTweVxhu8TWAcymu1Na9YnaYKtUXJAOkL2+RWRjlp6EI0uB1OPmryM//
03QMFlweoQigZB8zz9TFodB9NlzkWkovm7eco27M0j9CaxON9eCwKL/0slEjOjBijJtrs3msi4aY
8LYQ+2hpNbFa6UFSayOB01EgbXtGstMSca06GwejHzZ0HE/o6GYk6a0Oee+Ox8vhpVZiYRruBybJ
t15depZt4ZMagALKJNyCl3TKcH2eUXoli6AKtZiUxwdxPYjeDjNOLlOtdFxzJjzhh5Mqj8yHYrn9
grF/K223xSG4oyZuP9Y/KgGO011k8csQcSvJNK0InvZyVmC6zjkTYe3wI5odUwxl8Cj9wK4eelyF
LALpydU6ItklKtjh/WZSUIbSH+5Jca2C5rTYjpjvQ6Voeo6Ik/i2G/xt+lJQRZ0dewHjAsT+tgf/
gFLalzW4SF+s3PSXMEOlH4o8VfMG2PVsbzkMYXfVJum0x0GqvoHB7ObE9nNeAFs7Wjjiuqghftg9
qvGZ3vVMD0pxQYae39sl9+DTGgckMCdHPscm7LvmKNoAuWUKfs6AIgNXC8AAjushOI0GTw1olyax
c3wKxUxansakMMRs94/yfp3H6mHmOKy1OEyfzWjAZ7lMzCaVe1yIuFqr01mqYN7TXP37kVUWdMTS
Jlm2ghu76FCMLSiUTVb21dbD+lHdf5RyYKpISoolOkkICQAkwnCmox8zdnRzRGuogFoILS1AlbNx
9npaRC3WHzVWtcCHpzdFIrN11M+er9p4IjirzvDM1ri2EeBRpO3Kft09bo8pHuBDj5tXxCEpKDhB
dYYWe+8UE4CWlBeroQuHTi+X2se07y6q30qySKDJdp0okZpn6oCsOBx2xZ8gAoRfaR+QHnRKSkO6
tfKFwLnhFlp1X9cc/ncDRuCsq2eYG9NfIDspMQKrRmFc2nFUS+dzghfLeZJW2nsv3CD3n/iaTtKQ
UAJI7WXkEY8xjvYpkoKjoA+uh6GeKCyHFqqUZq1SVUgvjjqdQX3qIYusL4rxVtdM9el5Mv10fPgL
iRpttAv4n1grUD/Uu7wYYODtBvrHBoa2nHUJJyen2PLSuyyNF/Sl+608JVNSb4C6NnJXRQxsDbpk
GUrBuT4y3XvtUt83gpnGTOqJ/iVOXGZw6Fb6aBEGeORawezPshRhK/2fZLtH3S/ZQ5FMtSq9hY8O
Sc3ZSHCpkqVJrNWlKQMMS2iTKWq71N/QnIi3h+km+v+TZtCWC7IHPtDg+J31M0EtwSw9/Q0MkUJl
/VmG/7RsRTo8kUDH9cYgcXqqrVpygJM/DYiXhvR9Lyw6RfCxAu2IlBMHqVgAIUOiTAIgkOurrUVR
PO1dgNUJNrZe8TsZeACiT0p0FLMSfs1rHcuVljazsRdhQOYmxnvp+RMre08LqBT1ajC2nhaQvhfQ
eb1BV+rsOQMkook7GphV3xbIQNAzSuxz7plrFtMQECZunrAKDkL/FYb8Tb8MVNwhCCeI/5mpHRrR
Li0fUnx0VHWEU20/FiFbN8Z13scp4sOWOoJN/pgvLVvMIqibHSEYc+EJMBbztWUiaI2yg8hNgkyI
RlJna9ajqxUwYRjVVfNM1W2E+DrxjQwFvyDlVqsPZvscQmTBaFC27wFZyKVrdR+gHJiRcDZXhXJS
HE/HTNeCuWecn2zrLyBGlQJmmcEoT4ZooR1gAQcs5fC99EokqN3NcYoBmB8SWrf/k6sQInz6L5Z1
cz/SZv0tL8MYTCCDH2HU9KiN5S9I4G2Bj9+da5EdCUho8xOugWyGHQ3bpd4bcEJa8SKb3wIugwAm
gC8B+Fr1C8LtV4SFcuUh+kOqmW/CVN6JPYqYNDCqDHu6cb7iFQYxuKMO0vddkRLQLIxzKhoGpIzF
JPi41NCToVCP+I8KcrmfLXJ281p78PZykF8c+FdDqre8m/NtJ2nKHGCJT62sWSszvRryykE5A0rS
WbGTJjPNvhi9Dq5K+EdKN5kAbHulinAoeTi6CPEaFuckJHWbD2+OsUTVTnl7Lcv2whJ1wkAb1ipG
1o4N/cNLe4qinnJO7QG+Zzx6LzjQsnw5RryWXMUBXeVPxDIJ/px1JAwAEQS/Iqotpjx1rlI0JwUH
fWME1uonkY2sUD85RW7qWNY1nRNoieQgGN2tWRy4U4fFdOFlf5TtS93iRy/AhRgp1Bs7iLIc0yHt
CS1g5qCRqSXL+c6/weQw8n4DW+uZ/nspXVUdt8coVyAJv7+hoCR0J7SFp7KzhizdvjaRBwCM1YI8
nxOscw5XErtk9MV6rNejFlhluquRJxaMnNZuRyL71QoTy9VaVhdkSGUY5YheulT21F9l8tWfzJ0V
MXY/BcfawNGDzJUr48AChuGJI/TUHoRt0jXBdncBaAOC07fhImOZJF2Jbq7E9v1jNU9rptl3LwQG
b1Bc2K2cqv7vEv4KUs2rb2UrROZ+TSp5BgsIucxbdV7ihY6IfA0/yoeSGA5Rlx212waz5kpe0P+J
P7E+ajtzGMo1DGpM2os1/Rc//J7MLKNfihYWfJP184Guct/ybLGWWvrHe1l2nTZ37bo1mrb8vBCh
tF4whQryrJwbSV7Ie+b2NvjSfUKxs2/CCZDnYuAGuVjMscWsO9hCzJE6jqsi1xRKlcoFchn7zafP
S11Dpsx73lnh1an7350fYGVdqAkHhrdVC4LDSn9f/WWdY+IS0/UYxNfv21eZxaw7gbXAxhI4qwuX
lCBEotwUMwYXCvHbSlNRzzuQu935gzSy77GhXKev8L18HRn/MG0a7sz8HbTdlpuWSTmkPn16hWas
hDv8hp1oyL+/Yqn/jUhg1xeXniPcISSYxnCVmsAXc1xskubdWPGs5ykTMpFo8paDDz8LszgtQgq7
4Qmj9adk1TMksRgndTmGrxOocJSKmQbTanHz5Pw25IA3iIQhhXpatwV49mf8zyQj5ywwt1JqjxhT
25UeVHcABLZk7VF0mJWdnRlv098r/HqRGeIfDdvGDNZ0trQV4BcqkhCdk79L2HD5jUeQTUl/IaYu
Egauh4EKjxV7aR+jl6pMepyP7Bs/UZzYRlpUNGSaolJ1HiKk+LeO/yyQ1aRJCJ7d8JNiaMZzsxwZ
qkg1r6yTZCT5tXSrjzxg6SNIQ6/6r88BWoUuKKfPif/R8If12XHDlQ7h/zbthLFL8K24Jj7S4epo
gDLvO2UnEbuhkMRFy3Lzp0Qm+EhoGwY+fLEidMMHKh8pF9Qd4Qn1szf0ZjHqmX4oUyUI1jrVY4De
XT1KhbClIBUWtX/F4BnbBK38/0RF7xpeUqwbxmFd2C3ngoWVT+HwnFcyRQzZ6tvLwGmQjSZsgMdG
YxtWBQRgQibqJHkJg4hMXL2YrV9lcgBx7vvnNCJNfbkJSXZY1sDNEAqP6lOwWkGPDQvbxS7pmBiD
w/DYdtHAUjJS/8LmqKnXMiIWES3rOahWtZ5jBGZfOKWbozW5GeImtA3ioMEUy4TItRP8q0qV31TU
F2MrK4FBQmOu0KTe9V+bbBNrX/3NlgiXnacRgPxN/CLZ8xL64tkkQ2RoU3FGG6lvVHzURykwPLSW
4VGPTF4GGtHFP4DOFL8XXjpdEoOGW3J1rZD+RQHaT5KimxZu8nUSaDLlkQUPyJV1RWyFmWtn06mj
bi85h0UdA62Fdq7nOxmKkaD3I9r9Ks5pGUGVNPjYs7nhnt/q9EnaWBboA3UuOa2uMFiCRas/aTNm
wDFO9VrgFq/5VRy4grrHXp0+9aj457ukI8oiokVfongUjuP35SOa0vkMRZ8YhT8iJKFFNSqsUtcF
5NS2fSpXgTiRX6jdiY5SjmN1A27rqxAOpakXAJRDiZ7EsxVKQ4wtk5xhFvAUZCMR5vNi7rFX2UU1
+4HBFvlDzI7yZ/6ceG4rdWe2zu2ZQBidkcCKt4A+PvxOQvJEfV6NREBgzuolndPB6ub0k3gNV6zd
5gmr0+pvYUI3AhZ48ryHQojX12z1roIwjDXV2wrqHHYFM6VCT5kvpgdVvHToh3ceI41QdtGRAgwP
UUzKftclctx2z4AM7QC0ei5OI23mFS5U8XuNFqCzb9QkPtgZpyrCPzIBx6wIbUHNZuX7T9YuMpzU
iKWd5j6L0u9kHIUfs8bk4bDURhwP2j8GZ1KeuaOJIxse4ocA1oqgd7/HkQ/Cnjl9Usi2vfyz2agL
plUTdjq3xQ9XxIeHf8d8nM21X7MtEXM++qayqdXEF93DKsd+gwGYsRkFnVlEm1t/ILXVD78XR/3v
x3VWpgA9OUGs7CEW1B6dBoONYogpuB1rly3rmSBMzXr7cnBzzBtxX6cDeeAkjBVzjk8O0+zRPCKm
oNw738m2IguMMnuXX40rPuie5LJZSBbgOjE3dV8VjDBgjDMczuuf3r0p242D6aEe0Gy96BmNiC4b
qCgd5ELpjjfxCbRdgwCQ5JzyQIyhKyeomPtOb+ux9LEMGS2e/1xcl0ZBghrauJNxratU/Ydc/Fhc
6r823h3jsiwCyja+wZnDgCRq2rJdg0PTtU+nSdUTeHyVG/w1ZLMWU0TLqXHqE0e8ooc6rVBj2FvA
t+MDX9uuBFectGzif1PxJq5E1PXj/GHgu9Lj5fUwz6lnJXvbQr3GSyO84mj7HVqO02uR/ZZPfnFn
zAhM3Ztl2xwOOcRtlV0v000YRlzPe95UXaw4b2aE0Gq8xpQzCgXxv1gmuxrwJUQTVaDNNG9Dpazc
eQZjbg8SgeXHZ0eZs1RNzhyIi0l5bV17SzrMXQRWd/JefTo/272ltGARARzUU+YcjGbSBur65n35
tBRiEG7uHw3jVLBaasaglD9g663KadyZ2hrXsPKAdgDbBgy2l+/CJkv/QdY8k0qKMTLofZZV8w7z
kzRhADt5cxR3IDjmWWmrKfxkKVD96nL8dWDMG8J3gtQrvbhyAZXhB34gG23IlQH4HeH22/Xv3HTj
2dIgmVkVle+oZ7v5ESTDNFaA8gnueCplDZhkanrFUd3MeRpkJgyBndbDOAn+O7kgzHsZiHAMLdLg
HACAFjkNovqApVQiYEFd+G8pNLGIoF+pP2CuArOxHN0n2KbJDcv7PchpEcTt0iE4JAuPRjaUBKkw
gPIv9BswcDlwXMQP3ba2uchcg36eGuqfhpe5V0BXUwKQu5XCtvQjMsWb8j8RrpWLD5pCZ3LYf0mP
CYJ2YxruJbXkMdUaa1B81klsBbSviuUIjb2Qkjpe65Vy2EGkJpIAWo8EuouN7XgBoqA7SgakYwSb
fvo3EcfxFddZqbpA369v8VD9LBa7OyLeco5UFGQWd1MM/K8wCLiASoXHQkZqaWxGgqNYxobvrJgk
/sHBSR3olXfHIsXFD4vTqCP5iwy0O08JXt4QumMsDsn0elWfpr3SLLPuWZPiZaUPCh1IAgRG/zTQ
Xl7wtgwmHimpf19nkpHpbcYTgST/AxjkwxjjodR2HRiBIBWHLYwjTFMcDKNN7tXMnxssmimohOH2
kHDkqNrPePVOL/NbBa97btLa4MwAdc1J6bzgCFEUebe1GN9wAdxL76A3O4XmwfTkoc1RgKGVCoEX
Ir8O2/seqDb534u5A2Q9LIcsLKhndmMug9hL27oxHOKtT06HIkkzklZGm3lQ+ykqB0YRIfzO5sTj
eE76/Vkg0vBpmip0AB/HQ+XBoVyU4+wibcDrY644klSMsWlk4mA784ckI8htkCrYK95g+ZLJMEfb
K8DsqQ27n8syzsHACDEqhuBJVT7L3B+lL4haks6tekXA0KodFWjFAENotjLdn0c8oOFZVWLXWK5v
yRKt/s9yImaVJw9Beu/UgQvOrOvCj5lwhz5cJH1KEre1BECbpLAF7qCgSt6Mq7vqrOv7Q4E/obNE
QuikoUOtdJjLbyC1HYDFOLs7MI2KJAjNsIN2bsI4P+pKVjYXxTY6yZlZtFq48PCWnIbNkXEuzttu
ZPE1UEF7m3Wb3HRAOuJU8W2FO0R8iRxlppeIg+B+TzgIOvfb7jlyuHlrQD31Cv68poA4kIrUJe4m
iZ7hPRLolfF7gaRUx8kiwlnNNMyHSLS9HV3Zd0fDJ5xKcaLR6LyyMr1R3p7zineGqTI51yMdqTEu
cMQgH/Dn4g8g9rPfjrQtHaxA/jSnxCd95KHme0sDUsUozWEdeQ3oafZ5PbhkVe+h5B8lyqXaQOIe
pNPS+fkNPUAl8/Uc/QqaK0aeDjpr19fpndGyNA0HAQwbWvAa9EFePnIk6xOZ8twei5uQwJSSkco/
q18LYwiwqHwCEdrcBM2p8mD7WgmeYYDF2fa37967fzrwrYzIrraIAcJniRJQ+C2q02KuR+nSoDfS
YypIplepltGwEuynd/IY+6Cc7N+8kwIsRvbeawuMDvYMresVW+Bl8CWwhNuXjejgMtcrI85WZbsn
uwUVNS+jaKzUzSGSVd+WIaBLesf0Jj4yeTJQ0ypEi7QYjOGCu4EkQEFu4Ew9JAv77E+mMhOvFUSE
1GWP/2TH4rrOvtZfnA91IpGguMy73XRd6x8fRvz3pqCxOXCAThB386fTEOQAlddjdj5jCBnSRJop
e8kJmEvGT742keXwr6nN/AYDZFlY8nutWDKjZK/wqx7CQbEey6zItu11V7xt+dJ77L2mlpKAWBQx
Fx4ExeyPz5ztDzo0nKYBFGs95RSp+kR5bZwwY+5FM2fiw+mMXU7ATd7cbIamNENRR0+4LBkifYJd
sFrdXegBhcDHrnekOPEmxJrh7BAdSn/+Rw+ok15XA1CjJjeQfeBW+TRhVOy5JnkoBHXuYNjmF7Gq
scr6ID0bt8523lpmURtGj5kb+VEH9PC7qd/cm6uOZcwSBS28U5vPcf/gqxVpYIAQg9fyjETCAWbk
61cWlyfNfhpvqOXXC2biiTlEB82+9k9xubcpbfp1xYjl5WNbrFRLQWOd0jqJpNQnD8UC+xVLtxoL
mu2NmeT3ACudCtSQFgEtcuko0UlKG2qw1DCnLzEULPtKFNMFMkIZfKWi1ofgJd4Mch913PYiwl3A
EdTtCn+6ua1Z7J806jZovl0eN9RLSniZoA8F4W4pEblsvLDKoarxdUE65ZEcB5iqH666GFU1PTZu
VmHplJeSEyaI4X4kAN3w5l1eYSV8JfwcWhx7sptIQkKM+Lw0BGDzC/Ax04WvzOv+JKTdBFro7Tix
z5ClHATiKdRSmXhaCqgk/UMWRaoy1EHFBcOfwPqcxj3RfyrPJJsD7kqum7+JiXA1gYzMTzKBSXDT
784dRmgipcq1JEN//RhDFt752Lguwj/GmoF0/j8zIp1GSAY8HKBoGOIRHw/3eyYw0CsYW2xQgCje
cpbhtXxPFjqaQ/375WpjIH/dafWhiEjmcnmTr/oAohDJ4mPHKAFqP+4h6uCFwd7/n6L91Vn4quKz
j44hSyq3KmeLAh0w82/I9I0V42VMaG9sWKQiXMvCE0MBMJPB8zzj0hBFaaTuJ9fpuVUzCojQ2PgD
VDeNBO1Q7QfGAlhXuAWQRWGtB3W5LIseZDnWutEefBxiETcAwI+IOaQl+AWk+HIyDHGaPEl7DlSR
seS1Tc4ydLxoy0+VdbhbV+tx1wbOm888ePl6UQIbgRf8CWbqwcXFQeXHjxU/84bFBrb0ugUca3i5
5ToOZlNgoxA314c/Z7WzZodPukNvrdqUADkfJzDF9xxJFapS14qLPJOCqBxOryop6lFh9UctTVu1
kQ5ChuEH6xx0kcofWmta4mhPg/SZyyrUwzah1fO//LNi5NM1zYg78eUq6Y7n9De3JAkMFihlUzPr
p5p/SBHp6YDRPJwjSgnqolDSvpPFVQQH/kD71l4VcBbGvSaX70cdUIugZQ9apouf+hG19bRUT4Ec
5XKRGmam5bGPA41qmVbpTIQM3HETpYly+8ixjXbHIZJdMwKbPAAAHQENqfI0ztd6W8W+9DcxG8jW
luX0bP94s240401UOt9BrFIWubKBlw/1snWAVy59YI28ABf9URztEgCQf1h8vteHwdi8R7GbPUxq
MeNRRNBE5UXUe7bVQsn9a3hP/eyb0nPm8lyAu5iwezg4Whs4OjVC0lipdjfywT3bcvIeH1s4kGj5
duact8zAWyNlrhavt+HIdbunV/3z/fhLZnf0Bjbinl1pm+ZFMmhLG6bNz0blMEk7HXLCYYPMDFww
OxEJnT6XFfC7ynrupXgf5vjOWk5FJ/h6iOfTCwoIeCBNvIIckKHsrDklxkw9kObAKcePYLy1OeDB
kGMpcpA8e/REnejTcfUmqUAJ+VWOYFYOYfKTW4r3yuAAdfj7m0vSwXV71WF6yfa6sR3AGxsxkzIG
U/4aHUhH0htrQFaviOBBBg4emGrRxgsVTgWpy/+mEPF7h/y0gEGaMB7CyECaupv8Xz+FKtdk8+/n
sAJ3Mwca4LmINGx3KNH2kG0HT+PhgzuKLGemywm+JkIrSKxFoBZ3guxUOOpws/Tz1mL0QyXFwqsH
6kEsoxvJ8G5DApaYXAcbQAGCJ9G+xcj4mPNMngd7kn4tzklsYszPOTGUUqB8SJ9/P09cKZmb0+KD
KgDyYTkda50mKdNDeqfCVo3e/12+AVWIr6qyPv7+NpGreQtiyTR/+ZRYD5csePR5JKXwvY9F0pWD
GD0ICmU0iXvGMPCRaFwQaVnNTJZpQafuLunyhmNgyj4aMTavBXsQiWKbjdLOokLCKvSZp2tRl8J7
sU/m0JJhKj1v7rY6uazCji7dt+WNsa9mM36S1pxY46nIgBQLrMNn5O+p1MB2HwcoPcyEsY1lUH5v
HxqBGSEg3BTGputm/p+ODf46LDgYGJAwyHELvb83cv5JdxiJ7c89QvH0l9/L5cV+SQzOGhPq8oIN
/REXetAw4mt3YRSI6zxIhoggU6cw/GBSmmeKKgbsE4ItArQTKQXl7bcOzTcSNER9SSRA2mgkLpvi
4g/WVTfo+fGFqFh2oONZa08HJq9ELbp5rJEukt9pRW4AHAkYrRffc4MPWb82tMy+468P6PnUBmh+
cIi2ppDSnZsnuD0hs1Ok0a1U9XYR/c9fa7X2yGb/lhCsB69O2+yLbBg98ftoRc3DYxshS0kxCFgC
ckYGCIh6GS0GR6QmJnmtYQqluj/bM7pADpd/AZ1nAlakQG5bTrAAasQ3y3IBiaWsjHad4XnqGNxG
Ha3M0st+3w8ItJqz3K9GvAVFbOA3s7hrUqTAU9KIDpfcrbm8vBcJjR5QIbbRQUxWWrATDLq0ISCe
1YBMSpottnh22CKiOk1/5uHP6JAeCvCgOJsba3u1oT9Gzsv2l7JPF/qJZpdZb6/6gIMkwtuZiksi
BWk6zFOO29FgpvKqt/S2uJzUrPf5+CEtu7ochNSdvX3uwap+J7GIFf3BjS2dL8gnPTplJdVop3oi
kFRg7jBrY94sqrUVpptFjYl7yN344ri0WjjaYCCv+PbnvVP42N9ZvSIpaNQZLrylAYPX8mlMMpUv
n1TrAIpBWXJGhwKbXsjs1fKZz7Cw364uAgZrWc66icptg2bwRXPPZ4EZ3J/IdqaQpGM1cqLdqrKO
qmQDWf+4tii1EMO4Wv0UTyYXXKhbBs9yi2Go6qy9WudlZqwRgcTBiLaw73FE6uEYuSrkWDHy4tKd
h9lgrJegwnUxuyJo0SWvX77ImLLWnN5hyHvVV3JkEp5ohxori1vabBnaXcqh8ksIH9fREG8Gybjd
pOXc52WGRnwFES0SvF9Y+zyJroUzq5ycgP0+G7bNt7sVRvFpdG5d+1jaq4u9O6gdZavUw2L0sUH+
19ToMT9IRIf7J3ZYL5d1VLoqny5b//4wh7xUlzUO75YNfzf8S9rj5xSEr66ofgI/ScPQDAeSeXuR
tBrwxIg5EYrXviP3/DGCVUAFOao8Rnri+XE6BD2anLprUkDGzf848ygf+yM+XlUT30zekszmusHQ
3XO5xr/R4t6c59GfkbJZgtmSfAz+9WkKJXnBgYjrEkj04VPX37QbO2kTVrW0qlXklExaoLCbe2vb
wNeQVcgLEh/RveppcNetKR6HyFVyRusk4A9kTOqBVuUc/4P3zp8/u5x75zWvjMCPMXor6QrD4TRG
feg7Qo6qHwpd6L1xPTzFVVuJtMnL/YqGpk+Ap9/1XT7gIxVJ5RTTmTatcdOQdbt2XtIf/ZAMTcAv
Qe1BSnMgf5yA0ild9YxkZigySR7FtwaY4jIzuFoi6N1hKAKCuMgjKjc8XZuAuzsmKtaZjcnEg2VE
wmGbklWAlVIgBWJO7xqMxofoRwYpHlqXxSdJmSH4niTNeA4R4+TEBJPlHbABTu0NNm0qIYMeF+WF
+ZTj5MZlsR7iIZfZuRx1DaPq2y0gi0fPJ2Rjvob3Qa5QuiIZnpvRHq8JVdsPDXwByZPCOsneUAKc
KF0QqHv6UqSiGnbVPUcpFSYNBpFJdtiSjyTmVQ4OZKLN7KoflDpCAVNuLm+xgodRtsIEjs9SEq+V
Vcz7B0ARpuNFW31IWh0uWXB5uM8GuiJside6Ucp6Wlp7NjxHVUgUJ0QZmUt2nfKVkx1fCZK2t5II
f+MAlh8KqmlDDFbNbyfDWEXBMeRMul9+LrwOya571vyoVFipBYZgHsnz7XSjIpBNCFQetr5myV83
F7IbkhqMzNgzg5hafRj/6bmqg4Ls4LuZgj7TuZjTzm5nKpmFMBkJSjIyqe+2b2VPWPwinG9L+9vG
0OMzwWkumhXoUJBjEZ1WY8Y2Po05471vf6jvYkLQ2o0K0Me+3jbwFYpuM1QTTvgZ4ThRYUeWaSK3
Mi7XSbYh9UwuTdaOuJr0Nn2ObTCmMWrgp4XuAgggL5GLFalwqygUejdyKrPy8hxmb1JsMe8EhwIR
pN8vOZIDMYYdqn0JnxPKOd2TONgZ/g6pRxfO6zvAxBu5a8YdE1/1slyI+EONncOrVSyjhQ/uOJxZ
xPuK3SxhaBJ3vEplv/M75c0OEupGwCTWejGB9vVe5VoYEcPQPbdquvGUVCXUYGGSaysk8nyspTMe
PilKheF6sKNbVysGf2ZnACS+0wvoRgo7QhWMYu2pexPsuzKYk9HSGuGbrV0PY+UwFLwvWgrqS7WH
xA9tBpq0lyZQFAhqkvQSweTG5FzMRxl220VeImUxQs1Gm7Jh2JA04SPiEYzXABSaa6ij1FvRFMdD
1EvV2znOvRFgJqMSbMESk6sKCb8btB5FX7WDGqDWVsLBFt03a2pFl+xlO1jlB4TXhxE5qWBZndgd
zp7KPPMwvXdz8RZ6smr50IRo6rd14XScHM61FQqZDSdO0np1pgGEtVBD0fIGPnAuOfY7ztnq3223
wKRWmaNzFKDsFq4rUOArT8KPDYmarnAs4oOYOXwOB+eNIyeQ9a2GB5XTzxeMFllRrjZmQ4kretRj
YPQbOo8DONZYPwmZKBRJ5zF4BhPaBcWIQlEIBKFEtj2aXXDGtZqGQV//SlHw6AVyT7K5x44mxFJu
PzaVylo+sXPItwDKUXspxCZyCBooSBWr3lEHzCbDpMhLM9oCJzmmqWA8G14ovtTpnefbd73FeL6s
wE2r438NexGUBjJELRbT7XbjGHggKfRvdF+1OZs7EPL55AEX3YYEPe4pNBV86tjr/rXb3nghqV/1
4dtuZWLUxmdkDYDvo/Pzy4LrMg3VyTxT2Iwr3Z4UK3KNxZbgZJmncjjqR+RapuMnZ4GLwoywLj1b
dkUFAL9UUsWUnqZZv/i6qd9T/k2lvRa2ppscNtaaPB94lMwBi8bo/FxiXIgiPy7wyEPahy4psGt1
VzzmayrzDkqOp5+LAZG0J/lyRSj4ZA1NAepE21q0wk9T86k155bzjqo9VGlvcN8KM78uG0lagg64
pHNP6+jKVtnsdLEAZqUSGc0cEX8Fhu4MkIh7Zdwt2vLzJSe+804y6TBefY0bUQTpMFWba1FmrJml
KPMKW1rtWSB0yF1ZnP/exAFpcguStQ5EByBIIPqz6jxnneam+iE66UMP+8VF+FXOVEbW7vPlOVyu
sDzP+MVz5bzGkjsrLz0Zw6rdl1c9Rwwr1hkXAX5u/WwNPsjZYbM4vX3z1raXPkROJTeHdKZG2t7K
H22fUVwTdzMPXHH4WMkqhjsQ7mlNKYex4S13UNL8JJwh7lj4Y8rCjgtM3414DuV/a28Y0P4ryl62
4x9/45br3OeZ5mtQPIK9ocf1As2uk7qRuYTXdsYgDet1v1yR2B6DwZbw3HOybWuKWWQ3NeH4hz4c
F8IBXvVSyUe7s9FFiDsNLqvoQxLFPlt5c//FRjtOww/J1Vf1T68Ko/nQINJIdtBZXOp290gDT7mI
OspOvIIkeFhntzS8gafDvN8OQcFuMmlzZxSdK0BtRTY5PNyG1VpGWX19wEb2AcB9igTRmH6ilKl1
VQHH3BaS06BfywUOeOoFlXhs7aDJJLgL7YHtlMMBI8CdmeUxRcMSeOanwYKhIKzf9hGMZt0a+0e6
YsWApNyE9QN8GPQiJ/O4bH+Q/sZjgVHigAHLuTHVY9kvwj85AsXOWSZjbFddM7X2x4LVaGWnhxiI
VMfUQxoXRVK3JhXwXGf+Y/7r6KBEXBW71BdnPORfzKHpFKTqEdxdiXEJy8SIfqQgYmF1y0qxu0k8
bxQeTIbpnqvTy8DqI7Mcn5caOkyzo61xOMc7J3Nb1S04nmJgPEBSJ1IeDZ9iplYMR4DhJVHNkH02
GqypSmgcLz/ja/dS3Jj69hKXKuocOhdtLdnkpsvLWE8poxLap8/P855nCKl4W/eKyF/j9YA3Ka6V
u8yt55FdM8mFJwaq++NUQTWPnvycmZUrCp3OYcUMoWHoWWHCXC3/rJSb5YiAJnQdiyC/KqO3MNfB
fO6fp1la+UG9dTXOLal3b2uKjAjU4Lit1WoMffv2+2uADzcHnFTPpRrvCEj7XJltnefEQMtRtFDD
Dzi470c3rhi7mMCWNHmuXoKiUpKG3/4COzrEB6DW/iI5lc9qUxTwWgQLK/Am/SmJK8klOIqp6Cva
TrYDF7HcXEb25PHHH0VshUEPlTZgDT28iRPxtxkrCmnpQkUCDXjikIHkujxE5O7GEKCEO52BVOPZ
6U4uvbHpN+ga9AqzxW2qDOe65tN574ylqxWaaKEiHQYKLZM+qiCPYo4gUVW5HZ+P9Hwm4X8Xxu7N
eE4y5ZJ2v7R074dnCV+76kUU4J8TyAzcDuvoQ6R9BBZFBGBGEW+XVXgHU3phuEtkDnJOwDkIUwpM
FJPOitz2yuiFYt4Pfcv+EPCsxg2ELZCZBre+sG7Zs5IG+S8afE6Hq2ivYqa3aCgifeE8aSr/FUaw
CAVw2kphgFd+OEzQs1a+o8QZdbgAkQYzvuxEMOQRyaEEXWq2zCVRIPuaZUiteso3+hjGKfIoVFJk
4Xmu4oNruDBYHiCSYylrDxKT/p/4DRkfGm7lEyAcNws9Fdupp2xA6bEu8nL1bB3ElK+DQuodsnqd
IiSp1ABASke7x0lnSEslCa5CezLtT+P9ZnA5XvTMw+Hl3HnNTOmco+9uUTOpJwfnDpPAihayXwTp
jIS+5xzxZOsTbckmBGVHMJbAlpsEsXipu0TDTIN983BneFIPGYa4kz49OJYT9nH+WjB28Ra5xF1d
FoLpteJGDf0gWpFp9O8zO25hhw98oRkzLKENWXdV72jGjGfF8McfO9gjUIO07ZXQKBfNk0kpE+mA
za7buXOML1vu5vgpEUlv3uW+8k+J0WKzSDrhk970EPxdMPAocrRzD/nNZkc+BudMnF16Kpgqs9aQ
GvdZTixjIBq9zju9u2kmeaYW2QKvJu/6FXDMzTK+6Bp2jAZBhvVEgPwGg9ujM/2nkNS0Gl7Iy1lf
bak0a539mf7Sgj6UMo6XgJWR75Sbowjw87cXIk4evIBsJKDROYNz0jo8E8Iil7r8OkbfIBUBwLUT
Je1mtWwE3j7kFqrh1Yyt7ksUmTj/DmIozjwfuWL8PiY2HvxjEqtWhEcdHnCldIfuIZDXPIgEsJ8E
BB0uLZzGidWeljMFkxDS5zoQMzi6HtWxM/xPABQBQk6FY28/hZO2obLz0GnGXQ7bK9RDbwSO/VcO
IoSVG3K+55wwUit0rOTP0y5j8gauKanPY57wTHXP3wjmlRxSzT24MpecdUQxGK7EwKrpRTRBoimh
mCt+NW2/AyWdTUKLB5jA74ahgS/DkjGdMMM4JKQRPx6TJF7wH6RGyVud3WGWJvBBYC2QmlXYkTNg
TJcKGcYyxgZ6Mt1taEQF5E7EAAE4pjfg6gIdyOdSsv1HtCQNbmhkUNmbEIfhXuPc2p36BRkdFWvE
a2zX/fb1o+9Tu+j20mhTvgjX9Ub4l/vrnEY2VV1g44X9s9bCNumVjQqTVkztjg0bGXM+Wnefqn5j
xx4xtwKuAA/n5YtQIqOnXicfueRwZQo4N4XILoTuNgOuWqbDZKS+HzDYxzRIC5AqIB915g3fLwPo
ZKuvPS61ES/jhJODts4vTHrF8jp9o6cy/jrdvsBVcSCkdCfInbPkcngRRD+Ga8aUKHZ837PxRQ7d
8WGELQMDNj79G0djv7a6s9g4M4vxtbq0gXTT9cBA5jbE2LUKU42fYM0l2pKi97oidGEMSdsgCh0W
zp6J5ZLIoICmkoinX0UNGxGXl61vsA0wDPE6AZuywx9GQ5v+Wa6dFIiyUHnUYbDtLJmkOFMcfdp1
LW84ee6usA0u715iMROxBtybjurI5uYl2CqtV6tzwD36rQxHRcgkk/k6Bf0a183qafe1HuVFCQX9
6EDXF62CoIceaYg20Kg1pT9F9/Bf5D391269R2T0C4HQqPIgjMGqjs5zvXJSDgj1SoUDTEtySpey
h3+MjqaIMFX0Px0FSLtOuBmyokS9jXoP4IdPQxt7Hu/6B47Ol4ceFZqeU98eai1PGAbfTA3EI3Zp
iuxU2T9KD1rlkV961/tU2XizgrHqqQclImdlJHgEtr++BhVGEdS2llVBw7dT2RDFOPBzjAIsB8ld
dtxt7ICBIBgSjeGYqVQX0lmDpXYjPv8uc+ZMkXTytwpAahjYKGwUc1abycPVsg34gKeoFHnHZuld
zXDL5Vsd3eJoBssZUk+ijnRmu2Vw90Gw+qBbaNArdQNWHgF+2BnOXzoUb+OomQ43lYG9NQFtEGf/
NWCzMJ2vsCPYlN6Upfw7VIwXv90qrGKVhzhq5/NTH47jj+GEHxp/AOmCE2MergAoPD3RS99yMhhL
XplNR6TqdNZIwbO5afqg4f2SkeJ/Aj9VMRSCGrOmmwXWUE9ouorO4G/WreAejO22xibcP7eOmKQP
ozTsFQO4Fjpxl0VJoOj8zhyWVYiWVnIhmOKI9uXL2wIIIhXCH3xM5r7hu5u9qXOCZHUJwmGIrZ7b
CUsm9rvZ+gWhlp6NBeAC/5A1KtUJSSBt2+uqBzL8anygW2YZFl4o1sk/yzL8du7OedkthI3eKT8d
mHOJyvtmheDTfhsr3u9HGDKg29KFTTLBXSze8mVxR3BliyJJhhvwxDtzLglXhE328ZW7R5UOgRWE
/B8OiJZr44PE8Aa0/NYLPeSvF9w034jm2VztDOPbiB/Jq784dFKI08OV1bFeKRO/5VwL7AmYE/Ci
3br8YXzsLvnIDj52Q+xL7+RFLNdarEj/9ZqeMkaXy+FrOUHxULIaIphNjKgxApsJCgMITs/h37Ko
Njn5JYrVPPf0tGx+NR6xPzBsukp4gbtSO+rjAaTjPA092RU3uGP7Dcj5I/jgIC00nFNcbD39spDi
P4In+32n9zTzNzWUWSFPGp91QSyquXA6dwAn/TNoIzTiE7+jPh1Fr/0VR3pBf1tnI88993Ygg6Sj
a1kir8TTz9slZmS0OUzt0wlL5GoU0nc/Orw4428nmfl1f+j2MbYQX5zcKyIX5eIPCwwqGa0bT40O
rJ7/Rm0NL3oZLETcBfAYmGxZrCl7EY/+1wEVasc+kzMNw35EhuI4InSaqwsBdeyRkJlfXjA8xCnu
voVAlJVBS4h62kZDFxy3YgyUhSZMpTCDeK4hx5fIkdfyzadu2powyw7uf2rdvsh5Ggt5hpbUsYau
rKFQyK2qSiMwYJLWhg0zNupNZHIweUyE7b2ncl+B5BCmkGNKWsELq2wAKE59x7wHk/9qNf61Kc+Z
zlgM4qwLvRpgiJNPZWrnX6kvBJOSEcLSWazhrgLBLyK0eOUYUoheL1L6IQ02SCJG1nIytG0NvKJx
1TVVDt9J6gymmvk6qUbQAgC8PG+2aDSUOC/+tkrhnGDNiDphB3gsCf1GCgJWrOsyAlE7VZ5sk22J
/GSIseVCWvcwZUcNzhWN9hU4BzV80OZjFIpBjfqTjo3vghskOQy7YRwwrPQSHbmlnElezbkmU08R
Kfn8BbymPXCE+nKdxd19IKZtk4LYgwealSVwaGNiDgH2QJ1pWcCCs6ZPmxNaK790+18pvTMWz5s6
59Ps6RhFUmkgtCKvs9nQB1C8Lv39sAsQhofjSyR9Vc3R+MOo0g+0gK7ZL4DxxmoBfbnYszgVOjQN
K9mJr+T7Jd6/9fPSs+xabscf4ef3UlPgavsnUqOB7GL03qwuGEP2B93une7SvJVE3cEUfjPmE57G
qcABQrEyOtM69XB4l70vvJsQtjA+FO9nvlczSi+EEf40bWF1HQacjhTvkjhjyOaN6FDuLnS5/ZEJ
l/lmFsIHqHqh3PAXhc7++n1R5RvZLMPKRt0tv1Au0Q0xxusCgm0aDVdd2GZQtWCm2kuzSW57aWkT
XhQ5zF5ONAzvqOzrzZrXz9+3ScdsF6AS9cJz+aYq0WOZFxLP0FXfLoFPPqXy2hhJi6fERq6+GZUL
HfgTMGHBIytpjZ/BIs/gklno7vvsL/p68ZsL6+UepO/iONi5I+W78BdQ0dlN40uux0xNmINqGQeJ
QoKl6WVF6YPCPOCf5FkXy8pZnu77FY6WJnGLim13djw7DGWb4XtPPgb9RClOTDf+V2WZCrNJoRdW
UYRElGPLYxBP2DWnerq9TpXPc2y+hodm0m7urGKuM942Tk34M6kHBAYj3zmio3Dl8zburAu5D6Bo
Qo18FUftdj/7THqZQPv2hEU0y8rt4k6V/TvC/nzJKyTKdmHsQ6x+5geET3N6QaSk8oXO92Fw3kuN
Tq51ygTg4nye5mkUpu+6VYAygmvwALVn9U1gacZ7pBFxyHnvAEfqJTqJFv52O0uj53qnPZ2h/WDY
NbwyZw2yDMc/xLU3KzeAaKr2l9bKd3xe65Fo1vmnDJdeuRY0rIkURwBYsp4bI8sOSFNr9nxgIkCp
TZA8ZSVBTMb8zHuMpzPqD6oKdJYr5zLGkSTitIPt/WNnXdzh1nVjRFjwHvaLhQT6gQ+DEm4aCwoG
J6s8Tdc1+j2YOJy5rWKMqI7X/hJL/8Tks5idUcWZEE23XvC56/N/OrJ+EGQayfQXIuJsKcwjcgxY
OZEfFJrg4I2mflcCNfvLoLCYkm6O8P2Jili8oMIn8xQleAGpVgiSfKab03QNWLpBZLC41yUV+xeE
e312yvilXh4N0NgNQ5rTUFhA1GemHpa7weIXWSapgW3YASAaR1/X8MEmn0qTe165wyQbVaOq56xP
xhQvpQNUKz4Hx49aJiID3p2hv/51ujWl3XWryMf49s0F7nK4u49vbTzRjEsqUbeCCx2EECjfAjwR
pc4p6MYVwMbtztMVDKtiya8h/sKDp2Gkoy95H/0GrymihT7rDFPZVphcDDh8N1dqJ1hayeoYHpax
zhtm3a48oGVsiwoBAbnZRomBErvzbtwi/IIvwZT/Dp08i6d/Be2lzufCRyx9NmI6mZh0y8cC3mop
wnGOvAwa6o0YmMbOJmBBBeVC2acrJDRhz0og3UGNgJCXaiN+t7G946I6lmboPbUc4/jb9h0ju8Nx
PsgrNk46RiorHsv6rrd2bqH/BJRBDmxP2Oi+wlC9cFTSiCCy+N9aoSOku6FYKrziq4IisPC38RPL
DVpqd+2uV9loGvnCX/kEecWrxbRUMIDZXJL3Z6ZIlvsdgMRwrHqQ/aHYnjaFAs0kk1EkQCbmhVf5
iGlhHXxEMM++ve+TeD9uinn7uJXgvxAc+3BBLpD8tJKPBl7yfIEPDctGiEroH+BwIPSAz1ig0zx6
mqo7kzEQSTSZOfSsUYlKdD+4gjhBIaJCXB3NFsy2zDx1/Q62miNwqmRMD7y54/nfnWX4NAP8YYkJ
PV5oeizlPHYENC1ZGV+irbK8UwWsjzSY/3P1gmjSIVoDx9bTOLpO3qHRt/VyLHAbwviodzbxgxcm
g34gnNkIyFjlKJUh8NAqaKhcwiPc3jWWlY1GxoCJkSi6djyY38Lqq1mClVY2i+9v0tJyK7/5m2Bu
fZUSJ+/JXCdgtA+H2AHCTEs+CzxjfZl65kA+YlrUYz5SYWwYXOfo1A+pERkdPg8wMltA1M8lZRFC
cztJ3UfST5hS70h9vvTGndS9m1oJ3qXR5zrbE0n4Ep2724gnW+CHZAazVJ0E1dQZkdx9KZ3fOXAm
BnYjiKwAtLhqZpg9Yxsa4bAfmpQq8chPDU3YFiFVrQh1FGkR7lcsz9aFTxuU40LSelAhFKxBg19H
n1mNOatmXvcIF68ro2hNkgm+5CF0gPPR20sbwDrQ6xARNklULScxuDy3MJ9ueFjDmWOUeKL1fFRd
0o0W0FrlV8w9qIzC5tSRft/l0vtlC1rkU465kqzHiRDPEzmch75tzTTnwdyIBFrafTOL26wNhctt
OIDd0III5QZ66tHJpMWQCjn3L6wpfHZp/EsAMJpFpZk9ynryvJfmmUrSjqI/mwMxhavLhKfRmKOb
IM8FeIM1Nre2Vunow+Xm01HTEOPRwIoqtZfnSR4kmd0qkhJAkjiQzskxPq9OQVHin9P2MbcV5SPv
zNqKSKVjxCe6RkRKSpSiFkyRBapmPWuqLPuhpwKcffHjxqLrKNbVDmmcU/aABznfZ2nBELYvUmZG
5mwbDs52/MFwlCuRT05hFZ673OzAJ3l7Z8r6rOYBhRCTxfCakW+nDLhIhpaL20uWOvtFgTJRS2md
TnuhTUXwS7Glp2jcnJofyt8sMCwCm6mQaji5dqyrOogXx+y762y1DdnKQEiZIfhi8aOMchAIC/g/
3DjlYKcrEr1F5KjunT59MWq1n2WdpNP3gHM2viPJEkWqu7rtbnhtnHjPu1a8cNM3mb8m+mqcdgQ0
UApNBDr/zPJsSB3s9bIVVaweUyEme0LzNZEdC/mO+nDKpJ5U3Y7uRKeTaovP1wg/a2PuVCZ2J0P/
kMd34FwVhgK55AE56zA26AYFbVCpey2LyUSXsMjhQrC7dz0lrF2gvKeEUp+wZUb3g4xANkMWtTQa
Af4dBCXTJ9EvZrMPFk8/Tl68B/mH+E+AQkAqg/PA/0p7fJL1nxCN9+c0cjvOHJZRkNxEx+Lk25HZ
fjWbXQfpdqhDvAA6kVITcOytLnL8+zARwoI1TwCpw47Cr4agNJQu6B8+oq6cLlnAa1xVKYAsjkFZ
PZdpbcRFeqZ+Cj8EaRVoX0W1h6JMT8Ulv9X9et0UwQdRdxggVpo2j40cWhV5iV/fwPYkfz3NXWZa
ggT01o2uKkCMKEEo59f0oWfvrYs4lbyOsSOdxQPb1RROCV7saDJbl5b+a+hOBduEyBgVz0vnUDf9
cP3WwMWxNCOnc6iozmab6QojVIbepeeWtrdNt0pVGTlco1E/jjwjZjBe53ldHbvLg8NKqMHKjuos
vExNO1MIx7cCLMZqA/itnjaI4B2URqVgt0KzE/F/okMGusodcNQBhhIdSWQijkNmzmuQJ+sijkod
6fQXSCZmi/EK24+GVcNARmgarFhxpe1uhy+/NxVqg/gxmlod8Uv6LcxFZWUFb2zLxXGmoFd5QGEb
njXy7LhKhlEvyzQAg+wSn6aRwiNm29hw35QOAwcZA599E6OzBNYvG94FIZqubZzGu4VQ3QksyuOE
fN9fonp3EW3H06q2nImchgmfU3l+23yIc62JlF1dInhXm/em5iIz1aQIVH6kVeWyRPs5o8pWH6DJ
0qHUMPvYGQFVt11/uhkUBnRZ+i7OBj5PDhtpKUmvbM/zTX78kzECrROUhi1DC3MDQize4rv3/w7/
VbrlEm+0xb3Y/QN+MZD14FhxVn3DVCA6I/QDuzs0nl49qOKf9jTfV3wHaOTNAuabT0cMQL/bb7MJ
bwXpEOQho+eBi7qPalVxiwVnWmYfpeuM5dd9pskPahjP/fQN7aITY6ctjbYWONf1m0tRNm/DzaEn
gVLS1l3M4PMCWdmP0zN0pwDFn1BKhFN8gEWV9FMlsgRG0GMjl4/0kUX2gUB+dGKUARbF8fN7Xh2Y
V4X/JwXaUdkrQRTlAKbIIVVsnqTCmyy0J4Zb+I3vwhME8UGS+GITEjhcUTiHZ/z8EdjZLFk9SqVn
thTWzQcMRatlJSDEEkHEhLG7OgcQfeFIKRtq9NsX2hMsZF0ua6s+bPHTRFi+eYVKOVP7xuV2SNyx
cV6DfVYv9o0Vku5gEjaSUxlRuSv2XLCDYx6lt4PJRfhGNvcAmwviGZ3yMVJ4H4A8xpsbdB+rINIL
EO2NTkEOwg1E9bZvVin+XB9dfZA9WWqNpBsHI0KXA4QsdoCuX/a4xGv83QutbJVjlvGTlb5atqFp
ymynIlZJdHl069+Tp6jaMt6HKE+l2jDa4LHX2ppGwQmeHraifaSBKY5iYNLEUR59zMYdvvhhm6qy
Fcfk88ILSajBgeFd4R9sFKTUO0OAIW8HrecCotum0DzMCkygFBmZmo2y4qWGgYoNeCuN35ImGAdI
bECiJhDEi8DQSlutbjisa/OsdgJvHwvgLlP2yRG5P0mZSbLm/YgwJ/zx+3YCsgJaTY+Fa6MsOazi
sTlot5sCgWTKWlC/gkiSU8pN1HglbTfbaqdfZ/2Frd+FYgRiVYDqJGECGrJN3TiFFrWwsbASF02u
WmuUFpffLFQJGa9GhoAVbiH14Aam6ej27clqN3EeJecF+DniaAauauOMQUDubLcTmWAPqwaZS2T2
saBYy6ts9Lra9lp+PRqU3ZVK8SlvNZMpLOlobmiqDCsneN/oiwvKds7AMIqBRGK5LkSA3EZBtx1b
ZNwYEXiWAYuBLd6vHLLOCRbzrvSHAe3FvOBnHyoYyIjiqq6spANVASVoQaYctkt7xPbiB2l9w53o
+voxUZkYZc/GWt4arfbBFgmOkvzSAlE9w4r0hx9RX4MiQGUfh/hMellVA0CToCW6gSSqchaxae2S
qsa1hHyb33AIZkLj1qVZuopfYNU7n5WrQAuQME+3ec8J4bgtQmEBQn9ebMGxFdICuOT5Fqtha0JZ
4LJPq6B/AX4rCm4okddmgt25p9Mqo6InJXdvo164gY6bYyJD+2om4n2RS1QWFmkjAiUhpoqV+kHe
WhwqiU8KQpDm4WTJfiH40+wevQL8tcnX+ZJpNF+SbZ+pl3scneDBrDJyLnESsI7Zyc6vYDvMqQai
TefEdtnCjd8pPjhuNB5PBXF/L7Ceb6FJ2Ka/TNCAjBD7h7kP2fShm7zZDyv1i1rp1grf0rmPAWBQ
YaKDKGcv69bzQwZ4FSH4n/ASZKUPj4Q0FgkvFJHK9xwkspc79G+qXppxeLqPAJzm5YTqwunoxwOV
k016VLzfeIYEEimTFTL85vxNJevi2M8kjRW5wKQ/7UbpZw19V91Dpl7M5/3qywH3kZwNHaLG9FaK
9tJUjmETfvtXBW8yhl/m3XgrQum8SsAoMB24rtnZ2WR0JlVnrjylqsVgQcowUebw+6FDFuMvWfpT
yTfIxrICZAdCA7qpCOyIBQrJlx0BuMs68dDoMFQ8eMPv9bx595B4XYaNvwfTG+9ovovYik708lxa
P1AQI7A0YkEwmJO7V+F2ErmGb8x+6bdng7/8oPU039pmsgL8rLOISAZHDOpNF7L1ubhORYmgUlIp
IJOFo8I2isj7VlXZZU88b4go2/wn+re/yzXJf9/H9XmQtps3TLjBxJyE5FFVGRXZVX57M38gyJi6
b5lJQJHKEG6Yy397yIDn//RtydRRU8BiPitZocgt4DEeqbsLYJQ5NnvWOUwxNA3j3qloTewUXfLK
Y/PJ2LeHR6Gy10WEERZE4GkaIHSG9UgudSIFS6FbQIb9xFJ7fZpCSHKxojNisFcb03N9ceJUCnyN
QbykR1AY98ZT3lgfk2pJbnOX71P9bPAgJ1ghOTBudiZV4awqTqUhkRiamOfsqZKGctqrkZfwiOQ7
2cKoO0NJB9i3EwIML6hXbChZDB2rplBXjzNvSDLHAw/h9mTfDQ3epmHd8Lrn8Zt+AjJCdQHhoxQT
127hMcJXw3CUmO/xn8tV70QPsKmmb8P+mKSRkSZvTXGrEfF92jwl6iy8+0DPRVJBNwdQHjDz1wzp
Zdl4+v7TeJQ9XDVQyj5zesNvYHqJweDsXo2QSd/7QMpdCqMIPUrj+9Z9oMysNF2p7HoTtJX46kEP
bQ6DtUdyYLnzxTHdMcdysadIOc509turacdNduBKsIicp0KMc1ZeqCaYSbjXqtS+pKwFNaw22XPw
jUZqLhxUOFilYDR6chKWLx/ju/Yj0SfN+C2zcPnMwD14mQTg3fNzC+MKQkbcZ43aI1urMBK5qR/l
BG58wQz/NWMju2WE/97Y9RkGYRyeFhDsXPU771SwoCjMDkF6NhA3MrsBpdO35UPM8XAE9vjcTon8
46uZNJ5QRIFsgwoXIcYzUHj7xSu5oa3/SRnOWT9rdkp5FrSJy1tMaix+26Gf2/rjULynQ4VJqCRZ
i81JWXePMxU1IsiZ0th15qxs9jyn3M43UQYCIkvhS5BSnrkZH+5szUzBwsNqTpjKlyupt0ey7LKm
sXgX2XS3rdzGzAb/ETW+Ai+Ppi402V/J3ND6f2IeKTR3z3h12AMJi9YNZ1Q7GWtSqEqJTD1nTSEI
Z2y1COwi0o7CLxetkKCGX/cRKfGXXbk7dDN2mgZfwu6XGgDiElWuEZjQKJv51UPLTqR5NT6BaT8F
UsV+3HiSNO23xAm0nmiewiJXlG8boCrgM0Q7Pt/pfhFBlrijjd6wY+1jfSvz49vtGwoo5LBVF+f0
RJoOjiY56VHabygJcMVwPj6R5DDlrSVqNL7O5YLbddipVPwWvby9sGrzF2+m5yZf2lfrVaNutzT0
1GepTDXBZJoKSfQzcoEmZ5Ba0kmQKeFXilfRjlcXn59VmAFnR/BlyFn44iIsc8+8N+iN/tw+WSx2
yDSiIwpCBH3fmYTCHJwNKSp00dhVFoBH8/07M4fybTYLHljLBxTEWasIvPIw95I83uFozFHDDdA5
mtiCeD7Z0hsUZl9SV+EAhFHObYFYEKtYFJhopBOMIrOC+v8O2NNdB2NzNmbPPsP/0wP8JGI6zUC3
OpWOtWgUuU/kRu9/EOhMaw/OJCh6scB54HNUQ6Ir9M6sys/vXgDie7F1mqtz2uMLr2iAP8VAJ6bd
3831Hcz4AiPc+0mzUDl1CeBIc1cCxLgolp3wnBLLCCRTvKyQ5vQOo4BKJevaI5YUpcaKIFXGKpZF
9+FerGi1r7ht6hVaqx/c8SIU5X7dfUJiohVfPxnO+48TmG1mcM19eokhXXbqw0vaGQ1c3goN+iK+
/Hom0PW9/OqqKJi5iqWBalRV6M4C9YDjYkR1jAqEX6WpoFa/xy7pwQdKJzmC/AvXWwnNLmbDaMdp
1wuypn6aDigWOVyi7YU2ikUOvjkfndzf9jbNl2rdX0jAMl38RlwKowe4P9zJoJB4UcrecyqIxfY1
rdI2lu6tbBR2BBlxVzl8D9tVKlnZUrFe9oEKrxpoEf06VIJrGBLbxIHcfEsPx9oYhzcAl0Z3WaPm
RnDrJk0d5nxcPX8jEAZrJ/9GRdzk2Ez0kzHzGeGjtuSNYMvO8bEPCLnHjlz739+XSTt99GWA/vYu
Rm6P/kQCHrY4iqT+ZbWyaxmEELUCTy4EfyTRjcgFNS1a9OEgxfM978bcTPX8SQEf2HQqbgCYykFh
5jmFRbP+BAWNOcuf60Ti1V0I7hWTla9ba7idIYbuqy6H1qcJ2nwZ8noDnFPmIO37mXi0nNz2mYHy
m4fUQ3NRXJAHhEczKOUQAkOjxrMkdttIsSDW1IrxgVXEBxOJAm0gdhsKusQuqLub1RfNK/VOMb/U
dhYrHMuHjJd0v6ixPvezZvv3ibTTZhcS6rPMpeWLgikI24xo3jJ3q2IXaIQhYihJFZf/ivqVvms9
BWkH34GorMo5j7d0Xa5yV4t4ZE+RwiFGPqXeV4LNSwkhRkBs6uido9kOiLvcGK6970d19pwCZ3ar
B5ePPLSgGWOwkKSFCsn/LJMjE74QnlxOMq4yCwfr8RtY8aUl8YoWzAy9XRTKiTIWL5kVeeYwxXr3
Myovz7kwhakoTKDeLQVtUPD5AK1YVHtho6koaeuTjPmxAPVRboDp60FUV++FTHvlW08B9gIXoj0R
0tfbK6YHCIQb8alqaS0jBJPPXN1A35Jy9zgz7/hOabgj9ZHt50gS/3LlGv+Uy+xykhVLImEQ2zAr
bas2cEkhSdG0qaYIiOZ9PjZ9Gzto1jQURjRGQjZOJAXyjU2gwKs842pEFgUf2JOCC1JjRo3PIBIU
g0LQd0Gwx7WLnI2UCABxZvc7Mdjaz+TAvjMDjatHtrK/zoCSYf9pelB7QXTX3jyG98jtwjhkb7PB
YcrKwUhGdQj3HMBxVSJacS52lMdc77OwY4CBGc/y5jrrd/rw26eb+ySvNXo7PtqBtccbSH4fmWtT
2H/li3kqxlZ871srZFLmZvfzcLkZV+oJJQmAsiDccRu/oGmrWcVwVe4LyTFKT/MgdZKyu4eGLPNH
S/TdRn/cgZbUmSDVpTu/rH00EViaK2vTMK1cf3f4f1rOjd/5Em6oKTP6001xeUEuCEed9CukFuqk
1huIwEYbV63E41IBh4MO4dV23koQn0y6ZJvWGYBUn1tsWAGpMddq9YfT2nkV6N1FMJct160aor/Q
5Ib2wYtAB14aznlRKIF05RZ0t1WnhP4xK+xaf/rCooBO9aUY21r2gwiAaNv/63eNNVyI7Rfm/tkB
yCEnIvjJwdxyGUL2XiVIB4+c+IritRnzkIC4QG1L9e6/9jhNLo8bNCwooAYOkBa++jVs5Khd7wfg
C1kHZWZqmXNArPYUpleEyp2lNsff5gJC1ZSTO0buCb6FRfXYfp+0dl0xEwvrK2Ss+y2zVFj/05vH
xdjGOEMVVKGkNw/vj6EJNJj20hvJLc7Op8XkRFrxKfsRQZwifIQOs0oCCvecQZjDz5sNPjctAfB/
hLi/h0UszTe2xnRBFNsuAQI1lV6NxincUi6Jn/9Y+wmo3SKFxgTVUdGxZBF7hId0Ml1oGSeS4HWI
1Mv2wkjjXbWOqKv3Z76bW5DrJdj1b609x9zJwuWXsOZTxi/nrxUcg+vVQmbnTdda8vFQlyt8Bh7U
YJG2KEiCij8uh1XU/Wy9RIAJWV1NRwHVjvz7gx44r6Q2P8DIkZ3O9kyoMokXV9PEDe3Msiro6rLM
XciaV+tXprOO41VrRP4lrFVSjr4tKgmIdoR+8f65j2+Gb8KRyl/cBZbjpmlknxWLAPGQW/aJJeAH
qLJJE7tDx04PJswCqtKM+fGANXbRi563CtZlzw7Zt1wBqIxbJ03yf+JuO9GfsjVmHTjEafxW71W9
d8W9AxsDItT+O8yVDW9vVarXAmhohtvTAwWbISU2qr4ONub/NrzYI2L+LhA2XdvfaPwRYrKd+jZa
SraWyK6ggKBwFBUHlTg89ORSM8/AQG6QnFWctWFiENmTwciaHPdl2dgWx5AGVfOv2xaQt1gMx4hK
t2FgtRvOXOD6RU0SMqohdNjip0Kx7EpNilhQOp6qeeXm39+ctvnzfZIRt6kybTjdKKrYTl4EwfwR
ZjsFlp4ymsKf6yPLBg8OnjirAUKhqMflTOGUl632omZrhFWmQPQe34hkgaEhbLfYC+TJYFyu4wYw
953pmLmWCrDTlEXXXFm5BmRUDSY+yc3++J7OiJlfXwaeYrGNNir7NFMHBjcK5tBpMTnzjlybYFnc
6mLezTGTHPTDd5IPb9mLh3p9JZIsMUDBMVKPhpsedq1BjyVqBozrZqstLCnG8kC4wNJxjqCD4UA/
sZIpOforZEXlOKhP84YLgQkiTjr9SOx1QWKt/yLl7R/ezAaAf2h2cYdAGe0T3G9MOG9kQFQZ7M2X
UGK6FvDIOHUyty3oHXm2RyU2s60IKuboJskrjq2C8uaW35MxSsML6IWvJicKl9Gp87x8PVcHm8xH
CnT/9NX8eoK8gj+x2LVjRQwsiPgkajefVTBs7gIsHzT/Or8Y8u2tNDphwMpY/IfkIJuPyFqMXyjU
74H408AaCaxT1Sw6JPq31tFboy12GgLeyBuyN2R/4ihVDsje2+RJs//Oz/geqAJJ64eddHvryBoX
2N5vk909WcY4nwyXPk/ejRMQWQPrpgOBiBOKo2acGsjMay4HQK9ACJJHs+hhv7cwDuIPa/5oLMxy
At29EAEOzN5XDvh5nlQAXCfZlab/4YkuumvkSxiR7masICip6+O2SZeZYaFWSlRhbaczDOTD3LJU
cFakF+Tx1a9aU0gXZDtkZ4x0eX5ZuV90ihmQYdVTGFh2+NLsDPKFsK7XELGYwKKYTcqtbwNaZ/NH
ZUEL0WqKZzmTysUAiBDV9hAGivbsrusE0D5ha02ScQ/MWBxIfZ9HpAiNsV0UW+JKgIKO4ajXHPdP
nrXAdl0N+4uO0v+d3KTHV1aiWVxiNbAw8OxF+Y++StyyliSgSCAAo0LM4mRZb0ZwpvDlsoGASD+9
IbhwlQg6V/R/5SXhbkidKnx8Tup5JDK+TJ2NbWZrYMb8GgxdU/JkxfP2DX4bmTdSeM5ycBdjXY9P
ZiMmCz4bnz2W03G1C2g7MihMIRiT+6oiL6PVW2iGB5D0LS+K1GynQMt+LLZqtzuuFsDlir0Y3m3O
bRJgppS6c9ArwAB32pkMSRbupiLc7pWvXOUiwXR41siBn/4QZTBJIyyQ75O422FsPEu1AVMybKlm
erJQDFjrJKwO2k+w1I3watmI757rNRXAVFtdYJ+ZSFC7CQrEDy4fkDv0cHa+/atUHG15ITASja43
Dh/HY+Orbbq6ShzLq6T23cKggbQrpr55j87mQhGxE6greEuTCqjexqbMwWjGOaPBHM4N+Fcs4yQ6
ZAAtp9COT2AMFTBxQ7ccwHj8MJAVeePeI3goI3sBflOpwWZQSo6PeSAf/f9GELnMxpdnWWJvL1Yj
c3OELfIsVXB4AM6m3DYVpko7MOEsnzGzCvN/1gteGaVI0iHqeKzeCslzWxDrQkOIa4kI9UW7en6Q
lNVxve90oi1hDlAvU6j1oHZACDDW9jTajxjGVJey+oUU7PxfAbI5IaZa60qZdNSGmikKWMdl293G
TDRvndGFm36TOtNl+YpuM4Nw+iDkimbQjQ0fUObNgcIge4Ea+SOLvk1filXRllSpuOknZOs/HpHq
1ncPSYTkiqZIu68f6qxh4NMLajpxMHe34BQpQuIbJFmgJr1S4lavQ7AJg31urT3eWwnxB4ejYMVK
C4/eYqxQujfO8OhfOK5F3l7WB1mj1Nzr/rLJpijJt4FVjcuo9bTwM4aQXnAVN3hk/jTpFqkRjLcq
jbVCWBrvdQg1T3jtpwRgd/OVQ2PWfnHdGBkWVyewQ/aRLJC2QK5UkvWx4huUq4tsslJQs5VMxC7l
7R8Xx/OK6iMTP0ubZzf7TXMRT4wuWqJ5YepvPohAtxZsXyl+otemlWjANdrkB7BxJTJRUmYmgVWD
O7TXhv0dnW9lrQTk4fwURYXX/yKlSbel0Jgdsy11KwLDeCwYGFtB6XMisWBh3K7awQ5P4MpX2iyZ
IwcycbJJv6zq8GuWB+GthGJ7T4zLtRVYx29gAycXA9fIyXeYaaluVHb+PNHouAh+vsLtvTxPN+zK
fgX+qIGLHmrQe6d3sblqV4Nfcgb3lUWldDh4yOL68dfFjX21fhahCwBnhXr+SEEu5n1GiEfDrOfF
JnZuTdcOZWd0ISCRn6jIm9VzGaOuV4c5R42dziWp9CE15ltG51uU5MlwOoRS7jfmp0tMx8op8GxA
W+X6i6sVYO4i7UQWS4E+JJtG3bcuU62Z/q1bOIMR7rGbSEu9sG8vbW6huhGKXJIjpINUDtUPAQfh
ppgV7ZjuNAqP9qrOm5OHYoW/5PoCkECe0cpNw+m+uydCm1rJeL11qZ80p4mBrCveMaq4ILR9/H1/
E95LYBLk6y5HGsyrL37sjXHF9UVrROheFxZo8cDLSVDCBJ8tb8J8DVUozEHxPVHIDpGAEGEzH1vk
znLTjpYl6DNHVgRB79X+c545944jfyzqYWkR+ZRYy4r/fx2Nq56DRpmO0sXMURGHieAiQOR3XRCy
e4+o+AgtbcSqUQECzbrWMyLZmwu+F83jEs0R+WnknKcl3PQmNzI1TJFWvxrOAbZ14Ls9QO38rC/i
ZF1KoBw56aCkvkiLCvIXtSqf3EVXQcTm/9QV9/wNJFKPxLsKYac0sj3cYAreDobrNudcjAhq/zIL
1I5KmD/9mHfLLj4KK2IOWmRitcbAxYe4+oh5lscAysf38w2N3vs7IeaTqJ8oFYXXEEEGjJziQOeS
iuo5aTw70B5UIR9vgYnECzKvvbl+Rz7xNKqjQIItjY965W3FshYme7YncBASuh4FSCDG3NQ5l3rw
fzQ3pcCaK7R26NU72l/HJdIBdb5ndcWhQoqFDJ2S+C1TYOia1N065vqOXvqu7kwcfyC1LSFxY7h1
Zt/PYuRKYMwTe5BBRAv2gMYYgf1eI+94YbD3wOkdNmNw2u0c07Py0etFibzCxUBbC/sTJArWEdiI
98NXgTaHz90znNQiJmZNNPTtPWej3TtXQWsyn6xzOCL5SdqbmadQWFGJHQuarbHClUGCbYwrBqw3
ndA81kHxOotN7jvOt44mFZufU5kOWpyvH0zO5qd78Bl++nAVNKsr/tXha7S/y2Y4CiRjOzmnRHNO
VWJ2ZwuO3IjfOW+RH/BYTxto+sFxaTCkgYuhE1bT6NWTFuQ5A8umNBXsDHpF6UDi+QWhxBypRXQ6
gWHEL3hyd1cvnpPIdv+vRfeQQXh4GD9RS8BWynyfwHSwdt7l2KZ+SklxRejXn+2StOH3jD8DpNFc
DyOWq1tGqnxtJv49WPbZgfKB6+BNJ43aToEWUs5GQHVp349F5boVxFsfiYD0UKPoFXnXkvIvvj9k
dN8afCPbu9bIlXuAWk3NaH33AyR1djnAIcdtYGTD6RxivelFbZnd3+McmIxYvruZ+TlSAme/Bh7R
XJOwlEfaXrwlXda1RLqsW+5BWRaoKAAWQ+UDs4NYwKM8emavwv5sZUBaWf/jTK0B12qDih4VKINS
G2tEFKQY8LHL8iBfrV1iGIFaAWgBnxsqnmTlT6JE9vcovrgTDI+cTwBlr8mWSYUWB1XiP7jRjcqj
ps6mIG7q9f2Y0jOIQ8aWrmOollGTFQ2d8DkpFgXSTiwp1FBOXP4Y7Rm8GifS/e2VSlQgykXBaaZM
rdBNWxAwPL9kzd3A+XP73jsOZZWoVEH7pR2P0a58txdfpOZWXAgNCibRtu0FoLTROFNzhMZoR0Nv
ZiQSyMIcFhrfiqVpFNI0SaP8PWXFGQ62im26ZO1zU6fHyOAHXEsvfUBm0CTSUSjohRsVJbB/ba2+
aUfz0YLso9pmrNUiIuBx5HlMA1W4MdKxV9ZTrOqYbmPlM5b3qqu5gFxtQ65d5iZZBUMwwVbdo3lb
HIixjzuNttlf6V5CZWxilnaG26MEqmz9f2w4DO/2HmVm0bq1mW3eAlv9VT8GUUvwGbaIqx/WBgOh
CQ1kgCYXdvsjs/JZyNr5eDcvovTlIKZlxhOUa33VtLyqcd1X5Uc9aKYUz1fX3qhTYEIIWZuxeHzi
fjvu/JtOAub5GRYjlIsQtFvDb4BS0TBP/0jr83LhadpkWYFaoxhSGrnAxKf9/WfRV4icmrN+IM8Y
MjxDm0mDHYlS3IIOJC5Zn/tnQDtDet2WjYnaIMpZYJ0kVHo4Y9PXfR+7UKNcXuIkNWafomGMjOcF
C3QU8s//y2OGMMg5V01lCtTP5ojPgjt9saonarZ1CTjjd/dCfeEqVJinImjXea5kLNF10qtDw8/f
3mSZOlyR0PEwaX0Dtdp/+/b0PoCvSyZTarRRVtJ1zyD4Sghg1vWfkzmusg9oBN5rhxtbb/34SHBl
lmoQtS5XcNtqBWNlGSny86LOHizyxLCZ5JDuDiorlxm3ECWt2SX/VoINPaueuz8iCUftpBfhbsMb
dUNwfxPo3Rco5qxmzFEFNOViWXrQpWLO+dmDzyIWV5nccECtJHvHUjW5YRlvX7mSAgGIEKb+V+66
WBkVNCErC2vmY/bVYm1/EqJqy0kyFvUyjE3jJN+SgLqjEJoS9FeIQqqjt40JYyBM9w3I/7knBbeM
dKEHBt5qkssvIhNygFWVxzFQ/2xDVXV0h+TslUXYngz4bYyITIVjBYjOx+9AzDp6GMP5o+HkNAWj
fZSEoQ7pPWoR/yRgXZmBxzFH2Sv4cKHVKyjiiHeN7ZFSSllw1PUcDXgN42kPuLsMntxCNheIE33k
rueHlpmv2NWyheg8MUP4ESEXX0lzVdO/Qmo4bbc0djtilaH5qho2Obnsy/+YNYIeZzHgnH48hWG+
KBX2pVJ5ZnlZi1t9r6tjid2yRHeXM+VVp6aPadEo1Eie2Cv4ML8b9/IVQ5ua3iCLvSYJl15PannH
z40oibVJCkYyxolSKL+7hpLj0NQ8PMdXZYWWlxUce4u7m8hRjYsCF6ivrvn9Vwj1p9LcIjBzc70g
cD1rIm0c6w1/N4vD2zDj25BLbh7uCaGTFT+bDNBE+ec84Y+yWlZm0YaW4MUA8CR7tF4DUKZIu1CM
UlhY7x7eh/0wxLpD3yc6xNIB9+/8M7cuNr5ldkkVSMiu2AGBYrdYFBwvRmYHROqIXnIjkY2fqosE
pu/IVk4bGKUt9tBxZbRX9nPK4u4T9vs86KPVeDQuDng1gZ1QLUnxCgYzOu/OEUbEN8UOVLMs3HHR
85hbSnwdjXjGytJgGMta8GNOJtlmQiZ+tQz9j/BBoc0bq+nypSNSV0MtXtY34dRZKqiLwHAFc3rL
nTAN/ePSjh4fHpwsZisoDPmM5gqoPBd0L5KUAJnv2+Ju+19hl6wQcPRmnlmAy0jGO6y32u1Ivz0W
p9saVjqF9EPluKpZJhYz8mEvBc/j1t2nkIwlP60/kM4u/mdgJlHihtZ+O9o6bxMSPbEu/REPkI9o
VGLODH2QWfTfc4EM5WxdGQZ89QxedkbiomL9QkTF35nTnitG1nZ2aAtHoZu3k41FfuPLfgpXbK8w
jX51oBiqmwL7A73bb9WDI5crW+nXUf2Lvhx0aqrPmby3Il/ufZeUlirTCqP3drsahmvChSCGO7Z7
pw66CQ/cTCiuN1q5Uwvz5BvAauwmMEEE6cM1DZFBwzQ06yxPZQPS0mCT09oZf34F70rghwsommOS
Ts+7dVHm2/Z9FahfwX2YeuMr3YRwVHTe1Et4C/X+G1HMG3zC9jGKEZ56cwIaNvB1FVFw9MqnjCKu
iEsmVD2bAhI3+Q9V3BQMivbhhl3EKLXUmXdXb5E0Jw4b2UPRrrjGvcvhqoiCphnNeVgP6f/51DWV
52YX2hPT05O8yFPYnKPn1Z49swEkthHCKUw2bdKPlj8wTPyA0RBTpw+H8kPjueq1fzzoggtQTqlN
mhpQl5lNoC7e8XaLH3UTd1QRoMu4JyB2+mwrI9+Ru9bz7k7s2i+25wG4dxIhlNl86YvK0yUOgFDq
WdOro4qPp+HoTOxj2J4FPuRZ6A6Gqu0a+r9c5bSsxnw65n0xNj7lCNDVLfQtRCJ2VffScIU1/KoQ
h+jwAK5BKbXfQTnw/lH3wwnXFz4e/CTx4wHZ76xX20XzqlpFsjNbfCCu3faTwTzBt6Y5D/8KF866
DeseD0uZlFDZL/MUpaCbqdEzEtA2u7s7PUmOFc9fMnKLRcRIIODDy5Nv8E4ID4AxiQgF/NUfKMxH
aGipSMNiHeg2FDAapTDiw8zxaKPxbsi56lE9eb8JPSBHyljmrTni1om5Fo8jC8F1wPw92ZIWCQUz
2UfCnyx/4ZjkKZypw3WCeJ6OP1mBZ2kmoTQYGebBxLx+85aMurV+727YmPLulxfbfgBALdL2G+2L
zOIcCqi2Ykf8CdQSYyttnJhaX1fV344d0LtDqJdm8i8O4LziqqBiRAxzC/r5mIkUQua8MkxuBk+M
J4xP8g1tk/19GrgkNhMeAdS6eNEPuimH4tpQto9tcZZV0iIHR9VriSoTFHV3GPwvQHXf0zaZS1iI
8HfpwMc39h/w5AeLB9/nA51EOzT4uxg8WKhg+2ukNNIc+o2N6KbX89ZvsCxgVrTNqpJ8WY+LEBkK
WGuxK0+wTiw1OAwZe3+fWt6K8A3w0BsAS9A53bTVpQ+nvLXv+jw19iz8eZtTQ6kCJ04diycUnPZo
u0/w5V/wFNsnNdEunJ+LW1q5akqw3IQ0dN/j3UdJJJ6c054HXc1FdeN+7WqkFXRd176wtGGBz+UK
S7xIPFIwWmqBrb7fn0LC73AFlOC40pFVQ/izF+2O67LIivPxUUeOJ5U/B6li+eiP0K7qloi5Me5P
JDltM4yR/o16jf9nnT/6M6f+j+nEGS3hlBGP9Nfu2TT1akSN2KEEzG0vnF8uxgbQq6zxj4O7ep95
eVMAKJC2jm+YIsSvO+4WFagazoO0RFwo9zE8nCADKi28P7xr2Zpa5yBYzjHEhN2zyso7pM1vaVjE
FMwME7NuCiqOJSDdIt+/UPUoiqAl2RmlyqIMFl2nd6qco6JA2mPrgovCpcx/s6tuk+ILaCOpubdk
I9NTAN7EcldRUCuBXXhlPHQ5+sb0ltcpMVuYL5jPJckSJPUCvhlbrSxamFiqvtnb5E+B1vTSbdaO
OlmiJhuFWy7PJTy1KqDYvde8DctNg+y2Tfw0qXs4L/n4SOw+eP8khU3E6mcyyXueTpZq9TbpBpbV
DyDDL9Vwl6tCDqww6i4dbLgGUUvv0ekLt5nv1yZbuseTg86Aw10I7a/r9SLVYfqHVMd2BPx3PSEU
3yJOrDmWkg3+9fQ+uwduWn8epddp0O1YZufwTADX0RwEl0+dAljBDInQ7ws2ZH6bC4BaS3BAHOFO
18hLI4KWb4kIcEp8Jr9I7L5OhXvxre6Ogc8sxKQ2LYCN1QnN12d/OnuRKX6QmhtzzqF/jC6xjD2L
6guOn1cOBQL22Mdfc1Fy+oiW0I86svoenSb1ST4V6f6+cPUD1l51lmeeJw18NdJ5L7aI9sZ70flm
9rk+cz5nkrO8UXzbfM9Q+Vy6A6K/q0+LAp6mSTWExsug00PB7jw9Nd88wf+2jKTagyeA9iYJ1ddh
+5Dwn50mcgmlA4WD6DgefhKbKp9ERczoG/nD7z3Kpi3DASixAn2CgalFJUJQrKyztz43DH+Q2Ja7
6ddZe7F3PiOnREECCYvhW6QlT4ypM6ldaVLl6BiY1Bpu1cRdUAxNIQ4LhIov1LoeArNUbNf767Tq
bLG+O7528d3pMKZ1DitgVksSmwCIjFjE7wi/WyiQAMyMIt/ZiqhFvo33GW9tkoUusS+LTSEN0F8s
HdGDal1HgmnaLQqNJpMfsvnSor+jZvVdLy7uQtn03j6RzOwi82a/76Aw7u2ZwLmIfkyFj7bbhpsB
YGtKe967m/T1QCY3b8PRl4+WcBbTpCD6mmZyU5Xmk04jOce/OwawaSJ+jaSQ/By9wTQkjMteZhSB
2MmtyT0KCK5vzRafXOO8u4+9mZZjmygyNqyFEDvVvgKqSs5DiDoOCOYSOu81bpNNktFCxShh0YJ/
lwYvG2xKZ79IC1OB8IDbdXpD2UDtZx9QbOLi3gVuWyLChRMJ3V5wjokF6i0x3Gwas6vRWmu1Xt4x
660oLElFJNjSr/ZbGyNOOiv9llWubjB4cmrm8WCHvAaB9wIn8dz2HYeUHahLOQ6Eaw/tHDCwP6mL
hDh/L9Dcrwe7W1oV7TJxiEwUKSAzH1I0Vqgdom4q5Rjtt5t4O8vgGRnzwhlr9yTijrP/eNYQBwit
0i4QZVC6DnUtj5HnIOJwQ9e6TUDYXgVQ00M/UL/uaF1WS7P6AgsYhxTp9DCZe7bh38/UIIF1tMsG
mZvZdMsKOd5Dy0jlpH+AiPJpYDpwrkwgq5Cb7M/Cl/QKiUitqt/LN0BwuqfzhJgQhUfLRaCfiFN7
+7KsPctEXt8Lrozgpo0iCOtxkRlwt3mS7fJ9ang9YGc1j7sGxovTVqfrFX9Hn2dO0vd1slnu8OL7
rdIes2eG6Z++OARLp9kbaS+vBFR5wNODmX0HKCjshy6xgvZ5kqJ7iIpCr0IEtz5aPoLTS9+pFz6H
SyLC2qQgIEho5K4L+U/mMHbfYFlFHiV0DaOL+Gsph3CQsp14u+A0JZ8pLguULzYgn3o7tamuxvIQ
D6m0ry15DfZwRbpZOqYT77EdAcrAUPPeHDDOeHqaLfCye4ays/NKjowDKGZHKHD1rYBz/w6qlw2X
8LAJ2SOFJb4FItTfjdhY2aE/jc+DcJiMBuWjgr6Cs3D0FXIRXdgiOjFEn/PiLajESU26HlGOMr7T
p/f6UAFuSDWTfJ3RhyCaZjcIo2xnQEQVLRt0VVINwe2KyiMBuOZL6okCXZ7JoVDVeIgT1FNE3Gdh
d99lW0atISaGJLb6ytdz4TQHDBgxC6oooeh+6LTS3Bvg5SChB3YfB0mM0422llEaoDT1cMaSTbxu
iD4uGTr8tPSD0loYbkoz1BGywwD/pscFGIUgm5POaOco/RtQqgumrAY2SMXrByTj16578ioTXzq8
u/hCPw/TReHxrtNZ7070oV7Q2CyrbUKpFjq1B+MF0E8uuyWVPUBp0RMZclu5ITzBMSEmmgtmvx5I
c5RO3Bdn+XHhnuaOJZ5Rub6DEuniomyG1GHlvFAF9jBFItBNQaVsqVztrR6c1sd42VFEmhy95d67
TLV6YcLYKi8XlKpgU75U57uduRpNRR+ASpy2cjL/FOr7t5xoFltc1puENW0Ay5lNxDGCho1TmATR
T/SvJjvj7zWFwmqhYcZimkqIW6+q8Ewu/QenZzPdMCUXUMHAxqvF8TM6Pzw6UQrZRJD5WRSWKD3x
IIdqc+b0EekLUXBxLe0XYYN0kCZZE08ciOcFrNeyxUUbenzr0Fp2dljUMyp3h5E/sRudbLWXjsn0
sNfNMr73X9LFbrpr1+XKWMEFNxWJraOXFcoffalRVrVB9oZnk6H1FVBN8ZWcAyRdn+ilwhRfMU8z
AXO4yQtn5ZyhxK+ezoD7wt8CArPyRkHiXSjdbvOanZoHjemM6TEcg3Z6KAMQD3He23SZ5LptCnCR
1sQmiatZ7rRVE2EWWgawOOx9cF+mg/A9jEVdf3k9CGANYXQSWt6UgFCv+oMYQs20d9C5O1LC3qJX
LkDvGWIPdKDM9lJ0GpztCVu9xXDAbEPJpwAyYYKEaTNzRxPO/4Xyl1Q1IOGoFznrXIwf093tUbiY
2uL9f/5CvSIDXXSprRO8ZDmxwyZPgaZcAMTrkb/jFFl8VTBbzdgMAXraVZAvlAM17qr31zZe5cqs
LHi8p/TJ0bZIxM/X58wHgfk8Z690rYCk7EXjLPzoMWIKxlvp1I67hrQVLMN1Ts5aldegtYJ6ABcz
Zbpp2YJ2NLaHT1eiDBhARLuHQ8C5Dn74lFaLyg3QhXa/tkYJj15+Ib5pKjz+ljC7wbVy94Kvu3Km
QaWvA67BDbEiAmC1TGPE8n1TWHT3/cBAaIY3vkBpOtrUmF3qh8KLt4xInWusQsNaJH2CRWMfuus+
g+5jF5j3WrZNP0zND9gOjfCm8EejuMF7jaWdRjVzCr0LthjCdHmPHAA+XLEoFiY7IhFWwybXTv+s
DR6YT4yQPXRfS7uui9QOlvmJp5MJsKdQVNaYJwBkIIOfuV7+M6DKT1vEiWEGR6bglxRLn/sqnNZR
Lutua59WPN7D8+uLB5Ol5CDrAwyV7VwItWcJcuyupKj6ogPbaWR0+QeNhvTbaL7YLRCbKFRo8qs+
XBFPiwU7jggEffaPvYZii4uByS1tIaTyNJbDJTEZ4KD4Npv9vkni/MlN8slbsVqiWQ3vRHXUzpvK
wOFHJWFkCDu7uqfttg16blT2z11R84biz1uiDhMuwL3yiYiswzMvjmZLNXiKtiDthG5gBcfUvJvf
dIRGlK3o8RdjHgPok7ZQ6hRZgIuEvu0rC9voqE80Z00dh/1ld9VGkopTnEOTie9nKoqJCPRSnqiu
AoP60eXGppmj4M3fsq7DDfnMTSph3u1EOwkXRQIaD02/0BPleSrR1Cs9mhRNgSgssex8fJd7Sm+l
WEGPf9kIal4ISFMdSUClb/qzuG6wZlXyhc14ty6+4WryYI6C9XgCiwju/YlDOvDEo41WKjjparb4
jCaRsCPilBDeJEPE1BYbYph6LAHftPK0dRKZdc+qi3n5+8GafkF4hpwJGbGvCKa5PgzRuMy0CtPs
+9589twja7Pm5Ki3ilfOBB26AYx79AarMXaA/OfWWfe2eP/HqViyaC9/m2dKRRcvVQ//DxJEDffZ
lvoSE5kFUTRWKxB4+ksH73vrADbZxkZBwuRjJ2zZJ34DBGgFVGzi+amudLboPC3UD2LLhYH43kM7
2hARFzwScKVzjDnHPDOmp62S53Y4p2CoIy079svKnUVmiqlRMZrmc+oGhT4LG29XZ0vg+AaGFUTp
2MIBEfrxYzyXfhDIsIuIueXdVpguKMOr91Vum8jcbUrotW7XjyEuJRSRKKKWDsGJhz1Yc2ZHcr4G
NrbN26NgqPefa9hXuZ0mlJOUoBlG+5UOpfmBqBwVER1Q//IG2zU8P7l2JNY/cIGz704pwL+bnL9e
+67Etyc0Nx5gL2ZQdLHGdmq1ITPlsXmQfsHGI8m4md0SxpopDh8xFXwQtsDs5zujLwt3klj5i2Fa
XSRQCHf3YD2yZOaUJnMD2BI7GMW+xhrrV65uZ702lWzjeqWa1OvzMNBTQIC3L/ggvK5giQjC53E9
d9w6V41NtmUSm17YeBSPDVmKP9+thTmPS3elLLNxMtr/fq2ooYwL/EWG6vM9MJLcND3fEGiY8eID
528Er6j8Tbebr6y6epLNj7MyivyWewiHHtsXnoZahVL7Uvn+FXqJuSGEEyxv5bDh5pVbic09kM7v
Ubmw54cIGUO1AvEkqGyc1fgcPgVdvNAjsZdM/pfDSQ4xZsDW+E9XNaSZusJ1AJJjb+MD14X/fusz
2spwD7CU6q2es/9LY59Vy6HMTR4jEaR9xJEEr36W2oGmAkL/OCcblokBKpPxfeTRbeIk6/ak4fUk
Ld6iVi8lJxt5b7JYQii5fZMMRw/OOJH//bKr1KUi3m4GpsOJPYvg43Fd0QAVtr3BLPw/pZuUT5GH
FeGn9rfzpePwM7i5denOZq7eqor526bKRjrhrUH+bXvnv0vObzaO30Jqr6wThiMTUSsBCFVckIMy
JinLT6883DnaN9xqAQEba+0sABoQhCyG+KRJvfI7q+hBiEarHxKnZaDhZSXA6lQggjgRBcWoVAuC
hOFDbCBPw53/p3dB8LjzEPVjYgdQr5Wjrq+uBR1yyyZtTuFYXBngQPvQNLKZ7pw6XZM3b37kfgHp
fOLqPHsUgj+Xj9xmWzsW9TJ3eSgEGrCugDsHhlupuiVKq4Hlf8kjTweb1ymrzzn8ec2KwamSxY6C
jN4Jg0rMxIYSeMXo5YxLn1HVy7lbCb6py+GgBS7LsnJaZEeOsQG3IrcZxhqNpjtKb4TwxLsuvTnx
uf4OLIMqAyoOtJs4CfvzGm+Je32rc5T2pWRUXqjG0rIiwDsxNHQnMgjqPU0b+iDxkQGxhe5uF9GZ
84syCWVdPPvrNa3CepPC5wZsHLBeWgY2XGxWhb+5l/mf9si3HHo/fA1dnEJ7er8LsiZQ55MnkrrA
vu5eLjBwhAN0Ma21FXQu1MdalX1LJ8bayFAkVfsyJ79OPXw5IopoQU/d5eCdhRgJfkcdJqlfZAIz
N2aWuLiPrbiiqolksh3hbcW/LUauHP1/LcH3IZBLF/lSJ7XQbamolopcAgW/3LNgH1g1EZo26R8f
jPc4M6kRB/D22p4NTUwm6nHe7uhf4lTvgQRQi0AmeFJlXaJqaS+Nr1fxrJnUjA3/ilQYtysL+jJT
lG7LWh6nhG4Sel56qYzbm1ocMmBXsDZ+qwBBq+Lhs5KC3NOoOQRZBK/x09FzKFzXYqFjeWF2Xp/z
6Lb0n9ot2oJ14WAq0MKKzrfGBVkR2zyBbAw3Rfbc9vBku1QOI55VoMeDeOHYq0bjCIvsyWip/1DI
nBQJKsft+mt9KhfGh7mp/NqgCO5ltyhKo26YJmZNpVS8DKhKlnXR3GvyRJmKsordfEZaJxarmLW3
2OT0B9UQBGW6jIkOPmqJDyyGIhRCs0UI2gwoNkqrJ7uPtJ2UE9imbO3B2erWr7RAsogr19UeKnjS
x8yzj+N2OnVYput/M3DkvqQd5v+hZP8OT3/Ln/JnWwoiK/LZ2NfC0HMbhujAzuNr01pK5FqYk10v
Iq80PNL1sbxHspvbarQiLRipqjXkkX73n2LAfr8p1Ew8SRV0jXiwNgUfHtMIt+Xb5IdvxYRmC4W5
9/7SaK+GYY85C2ejvqpZT7bMl/R1ow2+z3fyjkY4nDR4W97yF0+VVVYu4qMwNIwZfB1P6ODkTr69
nqkXRKo5VXIrIRL0+Wb+HP8qRYG8mlHHcxkXIGqKU92wAwhdCIRTGg/AlPGEfcNVBeiKZS0Q/5jF
ZupnV0bcd0Vssgj6xcnTfFG8osEI0GEwMpFj6hOAMozePCzp78nlugK7HZcRG0dI+gtQcqb/PXRz
k5rnQO5bUhkL/a8/oRj97YSRjBwxspBnSuxc//14TZP5Sr2vyqFpLsfqtW5/qtPOedp4JfilbV9A
Exp5IO53Ssi1yzF8mdd8TD8Fya0l7YR+owGRSEt4uRz8uZocZJCLtBz7gkmLKsO0al6s1gdxuxn/
Al9XzNGIBk+5vH3K+Bb89cW09gQhazzxweLiPj0kkFUW0IZRMG2CTW/UdQkSliA9xpNgX2WoUTzG
fiBXAEyWia6mqkVq0OvPuGSR86IA/Z7MJsSzUP+jcU8RCm/uZdBK8zF5xW/4GekQFUJ9lM3M1FlF
qKXHdNKQFMSK03tv3rS9ITgazlN5NqXKRyWc8o5uH6bIBldia2ygZ5ZFfWJq+weFOeD183Cw2d91
PmN1hCi7/sq2ivvxcPA99OhAPG+dfTGREnvsPQQGgS6aeyuQ1wKcpt73YWYqskg6Lpa7Ni0g9456
MiAPm72X1HNSa3RvJXb1yLQxTejZKPEpVAo9cMGjdUxfm85sRyDd0Q6LUfoXnPh5kIavokwpde/G
pha7sWEXHaEXEGi06c9mOcPhckTBMikMo9diOW+3L4ixJ6FMmG4BYJNX+6I32hndO6ifcmRtcwod
EGFi9Xbtx3TzS6obdq11LmFr8G731ICITgMjP2iK3MisjT1BPFOt7hf78h0XkzzG1e/WRX+pLvOa
EODnNTTG92545AR5BiCZfLasP3JgS2dveq/GMQ0HYtc8V5V077TypVP0JzAZVp32Hkl6QpTw27wO
6NRybUYCoDVeaCXH0S9sFeEYOq3jCcZGAKf2lhKORWFpo8SGYa2G07HOgPhHB2h2YBYbKw1LMKcH
lMeHzXAODTRyJoqcDK94mMW4kYwWimtW4FGJHVcgmcqW2xgVbqVxB77F9XLc4ePxBmUf3s7EXHca
/4MDirxzTsXaURmaXZ8spEuVfa3ZfVjypXRRsrU86OfOK4t07pmyBh82H/7XKVQrJxTWtio6nZ8B
LHcEjk4EB7HMZ41uhI6DMg512yqAtZ/RWM41LTQqrgjw0NuWBVIqwBIwPyon3/P0cXQw7Fb51a1s
6ZPX6ZPsp6AEE4sb3VaVZg6+WHK3HvX6NW3WEbqmryDvW6McXVrq6A1WLTQhlnNZwk27gX9T+S9w
O/ifOZlVnSgMWzd8S7oU6FVEOfDNUXOAElQ9aAfTnZhCEEfh40q2cB+zuNYtTZt8wxQKsfGsYarO
yf/Y34dqa/5QeQon7BNIBGVRUD8iLpVGGDgooohpv0F92/NJqTfuZ+zPgPEqJG1Wz0EvLK/BcJF/
uDy+LuvdfgaO/IST0+VH6w2JdHDlXvFWTsq8+fp4ztIP8FgifQ2ZOjouCEd5rCVA503AwlGbSJsH
ihB0O8UMPWsI9/3HKU0WRrKjKjbwr0SiQgBgpzG4is2zkILDFKS47FMC8xrbCGk4Eh3mMqIY6K5I
V8ZCv4goUptlYvDGDYMo15PpqJpvtyORNPmyEJj4Fx76r9NXu3Z3wCHqI60JK0UJUF/15PQtDObg
+gtXguBkiCdJ73ImPHiuBL8uTVrfRk0rOJhBUpvqv5yblrHosAtRqkbNNtK1pd4CgKr0G2HYyeh9
c8uuPN2OUGlaS/RAIgKOrzx2zKxjDMrAVSc8KIc2Uqv3nNh3qCC1QRnVkQdBT6ip1+lf66N+XmBA
WmIoboxslJxAIKwVn3/GjTwQdSwku9VGi7ww8zAacVWEqcF0BZagOfD4PhqPgP6LZtk6pwzPdaKe
0ieON9z7bqgU/JAs7e8Wr+LCS+NIOSPclIoA4vBtOZ13bFx2/5QMb95bxv0xbp4iOgycey5PRcGT
Ws5ksLwwVlMumtUFG3v7tAf0BskGxW6fLUc+YeVP0mv2poF+TAs4NniGkLVT1E7qnEzoRVFp0ask
u1EBigtgdELFfKyQ1jrHZ3aHh20p39VXJQ03dY1cGKH0fQ+Nyev0gjbuC61FIry1ykFjDMAFC/su
ydK4+M0CGPZ/RBGPEV82iZTm9Oe/mkj7NysB1Ym3D4bIVbvIJW8IOlxXq8PB38pXwk0OsMhNRuKp
0CP1dOvqYL00nLsinTJSYmteCSW7N1JCOGZTMV9bpeLv9vY2gCNdgq9WqSGRoH4g8EDIvK0quluW
EBpgFPXQhqjuWyVR+sSeLaeKX213OTRAcWTSQbRP+ZJ48BXzbyLM1lTDKf4EhHh9Si2Vkcf3MvMT
ht4kNAZcp2cxVlCWlFuOS6CskZRntR7FS4O2JATph2p/lctfH7GWG5hsuxIf/M3oMQ2AOBPIHm8A
Oy/ANzdGSuVNFtxesw9eW724GO9cMXHwEThfXqdWStbFv4B+LH9BmFHFK6p09ok64GzUvi15leU7
coEoqYTKpsiELWbe6ZFYPVKAiSJVdXBqi0k/PdtbRTFGS9NmEhcMY16pj5TeGzxpt+Fdtj8Jm3ak
9K53S7g7AWLbnDlVYR48tBy80PeE9EyA91TXX4gTopwOWM3JvuzyZVYVi5FpNFPjZHb23DzCzpIZ
jJ+wQJyDIJrHHC9DrInN0ZWci1aAia1gFEGmFPSJJLILCmicTd7yaaonB4zUN3k0imbyTAktSFwH
VD3WmBsJClIBA+4ggv/F+xtevrC/16JBLVKs2f0vmt1OPDz0ixcTp2ERkKJs1+CTME27QcQphXQ+
QupovBwvFDnjIcWm9g6HpQmydDolvQY4Kgp2DSrCKQB4G/YizqYqD/9UPwGQWL8BWB8zyKk7ITdf
fJhN1q9MHM7DvZl9HrLiaHRLZErB2ILbngmSm3E/5FcZ2TtzJEZBrfOxP1krEK1hldsJhhmdAQBh
QSVkkV3MPrM+MylFQkMwkGK8ALOsyB2pU+OViZp8d7oQtBYXWKPh8JCIdE8Tju7vDgnEA3dKelvy
53u+TTM9+aCJFiVP7u46ikL/Spu6xNcwo20A8aewGZzqHn7shwveD4CALDBw6m+uDx6joAUGiz+8
Vy5D5WtqRJdVTuhQ7aCnbdDJMzCwlF9E/CVmU37ILDNc+UNJ3Z6aP6xSb2S+C2Eyep9LeOozODgF
H6uG/UwI2tK/O5XXjKofPVtrNcZokDwHp/wPUD253+S6/KjtvuUyDOTYv72qdMro3KqvPEd749rt
w28xn1YlfrDcEMnHETdiTXADAV0jKGLBSLQrLMKjZn+d2Ac+W+pc9z9F8akHWLHzFW18DxyFhmyo
6rCsTHRKvdYXh9XjdmTYlsBuMREdZ2gdXxrQwZKHaVVq+xlZ4JtHiDpW+Frg0epc2TChVeq/SUdN
/ZdkdBhosAiC4I0C9e3De3N3er/FLnRxFyYF8RGiwJ+6D0iGErkHifup3RhBrOs1oYeVwb3RbWTk
ZFtt7bST6nsCS+MZ9ukjeM1GjY3YBkonkusX2vAYPXOTBbGSOrou9P3ufZS4rzU8JY8IW1ayVtw2
LnpiGfGoRiMukaNkxVtCfZwoMdiRQR7FG2KztITPuXL8rhIRVICNCjnTU6/SYcPxJwCx2AkNR3Xa
L/Xv7oT+Cd7wHEdh0UdgqYLItiqOVZ0mc3CfDrX5kOOFLY/z7DvBcSX9TVY+AlBiH/8hE4hYTa2q
nG83j5uTfbOY6h9UBz2nHY5CpAJQ5P0YA+14Ud99W0g6xf2HCDMQzmxBPnuZU7ghqBXjliDsxFlb
dRV2LDU5Wk408fd2jfyYxUhhaeztLO3XspKEawQvmxiJMi28lxC15EtCXy3SEtvfHY0bwsZQXXOD
RjZgTuRn/OvpzVYZWFLbbG6dBN0IVMV1adcCQt5dZ9dtjf20l4wyFW0xHJTFFZg6aWQLGXEMw8Co
ZVSsdnLyTgIPBz6rLef7hrtz7/T9NGfI+oPJJjVTWiknHi0RFFunK7rBsau0qXRohVJitHOyPJCt
a3IGjBm0+vPdasOcYRi0oMzdayN3l4NdPdu512lX5MpuO0vJMPQBT0HdPJ0JJW6uiii18kUEAX8T
Znq5PwGI7PrTVYHjO8cOl8i8tsipx3JIr7xmXv9tTTcj0SHCv1SZfIqLtX4aOz06Btkp9ygrFeAi
8VEjO2VB2buy07neKy/pG7fx0P6OjZHBKfFY7AhMKwMIEEIur135BFUPVxeA+n+fWAN3Ov+bkSHo
09Xu+CHL9WJ7/prckKCgqsjxT0mUdbeW8SQoe+7GxLZ59cOD6O3OPJlUXvp/SO0JHePSXGqBq2JX
GY62RUEHrh/mgsbzAOsUrO549qoiiXpfntUEaB9VF0FYBKjtmzvXjfku9bzIuyQ2HZnQ08bzev7y
SAd6Biii3BnOu3bMPzT8mHyF8PBuWxKer1dX0OMGNc0m3z08MKJ7mAOpr8fKOZ2TiFoSREx2+/X7
JjOQcnFKA1C9reswFDY6ICMNirLoVKmSft1yIKJ4j8E2eMBOe/QgdPd88Fp1DgChHn8MNYGy+TmG
hgMcG/OSS2BhSqEK8JaG51RvGsIH+KNIDiXC6Q8FxiflDMUeRiIgiG4c/lcLqvVN77DFrkpokDaa
2UHYIpS8xW9Z8y94VaNBIU9PXl0r95/sDc7CDScrHkKcdBjbRXB8BK7DPTSBpDzI1CGlpU/NH9yF
gn+xMzFQyySKHAMaaLY3gKQ5IeM4axvc+6xNAwpEkMWrvsCyIEpenuzAVTTHKqrRU9m7Yw27pM3T
oHnzT6S5NLOel7KypeowzOcBhBPWfOcYMIr/np5QLW/3gIOzrWvOXrGFvaURN80akgp4qDvZJvuj
9Z+v8uMb6ESTwVZxxMrGsJinmGFvq5n1MNVSKTTAqTPWnf/psPTzfDfJECA5YCo5a4/tedyKQmLL
A+oTC3Mwu0s0Uzfc/l77mpIpBcl7oOPrmPjrQ8H2/ZgVopj6UB7bLC81i2fC7izcY7UrxoqsJvyr
2nJ5kgYHkcoIQTDK8CHLWYZ7I+cDYzXIcwXyFNf6BrghmzNK3VCdw+W81hYcMaEz8mQ+LBczqGLK
CYmSD+077OyHQXvk+qrh7V3crBXpVqOWsWfa1f4yXj/jYO1nN+A+Psq2aNerrQmOW0n47QhLpaUU
RakvMSxvtkj1IsBUQsWjLtbGXj/Filz3c+WKtecFxa6aqjkEZyECh4PWVUawKEzh2YiX4lmK3Mfd
pUdi8QY8yv6JS8HFlPHmELMx/jpCSQcDAHjm5BFORa2aBGzpWN4kb3sTh12nEQ60SmeutH1NY9WL
i+c6D9lOFOggDe7S8BpOs+EtxytBCxBZ8XWJl4lxULg1C23kcU64J1IZLezHRntyG+DTHa+qMdec
sZGpGRHVSKIkZaPoMi2c91bdQxi5l6O47jf1MydfgjlDgZATu9fgbviTIxRUIvVPGl3P1HMaeZx0
txzDg3+UxSKwtwpgszkWcdlz0s357JYmUUSmLMep7xUimZNXxoJa6WiA+d4L+L9aftqdUl3kkkOh
BwT/SkaTXpFCeY4z6ln1oRDH1cr5oJi/mUcvrnNXQuTr6HLGA+N/ThR8FoKGHjTanMj41NVfTNYZ
BuO/HTWlsQRmh194RQpcdbNLPzwNibJDH9EQSrUGRsrhU7lBq6cNlqelqKbuOQgp97R1eM+NrIuE
UU9p50DwGHRree993YRhCbw+cLmatU+4jRYGNpECxX61cecItOAfIVr3BiGY43AmrJZyPY3B2rlh
m51njvtDVhRpYcP5lFdHPLUIfOQFQUd3wmIVNfMENTtxP3RPJeJyes9FJxe1ngqY5ycicg5Xtrxr
gMEf9CZ/s+sXC88Tk5j7Dwi+LMKN8frwwjMVuRehgtiagAR7hF+shxqQNJvhHreph2sI/uqhJbq1
TnXU3Gbg4aMy7nIS2SP11K8SJS5kQw2j4AndTiLgUwEyEbKUjig1fV9xz2eEMizJPRIhVqOdTvPg
F7Pc6BdhbDrOjejM0jqwn8bGFX4R48qwZMhSRFZ1yDSvmOIIK8Q9NWne/7InmfZyYPgIo99GoQj2
dm8HCnkwl883m2/Fbij+HYez5H+DRoFIn66SHGnWIq4dcHv75CoT9DeqY3K711yDQszP8odMeBI+
Vsr8AK1RtSeerX0phpeBXAAGoj7PKxSLMlxpPfzDWguvFwDzXenNKyL/T+0RtfJr9HFQIu4lT6NS
UhfnjlYJ8dHUGL+yFqVwfQucT3z9+f4x9FWLbhS2hhXfH+fyytgVfChc6/e92pBaTgaJ8dNJ+HrE
NwMfsnF6xR/3JdbONcr0WPnimo6qg/0rm5NANg/0vvs5yR3Xtm1my1uWH1+SfyLywdWj8r+y00i9
xv7J11LJAIkxCRuJy+I4/tVv0XZmQFtv/8cy4NH7imJQRzXwP1p5NYeQo1TuA+iAJtFZPIe/whpP
pEXbGEYnkrpSgyd27e0kTeJ88NX64KBNMQltdMfm4Y+K4H7xeDseXNCGqaj7IGUMtLqb0UlOHQ5j
yOEhyuksQdzepge7fMAxWCv54xMlGlPppF19eid/CrENPGYAZoQsbpiUoPtu1xdPwqSFL2AeYU8d
2CaNGHhbgvrWyLPb7oFNLwLd9qiDXJDExrIA32A5RHTXVl7nG91oVe+W6e5aMnV+W2O5Hqox+HCF
SWLmUCB56bKhJDw1ItpnZnfF+xXNnKbZQZbmVjs/nirSavvxoXngTS+0dC6jODQ++lwmIzmdTEKq
Qfo6E9ssgGyPFn5Q0Thf0yVx2equ7EjHj63oIMIBlU4lSjJjGOuKpo6cGV/bnZQTqkuy6YrShTYO
PzcdQ2v8TfDJ9e5Xf8iYfatoW3TLqdo+TlRV1LnI/n3OzSJr/f86ZUS7d3DCEzB5JgfXjEx365lN
vMCX2nlTSa9gcXzaGWTJ13wjs+iZZnUUtt+KB9o/XUHpVNkSD4xEfZCwq/g1x48kh3OEJuKU/xce
UONoRf+QTwTGAKFJwEz56wchKBd8QIbWQs2YzYi+71vIjNVcZc+lJLgfZcZ1RNcPNnsqI8kU/CBT
u6OKGyG6KTxoZp3h7Y691G5dtxxsKoK2GIl1wFO8Xt9J7KcoLSfVVttuj2BWNCIBgbiQXXAERMfx
nOIWlMIAI9J9Rv+cu2Gmu8soLfLPqCE5zDBLWTY0pz5uXnCzJH9dnmLvnpidHadTQ/EKT9oSBx6E
QhHw8FLUVhGQh8krnDZ1xejt6ZVPAZ64AfOd7qPrW4Ia4dg8ov/XqfFlgx4V0YrjaB4xslMLjUzD
8h6nGZ/Dtmj640nTWsFthJy7QviK9fdrjbBuuSv5c78DWWVHMKGEnSabLMzfjfp50n8lqNG8fCIv
VZbpYy1y6KRV61rBddur/wMG9faIVRVjqD3CcFRvwZn2UTGkSvLKPdt8M32ZQ7sRZ57OxBxvTi4g
Uu7khFGX/qMxhbuswh7eeKY168xbYxwuHeyQ+wlaihwOaVytQYWhuTxAD2ySra481MH/XoD2+qLu
OHJ23pmULq2KpZr0F0/+7O6r5jb5PzlgdF9qhlPKTAtufTBWP4Fi4zYG2sflIqHM7a3VAuFFzIy6
IdPFcdXNRgCf+78qkrZvCUu98kDZtNTGzJmvpX7Pb26NPNabEnzhWVWUpXgyFW52yl4qbP/WnIXX
U2tY0eK57lzgcQ0ywg3io0yDvIl0lkwb9LJyT+oit7MYrPovvctSQzUq9+xpTgsGqLlj8F6UFHNf
d82yGYHM5bUdZ+Q5nMHjATKGsqC3ZpPyItaCW+010AgQu4vTVt5HtrtjdVQn53UGN/HSZr3BR027
h7M1wwq88RGMdEpJRGn9BedXhqi2aBJ3CNXusl7oeiLQOwV7ZZhJwQS3bIhi+EjiFa19CEbX4QrK
1dtyyYscvA4Nu76JYDc2M38YwIbRO1keqBRgCi1TuddL3oicjcET4N8A0XbUCQrw388qmu0x1fT3
yEafp3gtC+Hj9S2BfcvhLeD5rWXuy8UE3rG2aup7EM5XV3bNroBTFrPZSavh2ea1A284vWpqiDf5
CjTnqhqHVPrhPEVierQnE4C9Iv4+1azHuuzJYEflysP5eQrtefCj8e74oo4Bjm3NQttuDJr5JveC
42U628bGn+UeFTFNlVMiDA7G8Qzj0TgJduVLyMXS2/kAEFfm5XWFTf5SK0rYYaalOK5pcNe4gigw
0jYvZTQw2za5pdGSMgqvPxmZV0tOEjTzlsZNqiM4YzE2lIjQbfk2a9//i7PEV2wUSqrumsM8kFho
tJa9bJLFngf/ocPksVTnN4VrLYwwYe85ALzip/eUvatza1knebye/VLZXKL2DqJtWnbjv447pBsa
r6CH2DScdkB+/f59DWgpIPjuFi8TyXU3KjnrfobCQz+kmm/bsHoXfT6ClPspY/BtHTh90W83LnNi
tmdVx1nMYeHCr3cH4Tspx6Ga0acZg3OzW99TGHr2CGDihglqg0ibsDth8TRjgID8/aWCy7PzNiaM
j1PvovmszY0WowNp+mlIl4oWC9h4FSViwDSkjtcGVAJKDrqIghdlmQo3Tp0zTGv+2oU/UEH1snNz
QzIpnKNNtnHwY/RJU34RLNdGriNVJmd4fwsFTeG5lEalJsiMYF9xQ5GmegwcrIafE/9asxghSdjw
lmxNlJPydyNkN3kZ5jUCA4CsXjD0EmhyQaK8zf4ZEiaeno0XsxhMbhKqWKLVQLJE4D7Fr1mazXhu
ViGPmUPiTp5qM00rfQTayWkjkZxAJ3GeRMsbTgD23C9YlWZ1gfCVEST9fIX8BYdOjQES4UC1PUr0
Vf6i1QEw22QImavb08/+Z35SOvszgfuIpXN4DCxgRKYcNEX24lUeG6+xA4B58TqsmvYhQGBAIZ8T
l4wWLe/cSkmzBRopPdFLVfiX0WIZdI25YSFQEOgOl0O5D25QVgq7cdocoDVj13jOBEjFeXIZvcph
tMUnm6LqKATbuSC4+yKNsBJM5PCHAOKjDJ1oEoz8hVzUAJ/a2R84Tk5a45FE8wNgN6j68eBRRDjr
JfpEFQ1Ry61Klod4c6b1r/nkEHRIPbUP3e5mTTOcDB+o7RU0fSNA0Y8phNDrZFm3D644Fsno0fpi
j3Ofqz7B81OZHAVWeclgrYx94xcLqjQgHBr8WdEROfmA4LUpKiWCi8LZGggeH20l3AsGZ+9RmBFm
1GwshyalbfCS2IZ7w2b6aXbg4v7c47IW2tcgVl3LznwpYhrZQkx1mVYtnLuhjk5GvurrpreRNQfr
a8Yd4P06Uhrps/6iC4x+CSXG8kLW7Uz5O7DirI+VNMgNSlr10jvMapWemxwRTZ9w1IvGhSAV3tv6
73wD52kI15z/SeJXSI9GHv/GGdPV8r5Hr2Gl8Z2YrhyFcvy4BYF/nTz98E8hZJQuAlpZCRRqMqFB
2Z3yyZ9SdDLcR9nH4J4MlpIkKwmYkCpF75wpP5/tNL7/K8m+hj46r/kF3ulvWtwapj9hs0tDAqyG
xNIh7sowTuIU8on4sOJfDaoddzruUo589P8+7hmd2AZGYpLwxDCaEP/3p268Hs2b2cEa/e7zGH+c
cl1y+H+7BmQncL54ApBMeLmUwoDDBhqmQ9Gc1hKFag92PSkv3u1ZFDqwIwf1TEB5yS1UomRT5c0D
ZajSGzqXW0JOp3ZVKkEqWRJZjjSDMA99b8pMebwt83qs+oz2Db/lO3QQ3R9yP6rjzn+Oz7YJ9bN7
5Maka7D/RQkSQth3aYaZiQ/kJGt7qPZY9PY6NE0Mf/A9MLTNpFumngRyYgFiPAPmDKOwwCXqd/g0
4DnYB3D3leUtWiFW1jlq53/z7UrD9v34NxgCJdVHOeMuRu8gqo3D6N4hZ+AEtQumy7fcwNg24XLu
JFfHfCFrepAIcZLXe0EzfnOYSrCsBa6SWTANzBvE0RnEEEDUPPztyG+jOL7cFP1Z4BgwnS0rsmMW
ALVX8C54HBaMA7A70pr37fOCjOTtnuGXnBN4SpqZt7WurICcGzJ03b50GrBzHdTFOtqO2swlvvRl
5tKM7OHV3K0ycMZd2YIJZXIMjLBSEWd/ka7R6jIZ0Lf944GRjVeBLoZ+qoWq26UTGXN96EnQnhdB
rL/NUPVn4x00VIiI3NMLOECdD4gH9h/rKKtRJ3CoZupS7WSpIMCrXjaYHivtSscPva4K7Dv+Ie4z
eW0mPUsbBNlZNR0D96jCEO762kEYWpLPE2lbSyIje+Nj+Y4sLKzr7f2zz3BWPLpLaO19ciSg3Hmo
EOBxkaxzJqMVP/SA/ipqki9w5gBP281elWJkBLPlIGFLxJOaeRD9sA/VTZxcpAnGTdMyJWc8ldvF
qPgxTKYs80vZ+I6/HVnrd8NMBD4zhMzkKKIVLLgdcmhiKV0p++o733EgmFi3ElGplUwZJQLySXUD
Tq5EGUNJiigvsVxgBUrDWTDiF6lepqPjGYYuRcYLvmNPKBea81EUnFB90cr7gsWbQEUWWct54fYb
65XCuagj1eaIGip6UFzAXUTUmj2+B64jx8L0P12YsxKWgTiQeQfWDwxc2f7CQm9U9qOE2PasbEV2
+eaqRwt2nK7QXdsRAnIyh6brXnORfFSbXxMZQIdm/t/YNilmdgNKxPcXE46nIXytTpfVnM02Dl+e
77lWfUA2UCvqq1HmGv70ST6OT9Wj4d2e6y1M4ONhtP3tauKO8dPwoKYBFEnqcmKDDU1Y5FJz4IvC
zKV6+DcuRiuisQ8z3LIRxho4d6Co2cfQSYslpWfPU3mIwFc02Ev0n7uW6Moa1KZ4Oe1dB9JH5FCC
F0euVP+GkcVsmSubOhWR7QSmn41jKJUr5VH3MbkAOmhGPJN6Nh4tFgQxcJGGnVyiI6InW6nGpZA6
i8sd183Ti5QPkmsN5hHZOa+XTjrI7Y1lqjLE7W6Fv8z1tPurxBm3QlBtEU2SLTHsMfZ+SRyEOwPI
oTKqndRZAFLZ2E+My5P84ynYxUjey3L4i6EtrT+os7a4kP9nVUN+K/NVN8dbucYf24R1P7yj6FCN
/CagZn1j8TmYVkF51j8nlO8ad9toBVLzm+Bwiva4xQll0lMvT72wHXjs3/2nrrDgvAliVDU9rR4o
fsxHxEioD/SdE1LhXQx3SmWNcBIpATB9zXWHGOuDmtlS7fz1ItgtmGUihrdmH4rovGdDxe5yx5Ck
Iq6bvJnOb994qZkl3ANuUS0CKZJqWFqyztNOg1xqeCAMNm2z/jFDyFCCUqn4D65w6qZ6+kAfhRxp
5HoSlT2OGgAJIjaEVgnjMuj6yrECThRjRFUaeHX1ZsJ1ZRpWlz8R+Wexb+QBnNxCu3Hi12LJex1o
eDb+3wKBqQwOmjVOQu/XD+INO7Zhii3sevl5suHZjVuGGcyzI6irnbdD6Npk+FPt4q5RW8NnsEBg
uud4okdE+pRsLa0xqsDwdv4DOBD7aDreEKkmI0oMUvDlVYg7DVxjUmCmHx8eYVZ3xURSXlAdURBP
lzpvKbl5+0H2uKXOF6aIwZ8r0D2J1fYUpdAencYZzK5aBPMtxarji0gf5XH8yeOSJa/buzleYzuO
trCsJeovralk/NHRnBqMGV2MhnO95BjD0AkDe0cyNm146xa/QVG36kAGi4MWlWy2d6Q6ybTebQZN
8gApMbfRydb48JJElnw9h2fk6YsV0H/i/rxQm/RFJsIIHDm2aoMURGgQzuhf+rXG6NY5padVXT35
XES4CvRG+oOk1102zQhsqwoAgUi9fSMcjOXeJhf38GOGg5z6RDZIM+UVxulfYF9Ir8tMBGNcIki2
Va0Mc+w26ClL/SEP/nM/sPxBOOmOe375lThBS//yzD+ah8qAWq+uaV6w1MxxjqnfJ0cwgNe2dkQk
4blFA57xKk1zy9BrEwq50SpNgoaHqs1/1qVsVV9Ex00CfvrAZ1wtRdVpcF4hnADcEk7gRYOd4VwY
/wMeN6caH/6iJH1qGjY9qPPTHe2bgU1ry4T1xmPIplzyILFqwT6svZd4EbBAfcgbyXRPXOAXMJw7
sxijf65sKljE6nQzeL/QJxqtVX8SnQfy2NjilTBb9UNok24jQDd2vHzTUKwUTuYXxgkF1Qfl+fal
GvuL7CkMe0R46qiYtHhkqWr+Q0Sw9BnywgdQoKc29FizffSzdsnubhGSygicGwGgiEn376fzvPqi
tFPLC6tzwMkjDQXRLxeIQGVnpHmkvW3zZEUwjoNMkNXTg+WP8WKVfXT9LrvUsKwbS5nJv7ueBPDA
gyS/f7E/k6626ZSGWRSVY5dJw9ZqTh4JCOkrX/dpSV3L83k/34cSRTZzc74Wp/uMSKVgTu/ogITR
l3UkwCJ51Gi/o9E3UtsPptv1kVIPTMq9gZ5GNy9MG4HBjgt9nFYdARCXYSwHCVAx9bat1BoF7Ezc
9+qgLgCdAO+PO+8ixtC4IVP06R/Qg2qPC7jAxQ5hSBL6xzP0rM5VMqpcbarc/h6ww/dMNAA9WGbX
OyhLJNIen4xC0JajA7rxGcAxB85YhYusIGa8xYxZdK2QtVEgFXbVJSh06otVueY/d2dkjDn4xYAq
giDpZPnv8vSsGKf4uYgiFIf85oIc22qi125Dqv6N6XGITbWvP8xxV2aXouLPv/aO2+5Yyueoggz9
WIMpjD3+KVl+47hRNZsQWwK22+6x+Rbew2VMczOnacyS8WcWPBOpDtm52FqJGv8u7GLsprnjA/PT
xbacjkE4YA8wAnEw8uI5M1LSLueQXjLgtAWKj1Z2jY7LtOAG26ksnHYARxi2Luo2fLZu3F3l/SpR
yt+pbGCIUXcwVPnnz+K91Su0KhCQsNaiLeThefEhnHIIm9+RUOZAMizu/CMqRFzAowTCSurTE7BO
Vy0L2k/HHStecLvebh+EuEbJJJuK2ycKx+/dvBPsqVeJ78rTBpS4UOPXThRDpgo719Kce82eAg50
z4pTaAsJX3QCSFi3ciaIZtEmLzsLSfg7mLeJj9d4ebHozlUiUC5afB1qHtX+/u05yRm6yeQMcbAF
9VmPDtBbh7kvH53zWgsudCsnDG5f7vKPRfZA4Fkx/m+XIiJK6VmLh0HbN4qxWUjrQTNl0/CkHrrI
//neP0uJf/2/Z5WHXj54QLlKJ8X2x/5fNITY6tHTIkJcFRtlERbiD8Y298TQG/oUiY9Byv1ERoDb
Cz8pYuA+0qQqg6kce7s2y0dT/D0uK8WZ3imvnSybTAQdU5NlPekeR6dWfWUDobvK7VWBSTfFv+EB
LGnVOdRSk44g5+nvVjz0/IQ19IML6LzobRHzbqBP5TLQKWt1rrHKzy0Ele7IN2nt6jKg8TO09P5Z
zXN+xLa2b7w2hK/WQwJKa7KAD3UFKKGTl+KUq5iakcuX4DTyFWLsTfbr1dslKegVN32BdeH6QvwB
ybXvxZCYJKR4Ca9A1nA/6cBvZdI3gJTkZ3p0i1GUuO9Ok4nw0a5zekAeKhmD9MUpwIVHxcyYhxty
zNHnl0JHTMaVNcoRvExUZqKweZbtTRdjpdUZZUFQXTIa6etyz+zL4Z0rXu8hKP/7c9pMwYOHYBaq
mmkFzPN4ptItwbuiqEPQwUsuY6o6TLuhNFIT+X4ktd+4aGZ4kAvz3qhFYnApeME/Tfsyiu1gQwic
VVcPj708X4pdC9EylaFlZwG0k6t9/OU0GJd23YJaDBA8tmUN4eWUyEwEhMpSAsabDp3+gTesVAIA
WEZEtKEu2hUeB/szgbRx8eYSNlzg/I4pMMhk50MRke623PmsjHDmlaXuSwtMhDupChHeZqxn13bi
iJNqPOw0cj4gJu/q0tz5aBNkkCdXDcS9NCY3qNGgRc8Khe2t21LNYNpu7FGo/x+r/U/79h8Ngd9Q
w1LZo1NXtHhIXkreFEtosnwBgE9Pg4jpTROZadhxVkJVVWwUuRyAjqxzyEgjkvl1tZXoV4BpHi2h
yG42pFNAnLF+8Htej/8tkyEGD7tA4qQ4BeIIgmiG6GYl39mJJDBHi04uB57VprDABXb1B6ZN5mLv
u0+iW8+TdCe69R3S5T8QYxc2hMwFA1hWijMpU73m8vukNTXZpfZEmrs32APj2o3XE0I40aIBcQTk
Jh8oe9G8WqRVQxCds1dFCe+WvoJljM7To7aBOxxPaKl8YxfRxZKha02P5d0iQTdEGN9QHhn3NwO+
WpiHbOJ60fTpj7qcWTGwubXBxqjWm+HjoPmkhIvY2LkUqqsJ2vde2pNoUILOpZPeNA/LF8BMFbCu
xMWbrqyn+H8Zwh7RS2cddc75pQHrXn7RDgx5vyGXntbfCSMZsDaI7pMLNcOy8hrmNHHeszcEo8h7
MT/JfWQU6m/bu+TVXYcQfFQ7qqbzupVtRmsXD3bjmfb2+ptb+hU4oyuwC96+bU/UQhhd97173OaX
vbNWdNAd3FToHdEZsE6/eBARauKGz+6wFfkRiEtIHZLtBxWMY2FUYdDdAq5igeOfGfU8EtHiRaWz
dQeGrZ/PI1/vCvZpiQ7QrQ3EaU+fRLBApmIh9dpEJqhdNxr44FF3BYr9imkB7W83EWFFm6IyuiSS
PXIn3abtNINy+LJbAE5PNRbGZ5iY512jf1wFHBtEy6qyvOESDJPGFdHsrMwvi1d1Z5Yy88KaJDo+
FnlO7N7jQsjSGIlc4BP6LJeHarPf1OCDhhawJ2i2P3dYzgpfcogFPbOfrEeMIBHBW1FY24wv11OA
F6lzqglgr7YBllqd4UB1aiFGTxg3HOhci7KqF6QzEZWgkGXztNg5dSqCzhnlc2cRbkB0eW5eWvDj
xB0tJSHFRjLUKczs6I9IOml0SgLapBhj8ZgYmw414mCmT0mptD/epFMIeL6d7roDnuEmEfNg/1aR
lhQFrH2Fftytcr9iMxuaFseVe2VbDgWJEfmjGAxmazzoKedaniFNvJOb2t35ctAY/6g/FlgjNr3N
y/Hvo3KU/vNnmBfTgmnd7Z64QOeJd+rHx4lg8L9Ny34eeRYDubcvR/qrnGRMyqe88vt5l1BhEARw
I18oOBENEHQihqJvGm/AlSoiAj1T05H8J0bZrdDdpkI0bDmosR0B4Qw5oS67vJxjwOls9nNt1gFU
z7o1XH34551lqTe0eKhEdXwsT/u5MPMkimYEXaXR0N0cq4n2E50gQV+ZwbsThybB+/6TT//bbr/B
Cb7HKmrfZqE88J/nwyG4LgR0gq+cM77LsVZyrkE7NMen5VRo8Mctfr/Bml5JygkLsFkp+WDsO1g2
WFq/dzAGimPNhgopw0hx+u4pa8dIoVjIf3mB8NY4g6Ne/D5mSNwynn8B+n69ed/yyVPvxwlGKAVs
Mp0g2z+7ziEt4reLZPOpqqcb8zasr8x6rdsAeGJw+OLRqEMppP5MBxMw7JeTEd28HHTWArXxijew
hnLmaU+hHSOiMnubG1FmLcSD2PKAz0j1v54dHAop8xjLUGzZ3YNqtIsZ4l3aQ02cKlXbtI6CacKe
lfmKJ/B0qeqXNq8eg1aD+rZYJAhOLvVWhCkZjEczPwZGZWv59R2vLIRzwFKkWLsRn+BDwt62XIGv
G+PE6WK1gsEkGnqlIAhZRuozVRY4vG9Om96jtbp6+i1FWLbijy1S5mchvYR7IBJjhezE2AfLO0SL
UunJluv1wXDRZGMl+u9qcpL6zxEcvtfo/aH4fFY1H8UbuWFAG7Y/GW6CbQIhuVEl5Pbq2695vuTB
0BII3O42kcoLWybxsq/RVNWsPjcwVaKvjS8AuR8ofeAvF3iIuvG8ifS2mPupxxA4DsL9NhfXHJ+v
Ibl/6duTrSet7qLbytASEo+hseaDTcNTHYGYxJfvIAJoJ2pQv4hovXEt3irEZbaO9WAi6rxBrQt2
WQCYU/ijia+13MqtzQNjaH7MQuJ+r/GGaUG7kjGkeoerz21aW9gRVS7av4khjRlWpDq+GBIyqXHD
CHifwWdPEyrSKTv4OJz8UM5Kb+0+VRgXcLGXSrYK3PjhttSdDmYoPLX3SnMmjNrdntTtxbV80XRb
xDhPFzHs5CoT2YOtJb9aihshc6HlEM+/r+W4ZIE+QllYxU5u2MUKXzOqVuzpzAwQfhAw8wUGucbL
grBcv+0tlkmIV4haz9hOLBZVa0Ehef3autkKfS1zXTGtGy5vadNdhvXC1hWSZwzOUJ0bru46yCby
vc8cweAmAOVJjn1z4uBclrRdOk0JSnvc/gtydRQ3ZK2TB/EqjJx8QIpVdhbsaRnCYeSKBneF0RX8
DfnkW8S4BNzmlOHhm0rjxhLGJ40zCio9zu51riuLGlq4TUHkBsZsMfUKom601gLF5rjgVS/rlhYU
u0tVc9EET1xqHB/7ZHAFVtifbI6iM9FtKId0Uzf53+FAEmyNSWO6HByAfrIx45tTrkx8Jn/7Mgip
xqhGpciDXsd7e36b2E04oKeAYTAgBYu6w4Frg54v0LPH4QJBu6+gPcpwH+n9LB0NTfmOVKZhvjxS
IgCmf/P+8n5mQe9BXfSqzQ6IYKEAbzgZCYSvFCfureoJXzr95iFIHl2EI2PbDIB1010ZAQ/vieer
tBno34y5/v4xUd5p19Ja9T5HfNVGOQVcXGbNiIlUpzY1Cs652xFaBrIVP02UqNRG3zpYTzZhGHzy
C4QpWkuS9C65WwYXy8PNdz+JtsfWiAJJhCqbW2nlOL+g6aAAhMvMvnE1I6vrm8/6kDhOxTuPA37a
3TEEYfxA45ruoXv9aOdUQEADYLnHQlePMYKrh5LHW96MtpW+yjgTrAy6pF09OCKVEbIH5mM2V02c
t84loDiNAuLrkfgrSjY3j4HP991cOyam7OLDM3y8q+3qLLp71UqlO90HKLOc3lJqDxlqKgpqN3xZ
YA+5Vp4u1qBS9hUaCT2LDxd3Ey1KcsLPvPkXD91hbnH7yRkL5XaF+wPVtMuKD8Fd91+UI8StdoUM
KoR1LELFch9wI822x+uIOEBXQ+t+8FsShRc/hFQvnYS4LDxGkHKGGI38zqFldHN0RAXqe6QwQMqZ
e5pKsG2zzv8Ju+07DWdLLv4cCcArbuZv+zx9nF/mdCHvZla5tOlRpbus6/F92KndazP6QEYhWofD
1yU4vTyH1Az07ewCM1QwzrQD+fJBaZJcjx2JmtNWn0kkBJR8NLHwDiBY0zN6TtMEhKCuc8xAX0ul
RvqHFlTb8qK802bfPUsWq/htODJthb/2wvShezgjVPXW3v0gjj60hsOUKZ4ai0K+rTxjFkUSbGwu
V68Y2haJmf4qfc1Q5JxlC3BmNYF4BxmE0SGLy6j1qBvInzQ6bK+zHi44EjJrlX/YZwhTHUjm0xAm
iKJrPD6T5fccEh/dgGN1uEu+qxACqgIdwL16qRlVKU6JlGHjl8EY4nfge8ISA89jy8/ojlJ/75B7
DdmdhdqwDpCKMm+aAyJEzrPcwDXK7aQv8nIig4/G6oqM30w+YuUN2dxmSrRAfNTaBhGMkFVgAeas
K8T7f4+m1STpqMhoqtSVRNMAUk/lY/6Omi3bmnaKakfL1dSjniePBCbQuxa3aNoNeK4VmtKtrHUf
OQm7D35OjIcNr/BjBT+cLmkKkFepHUeIJj2OTvvnLysaUO0RmoHAZDULK/xGqveBFx60tKKq2JHK
VQylgU1cEVeAHwQiIhdCCa1ZvqLllRwWeffOAZ6L3FZ929zrcO/2kRIM4+zBA2DcpkLaGjTUV3AG
JbJpJpeHDpz9S7E6SiOWYFzqMi0AoYYtzx00PQbPFP/SGpKeCJI2NQR6wrvX7E2V+r4iSYmuTaGz
730LUMZAoSJNOx3jdINObHaxpnG7SZDSk97IyuzfVGg+5ryynUbv9XDwsZSDUH/asR1tBi7EuGYu
CgNGoBWWxmw+x9skpUbH3sE5h+J7TS2l2Ge/MeytsruJBCVq0mw726al7j1tm+Uxtsqk0PbTVkJj
ACgD/5FqWQqMi/CY50dUcrcwNNRxSSB66x8l+8oD88tVE1w+/N7WSatHASQ6ZvCw3EsiurPkd3aQ
WKT+5cK6fES+ddLkn23TWesR+wK57qu9qXAXhn7W2feDqyy8hMYr5+Jv5IeHybqgP84laZusGdhU
urwNHQVTx49vumpcCh6pZf3NTgWVTU2DdcH/59smuqwZPtrRg8O6SUUOOmz0mTaQuxUlOn5I/ZAy
F68VAN16ndltetq1TszJ33lXjI71EGKy0KsJFs2sdbZmynChhNC6SfEGzEFxKhKtDcEbmNFRnFsU
yyZzWUyp9mTSblbLhY5l5s+NBIUEdVBCL8kjyDdsAv5locVF1Wcj6PJ2t9npvrkRxIeouDQAbN16
3JGt/6U/dP7Vl0CrOOF7zznS7hncVcNWcYGD8l1mtGG1G9y2S770m9EUiU0qKIX3CAWoDjWO1hMF
eZmQ3N3ZVBit38b+jVETk0mMJi2PBQ9bF0TxZsl5uOCtnRo001NCT2zxCa7luToRfrez4F9AWxgy
LT+QVmkQjklCNrVdEyXkYaE44zLX95FKR7d9fj1uAs/M0QDG09yKkPGhdylataKjy0y99wtMgCo9
ocWtcyeHUhc5LC9SwoLsPW7NyqgSFmh4QqjxlRtOgcLWgja7Qu4BvxQytbbOTYKi4ZxERwA7uTXj
Yk0qq6Ie6iS/DjgQWUZoiymwVagH9Qu4DSXvCMyF8CDo7AJtNVzADr7inrgnh8cxwH/rGyHS1lqN
PwoBRE40jvXJJU9k+63bsV5blosSjl8To72iE2HCXTTf6VLwu9wJ2n3P19l9NpTHKcrqSmRj628g
G98/ZAl0xy16oxvIDubQI16//rc6Lx430uqnYo2J0SThpp58b7GqW1bI+scV3LhjNPwU4U+laqqw
6sjwewzF1aA/mZJgrrBrAWeDq2DWVTqvEgyB958JoIuSAzFCfhsqLR2vmkjolHMffNoH8WHPkROv
QZiLxkg+Pk2ANE6vpZFCsQzIpRePDYTwDqbS5hGwhz58PjmEkI9f8gv4DKgXfZ2YfNorY814HA1W
jPJ2Gr5qYrNelogjXbP0CIQKfFeQIFzKGitdRWfR5rtWixefOWyjGyTyhy3yXEXYPCmStxqkfArj
aiIWsKQSNcFi/Hs9hJ2dl4/3VxdikFycOJWmbT84wFj0eej1E+NjH8fyBbdKkRk38s8QdhTPx1ud
zdH/JYIUZ1xn8Yv2jesJnFU+udddZEoygeHLlSV3mFIrgAgQlKgNWbQNNKjEe+80AGszohz8q7af
2GEFvS9hNGq1JWb2mYkxEvHr7cZwDPwOIctevWyKoxxme51IxiT1QLP/2/JysmbtQXA3P0y6rtu3
rr1WYgVOcU8XmNc0Jmk09l1N6RTAiBKJJcOsmfMVk5ha2iicTSxlFnogfRndoNghDdWTGtyezBkP
PooHpXAcdS0e6D+UhLopSRkLkHsMDzJOxmcoQBnzkD8GMJumiGBEv4jS8Mc/1sGsIT7n/dJP7l+n
L2cL2LO+4dsW8aeC8eJ0HZtuQxDope0ndaFqlWn1ATqZTqEvZH7/PxJxXd9Te6M8eBG0n/idWFx4
kX5WRm/NRPKxMBHE/b3owJh2lLaEj2EUXDDHiKe0ZLiJ/CFFbmX/Ktk34xQwIQPH8i1I/ZiZa6cl
Lavtq06UCa8E3zeInJ3Quj6re/duyPjL8WbtPEJYfB/GMikkzyNLi9KyX2Q6xnVnVP+BC8hFO6ix
EyAd8jQ6bpcONwiC3bQZ421R93Z1fb4uHobEtbGWCnlPa/fPoX7ILAjPdcA5Ve0Fy3w2E0GdbQar
Yc2PksqMxocDkvYb1X46i8iVO5a5uaBsfVbT0KTqiu9k17fACBJAUuPNBdQSDaqO6PvANKQbu58d
bDJWJfGSD3WEqhDtO9DKgGc5QqLBetxs6Eyvz1ztPiCbbWaIftrRmk5SL04e5ph5W+dRuiosE5Iw
ZVcgxgXp03QAqd2Bu30Z0YCRNtZfEG9buyJb6ZgubRiWBQBT0ogSjTjPzeFwmcSbetB9VYkVHwGK
E78jJHyN0UqL8O+fZbGhc650j1SHKAetqAtrQdrwIHHZLzS3QQRf+SY/7hx6nuZLfFm061sVYbMk
qOmn5/fwCUp45GuxCmuRTOWESF9Mcy1AmN6LfJaTeDZNgPc6u8Pib1GaKCmyJgXpiewFfnm+qmBM
B6SYY9Uukkz+pvqOSYmu/j7yPKMaXZLqbN33Ad03UMLFc9xdFQpa/n5NOSFOEV+7Kyzz485fkp9B
rXE2UeCZMd/YWz38TqbcFZj6TX1Mhtyng+cRE3FkPtOXMmW0/kCq+Fddfx1fgMNruuQ+vE1efC14
BAJI1m8EPuLZMB8Kvo3lF91ZyMTxwlwwdalBizUSgeRvbABbBJ6ZLaClaWgrRkfn+xJwFNyDlS3K
unAeE/FoEfcT1IBX+fw69fxW1QXEodfhpfZH4uoQnQA20erEIPHF7ttEWmWDMH5pWxHCQygVDBZX
TzMYOg0SYDwew13S3sxJnsk5SuGjs9j1iKJEOlk7abEI1yVcR8qRuqBp+QBI4V4Y7vm54RowYton
6A3sizMT5N9osDipohgoAgREfb/kCj2+Ud3+jnVdH0ILvdnrqdkJ4EAdFVDq18VzJ+EybhM+1AFR
eSomnj96LFgh2tAhovi057s3p3ySN0NKYK1vEBERgm6iTFwZZWnKn7ma8n6XlzyaN62KCc2iqy2F
06gj2qmvBtLDFHEwotRX4Hkz/swCz/s2CXJzKTQInr3T81nzosoh5Olj0+sOMWwcDxvQX6I2qk6Y
13ErgMFrw7lNycp5WlymzCAR8IFdhSfdAbrgh4MjDlL9eupAniBFysrcfxIx8tDaH8G9DclYeCW3
760X8MR+X3o5+0Sd6n8G93kbB36/fgrcoeOu4ot2enEMRjfX+jQZzBZOXCNJ9fjlrlf0Qak2C9Bv
CLIPz67kmaCTuk8DMs9STzhqonOxxDnhEmdART138EU/f50ZbxPLz6F5yRTsjo+NKUSz3G8uUvW0
hlceQIScCzH6HIWpnEIS0j05DeziPFg+C1uWiv/BeVG3i8yAPXFTDrHK9sTkUUWYI7+6MMvbuJsi
T9Z3AhsM1dabRYFo7na2pX/yErus8XEkngUAi0joL9EoC/YJRxswYf3k7aeTSXuWJKTZ3vm/RSC2
Rydkbx3oyXvYr1sN3rTjcTPcsLPEXRtyE/1ZesmxywnNlBLJYFNce/Q+kLUhvV8bwGefDTPjbNDz
DbbzTaEsG4ipGFFcMuXALWgil5gkQqutvadaZtsRHyzy9mmhYR3vBLe/0ClgqohSWHhhK4/5qcVO
q/9RVw3mGD/m1EaU+QW3SWIUF2Zw7AoINEreEtvKrolOfTZX4NvtC/67wiD0v8JAkNC/4ZBFt8Wm
dJzZsUXRo+alnTYkF3eYSx7kRfHcqA/R5DBIaA5o8XpprRaxhdZfrcyeDhcvJLmCz5j0cdJH8aPW
7poAz1tTmm0oHY3Cwa0MZNhG0hu5XYJKawupg6M3H25G3ad7owTYNgO5RxM8mnCaM7EIRMl7gCqu
jM0l8JnMIdyiqgwdpYNh63GsftlUtivmjagBeC35Om45EfsjSgBtLHQvGapIc3QWXyckc8Zqniym
jgIpY+/EE0BR4+lWublfNZFI4G+l7R9KHiEtpoPIDdgNSRpw1+AcqJztd1IUffwZxYVklrfgEUW/
BSLaBpdrUkDrReLzH0QM1M/NbCVOvktNqUE8Y1CNu4HBnAuciGmhIXgNNgEx1lLIHuQoDwH9L/MZ
woApydXoApMGkNVCDY2LtwTHgvQ9y51lds3PNxZ8AvWdrEZnlQoHPEw2p8NhBce+hAqyNc3taTSn
FXuMEeBoeZPqW782uAlsI5JbyiwMJlE7+SKxURiQPxQp5c5OKhm35dRWGmbCF319BnAyzRHr3nRk
DGaYLE00IPm9eozhl+Tw9YY4g0XTLh3PhKYlJbR/Hmno5HCmzNiTbXbQ5sAMpBg+AOhayU0xPABZ
h+S+S8gRec77EFOtfXbtAiTfeJLUG9b6glPfFrSdz8YJMnMUmUDOcdVrWbdpwlmQmqwRvpSHdANM
RuaAnPDHez44ABluxksN9P6JiUlolSzlaloBFYiex+BCPONGgmIotyOL1P7xzECq9kliJIUVIcP8
U1jwGrhOqiiTnwRkA9SN0H6Nzp/UjOyo1i4f7Uix3HtGRb3tQv3c1yvhtGt8bPAWch/i0j6vHPj8
/Hab2VO4FoPqgJsY1DAnkpyqJdTO+qpRI8YXbmTC/IOFFFqnonQ7AeqnqLRi2B0ERcnEicv10WTH
iCqPuSfJFWIMRvXs+GLSe6oGuihfPRYyOXOsDh/a4/eAcoCMmHfduJ/HB3ChkScdZUIVLfB+sn2/
qGAW4WUvwNsAKKx97RjN5KoA5uSw/b0HtZvNTZURcBY6igjnKc8lXruAn8xmlfcZmvmPc/phwqo2
aPW8Siktg/S3Viro2Ref6IBmW4Vo+vkPt+ofCyQp2nzo99mlNKspQsRF1BNiX4CziE1xVa2f2E8k
sBctV2n/lc20BUgmC6PiuN+Yucm5DLxWrE1fmV6YXVPsheVTf/CXgiImzhs2g74ouxz26KodxW5O
NOCHdZ3xt8m2VWgKHtc6UgS84hQQQX+nDr1aeFeWA0CVTYjANQD8uRBUSi2ABsKlBsopJU7/KFPZ
h3menBL6rginHJlzErUcm5/I57eFuwnXWyK2dVsuPbrXhLlUg1vSUnY/frUIyd+cXv0uKwZNXYtu
iNXVxwMXOvFp35BAv3I7ELsFONNP6P1BBc2lVLm8YhqwzXp2MSuKXiqcJgiY3u3SxNQlGNMuc0A/
9+qnVgZifS4swmAWgSyTSoxI7JVTCeky5f/2bMfxV5rjEfj8xaA5fW6eahFnyzun49qFlFpI1kNy
3/6fYdvnrWWxsWWzm83RCk7P4KAQX7psqPeo5GM7mJQey87fBvPmBVYAktmaIVAwrWxE8urXp27X
0Q7/+VI0nJ6J/nzh7RQ22bXfyvmo6rK0cN/ZNnixlD4l8MWWVzqmOb/Y/sueagZ9nNLIujco5pNH
5GiMzN5vehz1qwqP1s84zcPDlsPp6vLrsjNM+viilGhUBCVChOigaD2Dj3nncLxfrscTQTj0TlZJ
1D4fLBm2nWYuI+UHLfhqiBHCKZhERKx8Vf/CNLNH5g/1pABdWVT0C301bokDmpen5mnX6yrRNDBh
4NcKOl3UWF6Zg5mipMePBet5DvEYq1cWO8OfH+nizISheLnBmJIZiwKxMYX1QYXwo1SVidaPt6L3
eYUKkUNrPwBnJXImB37QRabubdd7hYCNKvXOPhcaLFzdKxp0z+ByZuZCf5DpOmuW+EpdE4t9EQ3r
M1ryy0I/zZkuYP+mQA7chpEz2fKGvULX9l8+uoJbQdwPvCGr+Qug7g4py4xQEDYhjpGVo4curYsB
HjTusBrwOw2On7c0hYYIBSWmbiCQKtooFJRoUHvhwOXzagZQm5qKMzz4w7CZ2gnUDxvEHx3nbV18
vS9vE7LRuVHyxlKo6iAGQWwgP9qCnEyiIl3B2gedauDDgAY2MAHeaFqv84G6duP0O8b00NINEUwB
jyydXGQD1pHgK6OXYTvJP28AxNJFMDrh2gKpUhoVMBpTG5xIqX5mb5qXBjpkBCaFTRWtBsOAH/k2
k24vwyqDUkwtOylKHC5Uvcg/9coUFdwfDfbqP0oo30UwcVNvB7+2WDISDAbko8yKo8igfUg6T4Qx
SqXbzFzVI1trDNw/BZ97sw7/7pukTQmdp9+Unpleci1ezyENZv35Hx3dgtpLh9dJd+Un9fg3Az/F
7/cnA1s/1Vr8ACiv39pxUNrAf6oBwRqcv0ihHfrimDudxSeDC4RE6Qyk+OWY2XUyumqDndqSbYOY
E3GMtE+rg7S0hUFENf60FgwaFDYT20fW2MQ/L5zZWj3QVJeuJS16WY63vnrfTcv03v3YlkZGDTet
xe914Oa2BB2Q33+GeJM6cEiYS4TuoAjhAaMosjrRHfshxMamQrlEEgmj5CR+U27Gy+ujWLPNcKbd
9x78Fay2HuAlFSh5J6WMr9H2QCn7ylowGnRiegiGTgQJoIYLAe6zi92hEpbsOVAB5ilJCu4kVfqj
I5hnCNplUDmeZxRxIGTSckl0B3idlh/kAwsGAElevk4UCLOwr02c6OkapQ3i8VtW4WEWdnylngCb
FQUAYdVgCi3kaAmS3Cde37+xHVRrWiZwwVlX+U9JxI133EIc1tr+jtEEa2wHZzqRbfw7lxkmR5GG
RJpy8JnRdyYp+JTB17QJdwuxs7/Ll33fqWl23jM8qCt6KPWKJdHrg1nl0Guk+BDFHB+Tgynrt2Ov
+aPbDu+my+haokW2VbBmzqNswB6m67XODk605+HQ9E14/AQvF6Vwyl6/S6Rg4avtPoVxGMTvRUd4
dZ6W39TrLqqDHlnvhKTeaC8h8OgQjpYQbTIIsLce5DsLl1UHWPtHcfEt56UmUk8NwiIkR1RLHhsP
jK5z+q79R+NJd8ITeoFLONJjPKcGWtXJL0icU6N2mYD9I7XRC0mf5c6HQU3uZJeYeNYiTgjaUHGu
++jg1ys5/diZOghbT0c/gFKdvdYqahxR5gTdBdKjcS80S+gpkTq6/ZM+w5pe4++npiQFKbZ8jROy
TKESUQB7xC4a7j4yYicQ4kQXcy0D5+FG1xvSvfZZUPzYxhhRTR0QmgoHm0A0/9aZZSAnSpxgIm3d
JZaoW813iYsYtBN3MHC/dbWpl7nP0xVA+Dqp7s4ILYZqlReh8rX4en+Km3PyAZR0vTdV7vhq0bat
AQgHWkAf3MklLQA3Fk7MOEGwuxDIIXHFxl0YGyVnLZPNTeY0h9UIe/9eWc7z9Zr8VS8bI5iHzI5z
BcqE/Krc+4Cr0v9rbS23zfBXACr2KdEDdbC6BzHQt2efPvXp0nos7k/KW0Fjsy6wGVoDgtHCwA/M
pYvA1aPEZ+OWckuhjmWO5X0XA4Emm48d1m45wWTnAigqL4Ko3GYkrjAZ9K/rZySxT2A6SZTJY36U
OZX5chmufwgAP2e2SmqnIemvmJBfTcSM8hoo3gdd17BbwT+p5e69lNQwNdpQMZ2ixwtTLy6Eiseq
2+OxaCJWnFt/9UGXKPYVcwYb2Js/XKsQlhIc6cPgzkCXs7vupviz3QUA211aDF4Wxy5biDnzG8oH
yM5agYpd7T4HX3fm6l3DvgSkyKRssu1AHa/XvWFGpQia8u++PVkL4eEgqDHt6581lG8U28NKuYQF
4j6NoKaZA1akFm1mVAp6XaDyiUu2B2Uw4su9mRB07v7RLJ+gMXlEk+SjWfXYuiENju4u3bVsDAvX
3UFMfRSi//NkBWPAnNmRCnlTpyNQoyOaqCDUuI8UsZDp4pBH+6oq9w4EMgd3E+eHym2PB2uZcp7N
8bhx47MrX++QYcxouM7vipRdxotZMJaWMoL5ixfikR+2TGZG09jEIsVx4KJH8IWa2pA7XDHp6dd8
sRWCEqIXSVISr6GWylRFqzYM6kBQiibFbmXRlNdwZEE/L5pcLc/q+utkvKib8mypG1q7ZxSlztVR
NXYpUSCoZNEkSQ3EGuB1kdTbiZ89Szyc365MomzFA3tN7RGy2zH/PmymLzeupOxjigJKP5YxEl7H
yQXklTMT4CHD9iW7obZNoF19kpSUeuDo/5ZD5/SQTlTWrMd60CJOOivyRv6KKUMxPSOzy2etx31E
b8lYJQV7Rq3cU8r+v7kWMSgScJftBjVo7YCyEWBMOY1tIMZM1A6qdvn/6pr5Xr7KaB8lCCzcyYr8
c+KOLySxCAjWU4Ml8wPoTa02dz4Zi2HH/MOTO0YRadaS3AKrJpbEhUxgnH2r7rnl4OVGYu6ptZ2q
eJe+gjV+w3zXoJ1kEAez0c0tJg99xaC9UH5tkiVb0xl7IKUT1tZDp/bgFe02gcVDMuzYAzRoaxZo
vDmy/4cCM4lUayNUWJYO8ZHUVWVVrhWU9jTwbUIVMEZmrkolC++QRTN3pVs99GKFhp8v0a3xr4Au
NtU5pKa2XS9zL2tMTC3ldUSYT9CfiiW7wkhTmuDjmAwNSyXyZw3ytIj3jJNLV/SI7tMKPJEzicFj
vyPXwZPOvwsEA0eF62I81Ftutwyq1OTwDQH7efZ1Nj+Wk9TN3gsWIr4TfnQM3GL68aRaz9bUgVh+
blyrihEoeuL8A8F0w0qQ/F75c+QfpJMnSrS5VNTKZQ11R4UYgjeh9TFQDBTfo1ZUxDfu0xdi2BX+
sUzWFak/cCqtZtkNwQ1Co1ZJLsfUUAviqs2LsDTe2X+EjhIuo7wDhfV04Kisi2yrJYY/bSL+ods2
w3frwWSKMGtj8+GgUDXkBTT/M0fQRxfadR08Uu4eHrsTyfqCHpw0hYYmemZSq8/hq7xf+bW5lIMO
fk1qBfkA9I0TLDNs6i+LgImR0VpFIinCABRXLuQrYBGbZvth4da2FyAcMuFqKAEMnRBk9Ne5+V2A
nVP78leeq7skXzFKkgAyYWRzwzTLQPL5XQTsQ9Qw+aNS5WzMvri1o4735TuDTCf2cG1dofaJAIXW
qXWveQ5WKHd64c6reNjDwx4vSnkhOFKSQOoZVBUh8b8VGk3LZcFvH513ktqnwuDxue+3oquR//wW
aqqHdEeQURRu+5wELjSEJ7N75SBWqdDWXBvHA/YH0u2t12zG0xySYtdX9wLepvJ8MiecWTJJ+u3g
kvYi+j9dYK0k0qLSG7BlimqYTKBVNcXPnuUN24Dmhu+A/bLE1rO1S8ZT6psYN1xQqzRaBqJMRCrd
iY52s+wLW7ST/Hvj2mSWEcaEqX5zR+Trghoxef+UDefMaENLBVwHG+3vnqRMyzkFv3CzxkzObkkL
J1/n42Y6AlKsNnIKEnuEz2ZLIFp37GdoJWGakQWYi7fH9cFYz01XfBYg29aXxbiZBjkA4x1Ve1m3
lcrlZqh6AYgQw9++ODNcn9JO+ssaULhogfX/j5lehCCkntFwYP4NKVw+rja/GKjnBvGv/x7Gy0sQ
gpL2WuhLIXU6R6Wa21+m1Dq3+ECiIBFLno5SzsIkZe635zch4pPWVOXBdKdcMmvcXTggL5RQdVVo
Csl5Wx744qWZoaO/5H6Vaf7llvu/03I7LsPlc2QfuazP6UJ4ESFU4o/mFektG4uhTmo3Iyc3AHKi
YR/3oiQdHF3JR/nQ7FM0UNB3L9/lZL0DRsddXu3dbW9kVxy7HTLdYLfDsLlPJQQOaUzMAof2cZuW
m+Du+8oXCg15VLLl3kHXzgFa6Qya/VAZZHE2y4ACjGy8ipuRZHvrF/bl7pK5Gbh6XiDK5vx671Bf
wKv8ureUBAeykOthpFBK5v/k0OkwsrqKePu0Pfd9hordQEF2CZXMOL2pWeEl5R+NIgZ8cRTwNWKK
Tj6/KchS3Lx+Tm4pQNR6VeRJ7X/8UOD2dEt5fMCYdUd7x2dEry8OYuNaJr1iEGIGNWEMVAqtCijT
hsa9V36UQOe+UbfsO9omC/L7o4xYQfvfQm8UdXlcnDck1KZa/3SlLUp+zZ4c6YkT6Qt67L9rKlSN
gTlHd9nGmPxejjtisasstTSt33w1Dq53RgZBFW/v7Zqc5rZnM7m3bzJSYkGcF5fewSZKS1na+D3R
npnsmYQ7Uv+mPoNmAJUS/SKwz9rqGj8jMXzqkLDXiYps5zV6mTtsRUGMF35lh3cxA5OLH2p6hYT7
ANPmPw9j3VhgRkK7sLG+eM0hQk/zZkHBmyLoorwqCoN7yDgaPuklfcPU5/02ygBUESFnPzSY9xbe
VLNC2QQOirSxeq1W2QH1Zm4CCzovonHcXs18BrxjTB/E6Kn6yAsGtIgA6W7mYXbuciAgGMDkm2f1
t1XS/ShmEOpDw4ZEqfwqSjXSHaBf2K1H5xTZkchMxCnjUkAYvl5kDnGoHS+0lp4y1HyKPb2qANxN
5TbS/easQWRZvu44DhnkbCeUpipFslSY+j7yTtatabeLTLcUQKc6eCC0M7JVDiZj6oYTjL+Lc/RT
wRahTin27PNhJaK+ZsYCE9b8EErp73Ghj96wNLPbthsE6ItfQPWJgrxuUwTRnzL4uugXLCf1+ONC
bankyzjI2BukL1U6UUnQQZzxAoqy5rXlGC8bdKqsKs00KFLHbBVcZBSUc5PhCekLTPmuB/WpIau+
XQs731Jzjdoeud5nFn70+a9WI0ME4AhHheLp8nPOQQhpv34oZWRLzi9rMnftgsrPGeEcfsinyAbC
t1FTu42NSILzcrOiBDz8iy5SIHNJao6RbAloxa6Ejo/r/yypTN9yQVLlyGaRWxZR2SgK93xqpSxb
ajbk/1cxxJwduSg4dZoTxc4/vYmGQkybwf7JtBOTwNQo1TbLv10eiuQTTehYMEZYBZ6fs9fsALaj
hXm/BwnhVQCG1J4uKpzOke+zJ5Qn83xwuXbSSguyOhINJX3AXw2Pri2DWwQfTCJ5SeXvt2442tg0
E4n3rarXIwUOcyapfV6BmxEKcaf74m1jY7/KCXb60YaOyZAoYmiK36sqph1BjIoMfvn6OEXzZ1Ur
B150Ll7p46RSBuTK0u5wpK+dpbegTi02JSUWgb77UHrmHYhRT6QL6W7itipFuqdEFNgCD8yVxYHk
3bqlAH8hMsXeruov4bOd92+9bTGLEZx62KC6Mt8bvC+klPuHogFi9WsxuJL4xN0MuR6Ff0h4gVHX
3OqMdtRXf96zJI+ZqNlkWGyzlyPQ9qpCKwVhbR6aO/fGHQ2Yr2HtXYyKGHTc92QCS7A2lsv7YhID
N4Z7ep3/1QsFZctTKbp+UNv05GWwplJO36ApRrAroW7eTqDon0AbkfhqOKS6kmgGSllWjSCb9lpb
6+5QKmsg33lwm7Knc7EydjZ1Ik2CgiCwuO9k/tkyQgxVL/N9UFdbXYP7fmojHRhQHg19cb6o29zQ
WESIhm4Ploow9/SU34jFGnoJn9hvIFwmjYs190nWZDufDOrwS4BJXf4Dxh2NNAId2b/wBR0gvNzB
zmUqGPqMSirSSs0WPfDDyp5oOrHMYdJao07pYPM3x1cWBsd245DnwzQZDseLHVQzuE0c8i+WZ3nO
LWKNEY2eYjL6f+s0VMM+5nOz70PFTY1cQ6/iV4UhcdnVvKk2H/Mg+C/jC02nWaJUmE8bkXTv+ArK
Ijybla6OJ8KHzSPD0yZxGxtd0k4IoC/C7L+35Cqe8jYwS0inL8cFblavqF20q/HTlQwU8V+yfIEc
nqkyEmx5gsSv4cKVFWOMjOnF8yJMtTb7I4GUcDgtzwkccVm42DtEWtoK0rWwNCXyOTCZWun+CPHg
9tlWXXCigfD7IsD2jtT2SBMmARkKTTRltVaF+9m6QfkhhLxrld4wY8leyLNdZ/IZsf/Tzmj59BLm
hJiCwDYNM2HECkg+H8Y5lHHikQNMYQruUoP5TafjH4JSKjK+wmcyzh38Z7xMWUNhQuoDhelu+uMC
CGuN2OIxJVkF2xNfXm1P0IkH9uU61gkmxiglbCUuIZ9zscRVYEPJbpb80ZPQiT/aKT0ykyNOMihR
0K0kSCkwO5m973AeQtyhmrVbxfDn1KSv97aHFnD2TUmPT/06Iu/JIxz8swe/bZc50LIsxoTmkSse
GQBuwRV2UWeDKDdPVoiRlcoJo0BVpTuOkj5KxtAazAcaG29ErGeUH72do0Djlum/a2KEq8aURIub
mKbaLD3ugKPWyjupZlhvvAaBbIkUJsGgoD3FjOJngqLa2os/69gJB89uGcuzzMt2orZOgmO2cCfK
zUpsE4Xmz1i/29jaUuOXna5lYMUnDLPc06Vy3Q02UC9Omka0mjLc/Sf+NeIQM1zt9xJYC+/+tccl
WeNjejEMRRlXcy1Ck0vJtQLfH4j8ATrDEgjIIsckusMhMIgvyw+6vC3FwD5w44KSMvn12li1u3BV
QzAT+RLTDlsU41DQm8pLp1tAu6leTnqJqMKB0cvpyjZWB89KRVWFUA5m+9348AlmxfWoeT7lpqHw
FczhEnG1iDEx+Re6G2SY8DCtDu8iD2JAJm00Xb3AJ2PaAxHQ9YumkcdUrk5BaCzb9sYbnijd7rw3
QWKC17iw68DAhaDbxECAeXXByFBTbsk7g8oZLCNde7PsCPJqWpjvOfgKngz4Ykl+RIaYKU70fOfm
rYIb6YrGKX8RLxymd8qGwnAgP8f2WhFmbtR7YpafiKDCREt0h7htr+/Qcq72bddwngwpv9pyZn3G
gXcbm/L0Jfe/Tfyj+zmDwibm4NcP5mxfkWxkFQbadvQtYzzdE7/bKI4tkdYQA5poYSDDUryqGYK4
IOilJONnZRUOvZ4FyoVLSdkuJ03swxpo4HUJLzUBAj3TYVKkOkOrz7jfXoVb4yilKKyRl48jA6to
KJ6RoobCwF4eKdJeUHxETpAGhxx4uKa0xn2fzFRDlaXosYvKagJdx5Le3QD3FMSzGlWEMbqGmPKY
pkj1n5qt4RcOoYy5eHJpUDWkrPjvFAX/17hue/j+/FO6EW31Ri7jPGDDiuqaDk8nuWek5vXJKtzP
ZD3YFk7T5Zcwq/KIguouxGXhI40QPB9TcxTKdBm1q8RvOVZtta+cNoRKoOZiLGVmbV61o6GoNlIw
FoO+jm6Nx/qbqulSNyQcYf7ntfyDiUSVxRYuEfFfNvCiHEVY+EXVVsTLLHjsWUYJPcwth8WUr1dP
/fBY2g7XZLUrvk9AIRNRQm9USlga+OBjPRcaHbqBIrbtJecsf+e9QnjkRLzFlzYrpwtVbHWKlPOa
NseCxW9ohtduLzK7WwJDmNHTGGMeO5KfCk01ozLCzy4O7X3oXEXfL1G6mkt/JXRa0feGWlfjDOAV
yt0WBsemc3pmuzEXRcpVO3sLwQ57SpRjuOnn8/F3Dui4zkAkgKb6AMJSiL8w8wrCjmXHTZwtUkiV
Nowdlr4m8PzK3+hV3vQ08FlSrKBl+ph8KnKbLcytBxtoTZXNKxItMbDkNBYU+OG+2oO4j2RswCeU
SP2y+PErij8T08EAqiLGLTTz/039aNeyUXItA2SE2SKB7ya/ODCArx3g4LEMRlAYpZcC8cori6Gy
fudVUPSkGKQkjeWyDZeFMnphqRNFVXEx2tytibCttVMXDqofcjd+O/11jOVOK5x/7ro8wHq64reD
1n5x1x7Hna4CbmU1CojXTHNzwfzdA4i4SbIWY+s1pI09ou+JSZahqUW6pdw6iqFd2TgID0y4P4cB
lHRXKvZYx3af0mNkjicsB1hXv8fYFblwW8XYlF7y70IJbn6JKSKjanT8gg0LR2qDqNF40IQx4f8O
y1PlYGZDAyfkXv+OO/3l51623hOtvdhHRLyHid8mKxl4TSGe43zABPFlUgZMGTXA7LasiIq5Vm5u
hXq+YGB4Kd2ze3Man/mI8+L5Z7gFTN3a7TkNiXN5J9q5BcKRCnA5i7hw6zLcH/53lozUdFM7u5cG
sXeqAjpmwoTpcUCLAO5fSxeKvv4RrBMU/RP/ZoEoyl6qi3JTJcxBJQ5XqZUk/+zBzfbeI0yc1whj
3OBmFAV4Oan46gZuH+b0FVcDmGE22yODDEHlhh1iEnRYSgySnGJo/OC7m9ri1sIrxTOHyv8/tHcG
aZC3xd++ulIzTTjhtDZfkibw4rYSsVbmWg854Q52+kLtCjaESIVvH5TbNPzC9KmAqv4QlZDWHGqq
pkpT0Yfkm9NpfY9FCwvr5v2jMntYLiGAKKxMiK1H27/ls8twz4eCg2O+EZCJMEGYAXUfthZj2fGz
durYzBVWDQXtEszAX2ohJUDBSrOoLGsTUfdQk3li46ynxNkE8TK4/lMqYCuQrF/cCL3TU5JPmobT
pXfm+KzCTtUkIMTfntDX3ComjgvtUC2dMrh8d027TkwwA/VOl0HXf/5JbBTsnybkHFj4MWOyXyNz
rofy+rCRusbFU8u/9awMkqSYl8tfq0XEmb/PwjYwDyAoJR9rBTXxIQpp0G2TNdHwTBMH7EsJR0bn
L+EinHBi8cnSzq+casLSvxsY6DXQ6MnN8EHMFz6lNqfMu+ge3hKymvU0YAct/YcocnYfCBPyIXYn
mAEeEkF146CH71qgUoREoWuHm82kULb+0WfY0VlsFKtfg1Kvs/iF2WpsjbTV9w4tF7rBMqkQ39m2
Tq1ea/IpBnAo0xyxQ4kxe+j/2qtQEQ+0Xhd/FMFw0noNLGQm344Tpqob2nrYKrJk545zXxmzUxSr
t4doTA2vkEVCEuCXxmugVZl1Uk0J4WCXUMf06TWlGWfHEQlfqGScq5bemdPQ7s4K8Y0f8Kpl6qQU
mPaTh75p4JmE5sa5zqC/6t7VMU+nxgNoynDANUtsZvGWdlH62GmUxJd9iYN+ws/uG2eHQiv/0fEv
UN1ofu+x+cXg00XxuX0QwXrshkhwDHZwYQvuZRVxuJuGKON+1Hqlnzwj3oduztgLzm6BXPx/PQqw
oMprH02IXKbGl+rTDVwn0ybdEV5CCJ8oakLfeIf/g75p0mtcRPWX+/kSwS2CivfhTDIpYnxXLDXf
FRe7shTtwOvBO32JJ0CzOCjf3ylIqxwtX2RbF7HRLvMW08saJzFv3yCBBd8BuE6B2vm6V5rBbhUf
QiewBZmIu+oDCMVOgjEmL08rLEz8XTv8O3W78hk7Ay+uYeR1PDAa0BTlSY3n+zhlpt3lgwahWhUE
YiTlnsWxvPeRLqBN2FT8HEZBGdjHpDlPuTERT8sRZtHv55W57zFh0hf0jhI2HkkoiCO7bGzerA22
eW08agzlTlh69EbTzXHR9cYJZwnh2iEBlnQlMVYRFu4Arc1Ol8lcYtEaGSseYz7kl9BqbwGwNx6s
MbilK1uGVJi86mcDwc5aE25NVd8jEsRmNqhYti2lmeUMPtVNKPizY9F7Ft+YKBncPc1hUBBf5lhI
TcHL51w15aw3+17f7EU4Z3o+U6DQQW/o49dtMInZXhtzeUiwmmr3vPKR2DSmif8X/L+81EJeWn+I
38/4uBNWXLPTLg39Aj7H2O9Eq/agcfCEOJ0O2I+m4H4CtLYDAS3Agu+dnn/Hl1mf6mHu5QwSsnj7
W8vcMNrS4uJBq8APhqBxFm2ULdR/e4Wohni8h+0EObGPsOyIidwfg7pVUKmkd1LVxW06qhty+lss
qF6WB5sq9M4A3SEduNG5jq6craqdZjnivrHLMFplaTBTEglvoLUeXdq8OWNZUdL5g+YJZMuIeurE
iVlhJ54HKJU7/LTcRlqeRBLfeGh5LG9EI9LwHrglgN2UUKqsOXOgVXNnJy2x3ROHLHz9dXv567fs
cYrHlv6JDfXJA9zEx2z66Pc9T2y3/KExSQGpODwAlT3D6aanB97+t4tTuFq6bsLduNp1QK5VMT9J
1rNs+VfOoOr3lTAJu18wQMAEiFnQuX8VNtLbU/lgttcXdfgbO7Z3qkWrDd0xGrdJBrSv9EvUbiJh
FSZulA/flb/t43FvweP8mI967GtjvDimL4Z0ypzAUn8NUd0JEV41LJameJAhY0pv9k+Km5+QGcBS
JBtu3yibxK8XRVx4Kuv5L15q1/41xGMqoAAZ4B6gdpG8FDMEZR/OMLLj240RcC7BueevJv9FcHo2
2AGmJ93YhiErj6gYiRDBgjEE7ydAyI9ejdt5VzzbCLcL2xX8EjA9YNB2AMAgsYoAgY7z7l3LbJNq
GTmG6pjNyhohuqoR3gc3lF6fqahRMIbecamCNSKS4gm4st6Q+J+nThEX6/KkMyLvHFjg117mnE91
A4ublg3BNQlTDU078IIhJL/UyLq5Pf0u2ikhvFFRmVPjLytUjp3RiKdQd06KpuWMDUnRPYppDmlX
VQrLi+IuCmInPnX1yLlWkGquOLN1YBiY6fx2hl7tSYtR5TlTomuBYEndZbQuMxZW5/zGx474j5LI
xAkU+QLiHz965PbK84ZyEf1YudTbNRF+t71ebsIzclMyEb7WJi9dbk81Q+zAwF5s2y+i0yAtrlKu
f0iNIyEgxgJHdVOjzw1funm10Ty6MQQedThB3/X9rwakL+Fz27ln4Q3eJU9FEr+2jZmvp2zekcIM
cUH8tA4WewUoWVQJvisRsb+4cw6Q5wnf5GZOlgkMMBhWeHAJeLxeWIUvJg35ccY9J/o/HyxBCYMW
UhUEyT3XD5Z5ud2n6a/RbMOGdDHMkCFEdL194Fiek2gUbInu75LGujOsaZQDmAcPPGD2G+ygiaKm
Ln5tDKrt7rdvRPfXRJRK2cu//bBaxse0WZdUH2g5xekTh5p9EsMoYprJadMYuXTEISjlQW0uEJad
Fl1MJFqRB6DVmg1mnr74tlnt9D7c5vqs0qX162IuPSVTkSc9vZm/Ww6rebWuSdqGLBeY0KOJUjWH
ZAI3MM6VICzkaDmc28V3Mx2WtGJ8Md6Pqv/T0Ewu4R+22K50popuaLpj1MObm/v2JBr302OZnh1p
Jas005fmsQefXrpTLz+JNPUU2VHiIWSwjbmRbijVwSLtedNP2neUIibwnRoOPSB8oUzFuyh7RTBF
jzJVBCmFdpVa1ntSLuqTboScwJ3A5q/7hTy9sKdYnncoMDBJ78kdZaqTpISj5fuSFpfjxycraM2d
EGPd5F0SY2qJQpAB+DgYFQswKJmn50ee3Zv0d+L7iY+um+xSJ9TGQNotXq6tNhBnRbF+DS4GKuC2
7KkHptHvVuB4+HLkgQH/RHGZ8UGZWMiCcjaVtXqg8aaTYPiFZgbISny9Qssag8zb/Tl2Sr9EOhZt
qzZ2P4JjUj3sGiuExQtQLwAAdgXmRLx8eLJ1FFTLfn1TS68JNZBbRmMwXPbAP0avs/pWPPIp4t8/
58e89V9WBbitKDDzhryKwJ0cLgzJJog52VNz3ozUcKTqtRZPLys5y/m1K8h9pKz2WhzDmAlUHMQ7
rGUBx+EYQv7jmRsAjpeSxkjhbqWeXWjVp58xQYfPFAsrHnuUvJBpRiXx3pvuRK76DBQfvOAVEtK2
BjaAq3VNT4bx01Dt5cV4+L8x6FDKljLhjmfN45sgsqLEPlSPIqvixlurLy0OCAYgEpo9+FWhIW6S
cuewfPSMF9WQVY5F0Lu92IN6jmPZE/Ql4tQwZiexR+XC/S/3Bir0JRdfb36gQhmjGspXaYxTcxPT
gBtTqzQxbXBhXw0yFPOXQrL2UH3HoyJvIZgx+ceHSFn9QxiMbFnMbSvYLAXn/+6UsDQEI1ALreTV
NGkIqoliFygHuwz3Wtu6IY4eA7w+suB9D5DDg5Raaf60+NeO89YIUKvWnf//8C2IigtIHNj3bM9R
Ena7BC3rETGTy3n1BTpKF5OsXVzVe+TTGgKaswQndJeeuM7YlxLWxQnuCbNfdVcTcYYcqcBJlZal
4FzB5H86NZEMUyPHxM2yDEIYhtoRCFAnTmy870U/RDBv68DlHbHPnMxW+24Di6dcCUKaSgcGOrrt
zt+g9/ksQSLaGTSfwk5jY903BcmSOyVC6VvFafay03SPwS8vioSu2ILZZTiZnS0OF5+3I/upXxxT
x1rxacEMRyjJsPDSC85CzcPmeuf/n52KoOLjT4HtVd6hFv/DO5dRZoZguF6T8gM3KkBfLfiXgwHV
j+5kEB/SV0pwJCm+ZcNVQiiqhqUR8MvZotZVrJNm06tEKkPuQVcDwJobKzUate1/FOHGpa6E+8VB
5IsZ9/apy1klb6GWBiXpAZstqtdS0jTGlpKPxm8u3hwLM9D4IbNET2ptG3GoLy2x+K/wp4eFeM4l
wgvU8HNXBnmn3jU5MfKjILSlivyxj4GPRkHUiDr5l8J9Pf+5LXGudaIwKR7QrQ190ymAUuLMLkd1
h36Zgd244JUBSJ5+xmaCbbjoYitr5Dx1LZsHERvVcP6NxKc+b0MakbvfDWj1xZzzUbLgEVRxt5xH
ebOooYLUK+sjsJCY28WxBsAKdnzfQanF8ODqnUeY2jQfj+u50NT9c7HOqqktE9JfZZ9SbUQsZwON
2HkyWyk8Ppecf8VLmEdI9SwKfAzX2/eb71pMVg4pzADVkxP5AuvoRXElH71sYUhQbt79O22GLFYS
t5C86XVtyvnEQfWBRWveu0nSSNJ76gBzIm5hQrWq2SRVTsu7IFkUbEoLaSQe6Wt2PHiTSOlrAxem
DapmG9rT64GzDcQBhcGdZG8HIfGwJRBMh+G+LVyOIO3ZS6i1FC2n0SKeX76moA8B8xA0oEdIT4zl
ZGXJxP4sDDwWjMb7+zYX+7HsMRK3P2nLPuAkGuqc0l19wwQKAg+TwkWEl96xEFOOvlapWppvh1ZF
EnJ00UQvTdF3GeUIvU3McRAgcUptpU9VS9/nsg9KdNN1Hp86gMCx5rhzpMZTasU29FhrWWh72003
xSdVQnkJXN+A7+U0q2sFaQJU70JnRbdAgzr69SDMIR9Ngpl1mdlHuGov7Zi/Sz7DURqBtDEAOOJP
T3CgRYK/GbtpMFllO6TA3b+fqHti6U9BTrpc29aOQ7+Dsx6WXdXUQTpNPxZ+KmuKAUfw7kP0Z60F
+c8udawCDxZvXsUM86pfeZ+OROLRfaC5m3Yw6MtzSiKb9PI7dZFX04+vQEOxbs16cprxgpnHv2oG
rL9kugziNca7B3LENKjFYevgjLMMi8e1T33/qtUEZDLd779C5Ia7nWXcPU4T3M0K0LjUNnGtVYHH
uKTmYAR9F7ZzkD++8d/0hYsdU79HcC7D/wLP/zNbPhZrh88sbMt+InuVMm1iTW1CsHP6jMyxXq+v
g49wdA+DYGToRXvQ4YuxjicuWQNMiUzm1iGht7e2kMeaoPdjfuNmWrbCLdSBnRhqe7QBNrDIgP2t
eAd5ufh+fXlIMy6AqLUhkMAVxN8NI4r/cq0D1MaqxlPXRXe8V+sec++vcwoJ5NIr4kF4iTNW7Zzg
ieak+m6bpWyfivgEul+I/xpU3DlAiMK/NGv5H9kjoJvPdYgAaUO7z6E9uF8OtfY6BTpTqLV/5dcv
CIbDPV6d4hkOnfNcKe1XOQnvQHTJc4pbpwvHpEmp941iw+BLTHsh/9g7BkaBGqRGpoEMci3iPpQm
Q9lQWfbEf5Dop3nol6pUL9YwW0Ocq9IoFcISmApHgoV2kaoxEvFJ9vZVE8X8A6zzcNAn+PSTn6bs
KLcX7Hq6Cl31tB9pppinTBpLD5bsjRr+Hxf+B2gfKBIwjuyybxkumUUp0mxUvMYzqgHcCRAGVgoK
junPESyawfhu9iKPn1D64mgWJnLypISKeh55QN+sdKC0PzdXfAAv+SHmBTQIbsBEUS6Uldlhs2sg
YckO9q5yIi16uJRwfGyjJZ45jge/Jx9pn0t2aJ2zFPZ1zQITPMZ/vD+5Rlw4yigV416AoYclQVWV
Q9q2EgxzPwvK+Capdcc0iGUAlrnLhXNToS/4gH3F8db0bid/NwpgBYWnOfp10h+adNZd35uxoSzh
T7jLbWSIQsUy9g3K8u/VMYXNHdaxTE5kM+sxShFydk76ooPeIgDflSEIFsyy+GjW4lTxghFyhIHi
sWmIgtdsAodRaHp32TBuX3Fx0VhN3CRJo2eAgGeKoEcD6Uh1/2bt3OaiRNDx73W03yYgVlsx1HaO
wY5xDiLMX6/XHL85mAafnvij0sf7UFeyrUbWjWk0x8IxxuPxy/7XyY7RMpz0o3QwrH6exfS1K6jp
Qnmh51OqneJuM6TDlm6fLIy7vw4mRPu7Hc3Otj9EZx41hi7cDvAaFtKz5yYsT00fYvWdB9xsa8d3
s6fDI/WhXN4DakDUHvAyWMQTP9uazbMqBzEyi4J/B00r303OD6UoH67II2JQKgO8P8xc7o307ux0
G0tgVKp2llOzO1hieBaJMhlqYyNfmlElP8TbVSh1/8BSI/ePIJQm4u4AJaRUz2aC7rCqLZTzHcee
ImLPioIi9laJbgnExF1irwAQtPSOpVp6OhYN6HTg1PKzWdHCdeEzER3WGS9Vs2BdKgfzPd7lebFx
xNFyJ10f6ajzCmr6xtvhyCJ94aNZh7oaJMhFF20layT/v76Qw0yCHCnIxAr1hBt/rjkiVeHe+kli
TjwtDizD2RFoz+d5lR6JbzF7mauo/VpZVtWampjcaOQiXU/ZYdHp6BLZmoKHdudNqNeIdOcP5Gjr
OEUONcejx5AnxKdUJceZf284fsSjjaaamHMyOPvkZ1PPWDf13LIUUlyl6tLKnFfNRLVTiPeo+orV
11Cs5RYp/0NXelK49u0dooFqaITGdlsno7yt84tOtZ/ocikEo9n3aEX3aZoKOba55SISRhchBl7U
MK3NvjzKUd8y4fPu3aH+y6CBQEm/4YTrJ8jtM4nesylpADCJLIocxMKJf1FKFwv0lRnT9x8fen89
oRRlLc+ybY2e5QWH16kc9FpR91Y0+0qA0fNPyAqbVkGh0o0N2kci3aBhcsRFnyM8HDpoSSJOAsgz
1YXMQuWijzTffj545cdI5p8zaYQy9g8FNhC4AbchzROih+YiPDMzBtkYCBHbcZlVo30rbphbx704
IbGQbWPnHGZS0CSleatbrN9f6fXuV1vtkMztCjmcmsyV8XH1aFChNe17qSCtRWfpPY/lBovK3Y07
BB67kI/uHZzyt2B/aqXfFcZxIFtvqkul8D4suG4Dnaa3ElFEJnJ3oK0oo5meQKTyZ3K0jd/paAFG
WqoJlsF1lk3vm9obH2xu4+wmETmvIA7tKgpGfnCax2FZdEkj8C/OMAqCx9LuvuSZbZiI5+PJ7S4h
Odd78h7UxNMPkDH20e3DEF6q8jIF0H15bUjrnZFqPmj+zrOyMOmFsH+t7uK6Oj7slsqqx3YKcIiV
9HBxvCC8dyeNM8umSHFCBhgDoaAlJIb4QAZ/YXr2rP5F3ub/D+VVYe09v5dG/mte2KwuyKQJvS/j
IH3zUsZcQNEvp0EkMZjBlpXDLJKtng3iD1+TXGkEx5gQSmrjb1U2PCnGPGesAPglN05C2F6SJqgf
LD+c6SpPHk3821HoZNwWta35vVfoC7hqrAX9qrgi4uv7tqDbFsK2uI08LbXW5Ymx0ANwbIpBKHJh
lYG9vLPtCVQBYaMSE6UiY6LwTWzVnMEBTvoY5/yI+n0/V4NBKQoCXZkWY+rXMomk9wAspPubYV7x
2ig6wOaoOpK3d7wIhnO0Cv39hioeviGNiMJA0sKOhouX3sRODDrsIkklU+yGvJGrWKM25JswxzW4
rRfqVrvLb3ctJlEHxoT6MfO10Wi5Zv5BP7WL0k0w12UK3GPeHLj7YAMY0RrCcsjtHt8Ym1UxhqRW
SuGn96elWuKVrgqq5PdX5QstpdYd45JPXjtTBxQzT0F5P8p20I1Ybbtl6z+A2aQdnrIxmxMnP1B/
9RrIPYyrvhTyxGXhT0A22j2ZhbzvQy0wWcecUlNxFfQnhuDHgirV0J76JeBQAP7Oxv1/SlwtgAig
KvnAEVSl7IG5J1BR/ojtQ2ZtaAY5uinP5n3KcIMCTPqtFHjIFC9b3mKCVUz+Am0c4vGCESO6/2/x
5NXjtuHnc/TK9gvG0Dg//X73ZR5DQ4GsioC1MOZzuWgENvzubPrSnRy4PrEhMhQ1F5QBsUG8P5Hs
Anm8ovE4mYR512eUyT57DsftW+rhsx54AoX3ZFwYmxC/0A7EYerrgAfEHF82Juy72QyinAkUeams
/TmW5cyfYbPz8AfFiSV3v8IWujQvJePNpzujZD3ZmGLGBT1xbC/UuqiTde8+az2GN5q2aCtNW/WD
lyk+VuSy6gNlI39GmYZ4DWJHlEebuaTt63zTGs8fzxxndCv7PJNyJXVP+mgmpBPBDYs57ptp9Jbw
SICb/tobzQIJVimTW9i5rZ50/jmIOqiYR1aWzH6HVYJiDjXFfZdK0o+GdZy2LwgaY/qr5TWGqp0B
UHQnp0CNEIz/3jMBJ2flB98Ius7PKCHmptjcmHt9dGeLriD4lpnoUkFNwfv8+O1C5uAC3zq6Y7Df
YT5VlsFfMi0ESS2bNGf/C5nEQfw2qA4QEpCydYGENHfvITlZnf4FskmUtVWZYymrBOWg+ReyUFLW
phvdagFamsdxJq9DXNn67PCbjmi3jOvnFthwZ9DPKoUgoY1OvtNCG7jnGVT/9laHGkunWkeOdmAT
4z1wXYVJM2gM8Dka1uYBSE1+NxKkeehBPgbucs5LdTgxG+irOKOyFs2FDht0uxitfCfMj8fFWA9N
5CBLfQaNJuZ84zT65/xNiXfgeUNtxdkOpePpreQ0ko3V5DtSRqd8ZTs6lTpjxaAmD090OGf4w3qt
3HjS0QFgtODKaNeoHqjQz/MOw0zYZ7iC2+E4rg8THWgYJqVuxkN6yEPL/OlvMZRQZeT7sTKXpswB
mGoLpNgt4AZPF7gOJX5yVchDSAbA4lAKhHRNY9SCCDsu32NAKsU/2dlVJBJ6WsaMR/KyNFMvcNbP
Z1OqX2UvaD6Q5NBWdRiZvj5T6PMki7hYzi6v8IuGhpJgc1rEEyVqdXNz0fYx3x++fZ9lzZJnkJD+
X+EZirHuu3Bok2C2aBZVQ+Nhb80WdimEql5J6Pjb98tE3lFlMqrTIIQQdMTCRS+NVAQRtJyazFuC
VRzHGIyS7MP5VBa2io3GJLjsD2Dmr0StZNwARedqy/TCEGTgl6jRsVp8PiP5NfDNdJdZca0szngf
+uYwJC6OoyFM3bRV9A6OUSW6EpFJnLczyQBMkFGhrmenNEr6h2C59SrJ6MHH+DE15v2xueJIi25Q
dGPMFukJy2pUJ26ChtoOrojdSjlSMXYZ6DsnuTh0u1geueYPYf2Ojpl1eEpA5ETQZ+DLq3wXqhRG
oheRGPDKkrFlHW9GNWWqt/p83ebRnBW0aqnppsJlHhO1KxQ5L383uGXtOGBglb7uPopd1Nugh3oH
HPQzb/CFo6RX1XWIfKz7qctPpvDzSvRsTlg/0dveHSgibx2+j4S3BJ1htEZKab+DjDrpviCsbaLK
KXgfYkfK4S9PjUnla0FCN9xqluH87Xn4OwQ76y2QFUUhK6q9mUK0qdEaFcKjY9eD2nRzhCBLpRBU
2abMLXCgFZF2/83EAvjbx5mGdlK/zBg76b7BTLSDNvbzQ8u8B3PFK5n+VJEbPGcmS3cOE6WCf/oP
3RCQH9JmTQF//g7GqOlBmvY1953012GJ3sJI0aaNYW/kIcdYdSTis/Q6T9ki3//CZPDAcaHdzVj3
7xOpEd2C6M2GomW+PMs54nivTjZZ4RGwHcJoT0Z0XBu8P1wbPCH+wUiKQ2v+QDeqn4JUfrxbIss2
cEEagFjYjwpRORYENaS/jlWdkSgjYodWuuanfG9jf89euLm0UAkhbmA7WU5SIA7ncYu7scRoLdne
+ZC1wdDKPz1EXK2KFqkf+EpBpy8qudpHe1TgmaYODiHLGPquGRS+9OGbDIQiMZhyPmbavjKGgQ1w
siEf+CHKWlbdnR3gTDqidYjx/4u7zXP7wmOt1W4lfVI5HZB6GsF3vfDsHBV7by3VLd+mIGVmwBB6
ZSWlm7iUwQBzHOPvaX+Ux2Q45xUcpeMagBkEyVY21nK1XprMOTWvi4xbB8Z/lMzScDRWbA/4sKbQ
VDlUsqRPaVoCNjVfMUMNLtX4YP00BV99RqyzT2kd1NN7H/lzAbrpax1KVbA1+JIng5EfqrJSPz1c
k3aQHHEi+amCd/K/l9Rv4xAnBCt3QfXYuASBcuCpu2DzUaDApyB2j14KOiNMVXPXtbvXKtwgBiTg
b5cOPRxgz3yPhIvzbUYmhbmpZBF+dxR7E3E2MIRxcg99cq3q2uI0h13MylfIRwHee2aKzsUnmSiI
f9CdUAQFFzi+nyU6BR2HKHX+zJJjUvOpAlaPv5FmY+gcr5iqRBNPAXNMqA8vR0tF4RUAzEx/BYum
/JR5ffAJAULWOa6sCX6WKb0LTqlANZ0JuC8TMKIAP7180WyUf2mRJOoK5fUOlqSxpe9OP5tTDSJ7
Mv9r1iR7oGvGIsvtgQCG7Xuj+2j7dZ5wGihf8ok/VmLpYkwPOZneT1T2Qn577n5UA6qSbIgGIX7p
cLTgrAtp7bYMokY4wuEFGx+IhcocXxLxuax5CGeCyrLO+pvMVBBvbarIm+VjMy6fYLbWT3Spu1wp
nyPDU6IvgtkNRtpZm6lIKGCeajnJpAKQakmT67PQ6lbInECm4At05SBFiPlhNo6kRMUS82kYWT1R
RN4lBYb2Ef8x/ABxs8O/1aDHnRmtpjm4R9/bGH2yjVXsSYnuJsvSUmx1fL+WRSMsJZbpgMQr8PTr
40J4/C5VvkswhZ4GzU/5QQ1lBV+HAWMSC1MPu1w8u2vb7g3KpeOQkN5j01Vez/zTxb3nK2ekdosV
9MEi6Tmt1seiWHOI+dOPUFVJNK3ja5oMheL+dtKLFEZnQutOQiQFUisUT9jGXrSIebhh72KNpfMH
0V9jFYuFqgUtuhN9qukXSTT7zGmnzSgPDlYhkwQ6wVyP+EJG6DbjaE5d1JGfCCxKpRHDCYzIFKiC
vaB+h0kmqjPXsPBr88MetbqQchcJqOYXgMok4FWu5jHX95oXzvexBey3lm+7hckN6CmPtAGhHDUv
tX1NWgYRESRx6Mw8ZkvIHK876WcO1aDMiX4N16q/DF7W0xHZXp5x4ODFVOe8snSCJiyad4moENfn
2sJ5bs57GQWrO22RwjmYBf4/pkdAnu5COL0dJhZhHrQIeIuDukAPW4pHR7V5NmdUYqXwlHdGef0P
nLGn4LHHlEWYJPMIdgJJ3Ni4fXncbRj0bp1YhPBSOloZ/kAPB/NGEfkHAujzY7VrjBm388QaRz6F
atqFtXOEVFiuo/iueBDWMwjvkpD1GrupS49X5OJg5y7gi4qgqV9IAdS+kWUM0JyrsK1Ho+2hcu6g
tB0uAk/Kk26fD7GE8VktflDSGwy/Rm3oe20N2mqolYzk1ymyqllUH3yabBQ3Jcy10kiFYlp00IYE
ggQwRcOkgqNnmdLtBIaglCinDus2jokbP/AoA+iS+2hX/HOdrYGz5Se6ZCrRfZkKxPc8ZZ7ZVv/M
80SmnMwUGFl0Fzo9CwMrb5tTyzVgFzvYj4vKLwknRXtzyav2LpH8b3Ckt4Go7B47y89RZQcgh8hX
I1IsdHoqvg7uQHr2EJ8mhLzy/ypjgyB/mlgT+JlNO/gNsQ1WHeNLlyMMLpBwvATzSfasVxCO72Dh
5l2uUKRrII3qFANDGmb0tRoPfV/tPpE4PwgVJ5RPBstL4FUVOLVg8h+G7+oaBSejr361XCDOpkVF
3dq660QMwkQ6jhnpjRspz7VKh7hCmSOhlbPP5cMKgcnY2dKZOWBPU9MHzCY0MH7xIvo59hE7PNRD
4E5KbNRgfpnBTb/nug19SU2m4OCAS22eMbjXfAl4T5YaDhd4LcarRXQmv93H6rUaIMtQNS9RTkHa
M8UhpgzoQH5mj/TWoB2R7T8B657ZUiA+i2K6e0NEILQVMY0rTOgFQmWd8g/DamcAEziT+1nhUkIe
rQXgDxUmvysIvdabML7fPFiLIasioOWSInfN2g25YD9mke3SkOLF0kPnZscKGk4zq7v6OdK+FR0p
PbGywKrLHWH09ISZBT0W4GvyVDH81L6oIM6g4ooFgBziRv6ToFl4XnPB4lVBgaFKd8thTty6iEzu
/46UL6ObYludB6TZ4TgyZ/qzoLkpzpHVYIlkUl+7Po/cfi653Aejusxt+8EzjpHeW4W2hx+VLaXv
rjlFJ2jlj9sCq20Rj/gb2ixKfAY7Dsi+amvuIOufaFgSKGHxGZwg8x43HuaVWdby98s3Cd+5H6B5
RxGwUYTOkir0WxFD533zUS/pA8Y7cxh0n9/o3GxR+kZjXnf3bShv1aEnyxYvvoaVKfwL/q43VP56
PCwFk1boFLmzfkUQnoqQEGvOClcrLWHkh6EAW3McAVYL+Kx3VmoNEt0FvnaoOP5SfGwV8CS/Rsy1
NpsvlIWv9kqIFJxSeWE3iQPQvnzZ/3tqnUrw/qEg2E6ONAfiSkgd8p8AmO5h69PbN4BISUHKe48e
Cc5AtYc6Beb9Gak0O+hfm9VI1FFtG7X9vDSMoRfEeUWoDtNNQcOWZZpyE5saNKs5gFpgn3ELXKxI
UoBhaDU9XbrjD1Z7xaw3POm42cO/Dj/jNTeOy5e1tjeAhewyUTQj/eQ43TAewoRLAyE4dXFQokTg
UlAE7YbOCe4pz2BEF1Lp6SUHyvkuVqJs0BSAWnVQAI0bGONbigpDYddpalPq2pLPz33rZPZ72Als
xj9I+9P0PDEPdz2DKMBeuj7rkeIHCD3y9FZcbaziv74ee3O89mwqN58vx4//effVWV3MfZChqP70
RLGT+BISdH1IJBJeHv0vinsYtTxsN44w647zW/GjsO+vc4Y/YkRhrdc5Q9YDl3EM0+lzrhBxauCw
OtR8rcxokHgE8IUu0Hn/Hz5X32TF0EzTmQfayRlKmvV38OIHhbTOXb2tpfewCQ63FNaKatjsLgxY
+lswBZd3M75AcKbpAym+99krDMhIFvsl0JixtBtrU+bjxt8/baK8A/OSWOpLvoFf5gRRFa4NdyvR
e6P268XqZFYO8AS8IJp/J5owQ+c5ZePXSyt+9VvYJ8W4PPa+Ydy80vrdtKfFjPvDzX5r/Yq4Bh/3
VrfEQjPKPRFF3P4/AwI1Hkq/KSgagkZdoGE2mzZ//biB6SRZ7XdkTL4q3hPfqbcNQ8S40/Dqk95Z
rGc4mjhazGqVzFgwa1c2+XTEB0vmYO2mmi+A5C0AhLpEol1b+ePyg1SANiARx38I+Sy3n/pj6aJt
9um3agHRnA4emFYwyfJsLxdvsRQNnirNCPJX0PVNLzGJHTJMiz5rtBoU10swbq4FxVK9aCic5f/B
yv8UNUN1GZCMGYml/KgzYErU5fd2ijZJkj+cgIJf2aOvdCHnh/AiypYw+BqJDJMz92q813UtJiCk
o2EIpewHkOUelfmdMuFQI650Vj2/Hba4KYURyZQJnfI32P9/6/mo/pXP1o/wdQ/rSgygJUzItn/F
MyVSv4BSbFvLkocMhAOETJDeRTjUSaDSNJWX5xJFRfMOhzEnCUUWcjmbThQ6w7bTN/oHp14qcm5v
y/o1CUqkyg9DoqWt6GswtrVZ8xApAn9/ep2oG4fUlT3fMji/N6cP4bWKUZ6CQCLV4VZRPXHsl9GM
oAtqeidtM2uFIraK5AhrJPFBXsscYRM4/d50Qxxd4ZDZ789TNIrC069p0/UI6bG7VJzRGyCEBsJx
KsY4DbWfxxCYdrZqIqeD/SEyy7gax/gUkatWrPiIrH3D+3HGD0vCPWKqGt/LEZSjYJKjNHMYrg82
Wkax6n42qeNbXUgqvof5ITJq8bkegovNvxUaZ9VqlVN6bO8Tq3vXDh6OF7cwSNWi9bsuB0rkGVDx
0DSmHk7j2Ub/8S/49UtLQMDOFtS+r3Ix/OkghiEcE4f7L1WgOSktijpUP5BuQ+H/fWtgn1dYr3RI
IF3CFN7cp+EkWnDQ3vWXixDyq5eXnLRFrxI1Zc0jGPGMeVml25iNvMKye0c6gH+b5+rPuWKNbFAQ
S1dtMxcpFD3ZIj+StNZwm3MJeCDJk4CoOHnAVlGWDuidaMgOYVGdRKaHVeQOxrh8DIKYAeGpydhO
k0v+Z4jmZJkBw32x1F6FXe6sSz0haPKWwOoUOG7G7xHhTRJwI/pnftIROkJ+dlTqPxdA6ADq6GMw
Y9qJLbjSOPebHb6HlEZ/i9CwzObQbIOfAPdBxAmk1wahmtC5xb2oA+MSP4vOt+nj2FVvedD3Wa4b
6+FrJouoQi5hWlWHJZ8Eo84qm9FkmBRAMWQQN8bdirWP0gaGozmCYJMklAJm6nCHishsGb3psGFs
jgfFMG/CiKgbpGQ4fhXwamC3A/zd0yxju0vne/hzEGgpIdZCK2RuAoof27sSSMGDIRVAsGZrPcHf
KStjCAAYk9F4J+zzgtD/RWOs1ol2KtUNH0MfEmL5eUFsZ9AERaICPnX4q0n7UNbpDmD77p8gQhLr
+HvZCjxzHH471PXiiX4yC3YUV2TkfGeEttN+A+Vx+bygneOdy0E3yKXZVjIScUUJlFiDqJpI7Sqn
0WfAY9TLTeDj0lAHcEU20bIoD6y0E0Yz6E+61lEXtqXrDv8X4BLlnQ7yp/z3DKX7pa1lF+x6qhSZ
ipGf00AWJ9YTkVGnQmxQCfdxJtaA2jeXaO6XuyoEqC0jiGXxgGlv8OqluhbyoA9pWvM7qkbPMqT5
Nj7DXRcAAvC+9qEjGkXy5c/5K26a3uZLryd/xlgBKyiO3tf+YCh7Xm5Jy1GSNI2lvfflshMQ+Zfz
9h+4JJcTEsGHrfLRNDYCpZQ6EPU89iTj+gfE5cS6+dO7wF6pFEPgzwWl5RQnf+y91CT0t3BdhPK8
rZSCGZZZ44nc11h6drTsdHFGAx3ehoRWQdY/YCWT32eucWZqmSM2GvXMFmKY7q4gCPUOdVcebOe8
qNJWKWaOyPSB8RbkMzCf+UR+bh9UN8LvYJIW4/g4pMTsQXif3TBHSlWTr6AmhfXXs7BYsiuKoDcM
WIj/HzaLCyxsIRAFHgeguL5uJG/K1Th7GHoFnPXOo4DQ4bf+ONC0VE8R+ASfc/lDJju8M+5tbvfi
k4IycjOsXnf8olWGr5cJD/65v+gI3mooR6J68JNSRiEjS6CHs1zHd6I/ZuJzuzdCV/A3EkI5q/oF
d7Vv3EcEfWMqofx98jJmNtIPqqI11/UAJf43AAZ56NiqBQRkcV79hrlDL7lfKq1MhC3TwKSjU7U/
yXE9mVhfjxTSmcHLcZwKEVSE9x0VHMH1B/AMneFpRk3rJUub5EgBpF8e8I8iSoXiG6xl7gwTRgP6
oI4ZJpAKh9l3tGZBJjsEPGvmdV+awso5vmSW8horm9L5YC+U3R4wW1IoPc+Lm5Zl0OcXaV96jCXV
Ysv8c21G4o0kImxuN9ahSH6IshMvQVFx5+NGbeFmMHUAUfTEzV8/fggzRcDAiPROTbvvm4ZhVOmr
rYbkd+zlNCxW6clBcXC64I9jQJnlbyNyw9nlE5mm5Gsxq3ZtL2MrRgCtHrhfWNvpBZKJLKhlwbGY
rF9cOPZFhFXoJBT711YuylMxqHZf9iLFqjqEk//qnxahzq0HY7zbgcBLloMh5FwvO/X+N3n8oO0t
0YhDyGfa8/wuDciqHsHzxN56gikBhlQKEiIgAd+7Lp/yfzJktIsPSROoO9cbBVfnAKsftm7Dw7+i
H3z0NiVn2YB59bplsbSyiymGwOG3iw+Qf9v76ftfjvE90VGgCBHJGrnZRS45q5EF15EZnW2T/iUh
LN5/9Nwq8wi9m19loM/UxHCx8h5/Uivkt+sFg7naDIGXjLkeVoeFs4oobB31ohbx9QSI1dMKcNGW
27+cE2Z5FKoSmtJxZXCflIZib6pNL4Ip2+u1ib6RWBvLzrg2xI3qCXnEGVmRFNgV3hy0wbT5ntvJ
I4HCFeIBf/mB9wdL4bIi928U4mz1eXDGkJgn0j7/NQmqVr2B/C8ezywyIJtlAACimq7roHk0B5BI
KKgMAuM1db68LlAQbs4Z3b8ieUi2ZTux+shDcXeYDAtjh7IzPPJ18ZF+bEN6yq6H6LMojpRG7omj
nNBnoqtlNviiSqP5juh8/NP/6bEKQlJcWT7+xWh1OFwu+mnCs/Nl6+36L5NYAmc1DDHU5y9ixkCS
gSUD7cNQOO33JUFVzwURfbnQ9tcqau6Bus7Am3VFYx41B0obyQnJEMhvAUCoC2b6HvusBw3+Grle
q1g3vtXxDhAZJlEThelFuklHSp13sAE4ZuONPwZBXSRb1hTn881pXZEABibnRf6ckA5/79XQYW//
LcfHDBlY4V5k8HvQNXDjfyfoIj9HQZWmTHnafBv3LsUi6ipLHzsd5OTKRUMsRS5AjBffVZ5NvLam
UVlYx5SHFdLt3IpC3kws5vKIIcY5dXBME2O/eot6yJtqw/OaGZTL9EQ4TS4KphvFfkKW5yTZF9sv
0Uk6yNGpjZ2nolbjk/w1LWF7XYoLb6tGJA61KJGXPGz4X/JRtZaSmYYXHTsNH7qY+oC3kI0J1v3d
eUqsUH7U0yqbu0/6N9/1IOUysndMo55rseEQxmDwqhxFWlkIsNX7Zx+pgChUV2fiJon7CIhxvsHq
XX+RVwI1HTMDmXSDKwDDFJuVuCUSqqNcCQ6+SQQVVA77OE9e3WtMbmHim1dql4OJMBq9H2rNolA2
7wsI8i1YYH6DAhqJvv/g4Xo1dVCLWNP1eQcvshc++97qLZQwVYGYwis1CRI1n60btjTKK1uljsLN
80XP80OUlvGvepgz4/qCKeND8uQycou7Qi3tj7ovpn8GlN+xFspxfMnVCqfQGcO+7ygB+8ohjP9R
wcFAtTcw3FdmmPA8BdjXkP1Abf/OrfXjol3dbiAJDYNxe/ukEceHoBTQGQiPMbsPsovDK4c4EaAN
v80AphiUo29xUdy91oGcQCYEqfwtWK8YNRLzVujIhNPAYk2DptKoaUgp/fi6M1fYenOGaOLZBq4r
ODXon6QNH9oPaMRUSog2yJ/89nCWqA5kCxibISGN1mcENhQVBrenvurLLs0DwfB1g3oK8/TtdmXn
Ob3DCv0FV7RBvYYTRSsGYWA3Yw3Fcg0TiNRK0j5hZUyHZ5c9vv+ojw03yPWgOy7ZXBSSSBNR6MOQ
yUeAEtqlttU4jt+85jgV/BWK0+La+P7I0rI1HqGOTxJ3e6YybKeiBXPCuzSrdvzwaX7Ql9xn2m92
jV4/4pBZvn55nFOJI3JpN7Gv2EqWE3UECiJXn5cZy0uRPN8szkNZfmkTdOAzpIIven5i/P7ImBGQ
Dy/5lF8iTCCzyYokNB//+wHJM/G5gdBW3A7ysWUfXgwh0Yi1iUw5PmRxuVGxNEwQhq43ArR9yhjX
G6kcR/81GC4b6foootCzcVQBz79pPJxmOTKkEt+Bvts439AK9ORBnykm1rTXqKQhti5YCX4r5U4X
dAQfdlZHTMYPgw//hOmUwhhS7RhL4JQgcqyz0cWYH0BbtfLCAp7+Y5bmL2RihW5acrjiGNvPjteY
SRHKhrC/XFyUBl+7SBipUm9u/xWOenRFIVFC7YE5ajIfAiRbO+O1txsTE1iYmEmdN3x4jM4WOePo
yxRQe5jejHK37L3Sb/Eva2nlDvGVkKsDCD8PsNVDF1kSKwBOoYlKokEjdC6kd8n9cpCgVWDf0Iqv
gBpHUgnnMLpoXHGK7DjoJAAjadx77RONfDULKqcW8Jbb9vr7RXniYdD4RjN2Z1Od8OgdgBn7oiJb
Fo1uPaDCHauT5vg3gxMM+RmKr5q71L4vrSmnPEVCzDl6LM/i2U+pMK6bBdqc4ArWjiOv6P9VOQi6
zDhBYuZx5CZgMHTdLkgxzh9907FLz7ln+BuOLby5R9X9j1jd65JVoK3nfJezslTDOiSwonuY3Pqd
U2WBoRkrX18vvl/3bnQ7Hiv5CWitC+gXHsKg+Lo4KGRloA/W1tv1j6euwPtKmyRFtLxhVH3JYaTW
Pg6uGjwzJU71iFLPIwwcfKrtr3hBIiQ/P4Hmu0eInhUT6sNNreILN+b5Aim5mauggFOf3I2Ioef/
1PfhGd6yB1K56WkYEPAsiMibeudMucDvVtVMUgal6WDpE7wlknpuazwsUnHyq/dc4WTYXTfs1iaQ
MD0WVU8vNBr/8Ci+b0aTz9ypRP7uXgC+ZA+Fw2Lh+sjhj6OzUl45Dnzw8AnJyKweP1IwiL9lWukj
LN2LFDT/SIifJM4uOiV+6kziav22aUhkrKk/P3hebPWXHiSb8oAB9fn3KFjHHCbNHL2s/Tq/4DbB
d7N+JECwV2HweiHt4e0gv1UlgZOxTWQh8W9Wcc5LC0TlngbfhEFA4PVS//RKGJNlKjaDotfLV/1S
YljuszJyhurLuBoVZS1VUHspej/D4f9L4o3ZOS6HDY6LqkDy4er7axjct7gOvAojc7pfdRzjNCiI
Y6oyHX79xM+IATVcNyPYTU4ySh2y6zqo5NP/u0KfmpuWj9TynyE9B9wRKjbnsk1lkrmSqdX4LNPu
xqxohrcz5HuLjiB643sgn9Cz9kMILa9tH7BgsX8RYvJZ+ePjem3DpAPtzVXF8xNky3KEe/hHmo57
GPJsCvkXjp8Ij5iCbT1wcAYlGIY2yCkvDGgg0yZswkMEfzVr4PXJ4lmXRUU0vT9XETkO10PvCXEP
i9c4D86lflveaIsqYNAOyp92HgxTabJywQFg0KB5GR7tYcC8E/husXKPylp5ChUMPkOUIJ6i4uQ+
wUn1cl4RosOpAw1Wbl5MsrAfHcbowKEAicgVdLbHNbcmb0/gTyGRWeRmHtqzFzaFESFMOV1WU8h4
7u7VvfkqKXEsoztJ86ICe0QbEE7YQSOdGLIbU/ibQmusuJRdYUZ+MQ4822nV/Q8KBXk+3vejPDh4
gOuzxajjDAeoEls9+NbVg44pettLtXGG0IZtddI6bKy+6yxlw/r4L12bql1tcOT9uyFO3cXTTSmw
devMo80z8YNO6WLdFj/H7GOaqQf0aK57hrhsF35hVnyurOcEFPd9t0Z74nyHQciA2mZlN7C8JEUq
Sxy27vfCJl2lzh0GDw1VkCzyiMu43YF0CBbgVLfRaVHxM+bSSuSR8v/STVJvnYqKHpsLGCPHFxMf
sirutknbwQVqusVEVGS0H3s/DQFkgbj57wfQ97cMzaikGUpiAl/bEr1pW/ilB1qbiGvRbtDF05ad
UQyu35YYj8iEVcI2lUssfpiCSbAYSL92M5CAHNcjuO9F+fwsIUOXichkXquMcTGXwfhT9eJU7hY2
a6j7TkYhdP8YjB6A0QyKwxcRYkwHAaXx4+/Y4zVRNbzKNctbZI62OhRUA7jQGJhAJ8UYrQu4ua7B
JesIGdWCVU/hf8BXF0rlOdgdBewcyKS1BUXeR2qoAqctRRn6aHA+hjy8wov+2MTRzyPlLv/pFlQ2
fbICGEG4JKLrXH+dKrT3nwIazVRom3CA4BdrZNk17zY+O1hxMRmtT8z1hn+3O9elz1SrKmFsmxNU
WtvTcwsjcsUqtgB7dnypmVSt8LUWnf1EUuG2hjbliLO7AZ2g4VJUMVd3wmMraUURhLiWtX+0rs6X
4tZtLo2abCgytvlVHnLq+zDinIbH7VPEfxiuLbnoSywNSJWXU5KFVO+6vxE15+pWHGdYonEkOdiO
LHsJg1w99RsNClZq3uZml4fKsFam2AES2EpP3XILNcb6Pv8mU0MEOlgGSMXbMDED4MafycFj5chF
XfbHcRa7u+Kh1sSd+qI/O84rC5tONuHYtdKlcyz0QzOpDRpyAbucg/P8efgch+EIcw/DI8AliaaC
lEsrjpG57ToR1gFpmpKlNXHjR/chSgT9ysk/N6x99s0jYVoH3CscpZNDSLu5bii/6iz7f10YX3+B
KAAZyKwrwgGacFU6flch5ICrv9QA5MPyO6c/KZJksKh7XNppG7ekwDL39mfVmWDE9I/nm+IJRMv4
UODkpH4m4ecBclZoJRaDt4lDtZVPTHkwiNeZXn+cXL5e/enGGlunDPJ0yfhLQCqXrXKGzl4dVre9
0gS5P6+eNlRGXzJFztROpTrfc6I6QzylFyZZQU60ShOCuE+piMUqjX2hiBYg2b6bZZLU2JopqgXj
F5TgUeNAazTI97fGnfCckyD8gwn4w/o2cBXFPFAnHXiLvKDEVJD5vnVHcz8soT3NeE9+ZeizCwd7
VwHlKp6asMxEZyrfFLSlGfy27wuMA5WdR/WnGfl5+6LrNJTHaZ6FdEEFZxJUsc9VzrJf/17JFew4
Eq2ubfUTWPDS3GJQi3f0TpiLOZ0DVG+14Xam+Ygl0481s6pzu2gDHXAWxX/KZxClwcCLcNCLpDdm
MDnBiFDDQxyqgGOTaKuEhqLFWIKXDtQiVYWgvir6xgfI+cwdsZ0m/01Wf5Utuxrrw6SiDGCy7VgF
mmV2IY5y59imQ+5Ku1LWLSrkuXQo4X/RoRYTDMhSlYUm+hPZJoAnHqQPJUOSHLw8TtUXBTes2ERx
XLs1tAt5eQBESIPo/x67j/yCyFOh8SZ9kZcJPfi3D7ikOoB55JmOgZJtV61lNdv0/J7ZNRyQ7jOE
bFo9+k3VSgaEjkmeNwsifo4fdh50ZW7q8/SKwI6ckJoWbiThREmQT6w3TIoUUuV6mrOXRwp51RNx
JO4rpVATKjM7brRWlp2mH7AalJj/kq8CTrnlcIRrfaOGBeL7uR0u6i1Yx3NuO7XrV4GP+He4B9SN
rFwSZ4vvuBvhiFzjmVYFzVrjUv3Ew13EGtaYvnsu2ieSZg7L0410TifR4VgMo1ia3ZiJ+BiyY71N
wiQm0wUWzSvBilH8/WTqTTpEMPqW8azt2QPL1/3f1ni6R05/JQHmBQPWK3Yb5OxwaLFiiplmC5GW
orKJy5YjPFeUiVQ5ZQNEM95tC4Mz07nO33QRbJYI02LLKnK3fVcUIJbBd0r1EgfWQIb43Q+9Q0mB
Q6Syri6hyucXBTGE4sngf+weKBOUQHTp57/EK5OT83b/+liJeRMJSERPDNU4uvcOsgV3/bl6y13A
eGQAJ75a7zPe60i1Cj6tM5dXB6VZnw8gYIQW5YNcYIERGoEnWqGPUOdvnsYKp9pcya95+Bi0dHtB
VOSSJvj9XnvMRyJU85x9OZ+jcGK+erD+OB+oy65dODLWD+U+bHOhi8qPJiYWYEPOXTaSHfym+eBt
sENdri9SlQ9+9hcL5xWtzeoo0FpKV42SOalvTRM2St5UUH47V8z82ty+dadE3xm5v+WPUn+iN7M9
EjDt7dY4jDDeS+E/w9ObFQdrQp8agQ6E7KgL+qT3LIHInmkVSi88Obg5WLyyv3rQ8CT+8k0cImqo
s4PvoOl1KBs1qXntAKgOvvRjMTrSe6HrP6v0Mxcsg69Tsy11sQSH0rW6x8418iNvR1lyfXaT24J3
JTuiHWjIs8qg8TbXq9pUubtsRfjhIpcwNAQ1nmpkj5uPR4ppq2smtz+hEf7jUMG19Huq1p5toprK
JoFavcPLthPoOCNlZFjUlsMnVyS5vHDNGbt8XF0m0LaOBz3b/vKeZGf9LzFviH1AL4XvAQuFtLNp
to+6klwlUokLVMoq5AYdXkeVQZBP9IvWmfMSsw+IDGAAei+LmQU24uGsHLlcOzpyXi9UTvK1cqSz
vnZX8XXFIpqlrYplGYv6Z75nGc6g0Ug6wsy04l2a9yLcTUyh47FvmNwl+/eF2P0rIGcCytGr7okB
WJXevIjOflZNq6FY7KjBMeNgt64z7JsDYe4HXWT7Sxe8CfvY9LiH5UqNnt62RbnIW3Fghah3UKqX
grrhcjRUq6PLMSFrBvwQn08LnhRysLIyP8Ka9T/cH/Ep0n7ZRCWeaUeQloe51ZUbDeU0/1EfBnjy
lASG+lkFYlLaaMShlI6cVEvG0IyRNU+naJ4opff6quCdQfd/2JSxESVKQKm0n7yqvczIT/azkVwq
59rE9ffsOc5P1duEGoidMznyusggHRWLIFZixs/pWWbhegwQTZuyCNPU9s24oF8HMuaKpUQANiTR
QDA7C+/rj2Cg6muQ9oQkNG5H8HoP9kU+YZf8Ho9nJc2uMOVfZFs/4UflL8CyO7nKqpoFKWbJYBut
2VtP0kGsa5ncmKnoTjzX2bEk4cZQqIdyLEfwlRi6dmfRJJBP30M7Q9Ki+SfONv7HvEbcD/u+kGko
Zmv60FwnWUsmOE2F+BWAhsg1SpPK9pTTQxnp1XzBvNLaFCKvwnQ5ZeKijNfrxCIylCWW+wjXoUXs
7i9cCakFP2tQOscF12/5Axs0GLILZeylj5GDqokhxUuVii7grbqFgDI5pTqpuq7mlFYjNZLxeXs3
8SPqYBPfCDEUTS75Y7Rg0ya3nLfDzDUJYrDm0vHko2APVA+RNMA8W4NXi26ZkhHJq3ENVS1AAqFs
exIN6Ydc83YtQoBe1NwXdOp3onnxvOSNXFgxNxdDNSjYP3RsLFsJZ8Zp5TLig55vIneIsiEwKbBV
b2GKGMM1dY7IKzdKjidJ7JQDFA8JhjkqONYBb2IL0xe8Y6rVEoQ0xTxf66KeQkGaEY++N/LnF5Bk
pnXEb9ZHh+x5uC819NGCWyJZSMn8IrSnuUDWrhdtH0vLCBiLvZ/V+bhSwkL7BVxnWfaPZkLkMCIx
yGpYsYtM0YSsBSMQXPJn2ADVYhFBz6YEZtlC+tbZaJ0X8n2mSnY6Zaa2weRZXVSI5dr32rNz0UYh
qHCogNE7SDM2NYzBzuoaIXRdXrNLs82mPnxSDFHHGkQQiCLkqbzdLGyteT9tS5bHk+qzYshTrdVI
awHfGmDs5CRpn1hUen25mJ4Sy902LB0HqHzpXMSq0HUfvRGbaLALhuP6+ZwyUuW3E6F6WA05vdmh
RnCt0i27pm2C8/CT3eYjFuSUVgOfYxAGuZYzWwmCneDGWRfGiuVZOZYjJpXHFLQeOGL+12TBvKgM
9iM7hC/Dbr3jn54RSTWB+FI08RQL0WcYvWl9rlsRZW7MRHZiwpqupOG4dcGMQnkRZwbFGk0Ywq3d
3B/pWlwFQdk6zSoV4i6pZ6YPit2NvCt57YPDYi8O3vp1ZkDTsDY4BvwZG9Tec1LaI7i3Byzrj7j7
tdESQpvYt15lEfzLyFwQQ6PX+js/lVAkKIwSpESqu9uvUh/8+VA/WUKElQB481d7G7VCkvWUYkvQ
8AQiG+2y44inr4eJ7P25aLEpXhARzaKDgnokF1/qzPmhhRLIztfcxfOJCXMJlwJViwqUawsMHY6p
Ym87a6+M2w/0zdUohpk7KaqU3J7Zd8em2x2NaDNOBJZ7mDd3aEerJN7eJY7qmX0wMQ1KmQxoxMCS
MJOUUmRa1kbXdjrFQVDHqAmGoW8EKo9RdiK+2eAcTskjxfFKinp/RvbTHRNIYs7GbrL07iAEYYac
0TkL3wneJ7Tipp3x+t6SwWWLzbMKRJTHLqho1w2VAPGJQ1AQbQhzfN+lJjXmIZMa+Yk51zMgiKhL
skTFab9AxChpCjo6ArSt3XihZdMbQfQ4T2n/44ukdpL/B6OCbCMec22GzkYGA8YGidAetL9xyDED
/vWf9Jlj123/xd0hDyMKaOu4Gytf37+pTWlijngc0jBKKvSzE07rDv0vewBl/2QwRcOpEvqJiQKw
OEGP0sS1MgjicZEfFNkqf6q2Ygydr8a6HewXqG6F2YHud9CWohxYyR2YUPpqUI2kKDiBsq2CTVnz
7vXx5BlOLYMcHsxc70TmC6FFAphVskm6HcBJpWadVcuZEuw8hvMfOUGZGdUbt1CHRyLSrPLKz/qX
YwLw9+pWhUSBH93kTFCt2wa1+YwWy2cnojlE00uJd6XH9EvDmd+yC2A1R79j8fbXZy9joiCoiund
BFhnU/kCAd9o8dZjDot3PHAUqtMPwBjuzbF7gh86i2Niw0ONEqwbWfVTqUHAIZYmQ20XX+LvQNfw
88RojvI2Bm4ASrsauCeTEj/LsifooGdcHg9yhfsvQB7g+AMi9jIjZE+nbDRU9G29Qh1egC8eSMUn
mB7IJdLETEQS16YH9tum9B9+pRJ5s+lEPAtOibGEMKSiLO65tzLHPmgp11DzZnIi/3Zr1CWD+YKf
18uu0/7dV8NiKjo6NyqOfXoYnodevRDDwAZjQLc1KHKeqAc9FC27SmRemjI4G5Q96z2Z+MUPOIKl
o7pbkoJNbKyUa8o1oHgcCBAJ4BBiyDXtv4vaZ4Ut5cqOxv/9QqbuQoryYgXD+/sRtOZYWnU+UF7+
kwo0HwK8diTA1fI6mUzELdVfAvQ3m74WfC0Jj42pffRV+PIOiauaYkYemjNXSSKXiDEFsy97W/vn
yaOxO2iJwvvioq8YStWDKFEyTSju4fIc8Q+KVOqO3E/7DAhfUboXtRklzktTzg9kX0ibaMXPy1oK
oNXHp+CfqsCBpN9NLrRP6gmmzlcNDLLHVIwu6RvispdLy82rhhgWHysFIclCeVlSlD/Q7fsxIb4J
RbfmyweO1nZqtiRT53OP8lxUSQxTdrmnxLShc01Q+vXTYmG8txPG6mkrph97jzUE5hnChYvK2ewd
SWd9HES/YRlIzMbB+8I+PEUk0GTOx9HKzfvtz8rBywHUs1JA1eu97NwIjTiUex4xDVD/jStmK2BO
uKpN+XFyLh0tOgfUHPAhcknJeNGuj452G4Jy+/mLaS8Z8sTEXYrT0CJJ09QIyOriAbUeNXQaDIY+
PdGK6KbCWZWmM5QTgneMvQlmgcV9/GEDNMizcPPhP9V1BsnkB/mIlPxCBwyGK8omz8b1f0EPJeyg
4XbeM0MlaTQsEIMBJ7KLbrwO6RC3uJYtglEDvQGJh2J56E+sgn9S74WelXcHUJLQ8eGFNlp6yyoO
BnkjSPCIG5DQlMJoTNb1UuhrD5Ggqf4ws7GOPJztef+9gY3JwxC7SKt2riPpv81Cp3SBNVa6WDEy
am3mKXL13cRDKOTh90b+oNL1k6N1R13bNfz59DTo995Ue0YJZ7F3p0ZILeRDsfENXXPpiDjHGfkr
pxFMdj91zo3hAjLop2eF/gU9zfr/4c1evR6/a7NC7k2wmYWvS/eN7B7jo4L+z9R+xD8H/Lck3Uqn
6CPTfR0aTMLhvfCxrHdHNf83dcPvefRpORjliKcpGdkyW00Led9xqL5TLMSsGxnqgIea93AvOlXa
Vaz16Vn3j4/pFaUAz07ou8htRos/2MdX81JUHwpKjSe/UQ0Qd6E8INqdSZjJRxyZVJTBig12a74d
8/p+PoPfwV/6JJkEUgkNtUpxnivJPlBSEVqQ6eshVAyKbUpKdaDrFxZ7tQN9tuPSM/Tx8njvSK8v
1YJ9dN5RjBlw389W0J3K+dQTFirGaPWfRoPCSRsTRiE1QfH7VllTJGpKZffPzruqhYSbE6LWKL7+
ZkwQKOwfCeCjcZ/kGgC3qEtXGq/keYUZD7ZqZb2YEO5lZC1TmQW4EyIEU/PN23YKUZb5Ls9ntn2l
bSmhkgFCcg9yPH0fO60MVnWm3OfDnf5tuzvFeaVYKEjMlB2yQtDvwAwbCwXDhDl4eb4SYhISOrmT
YbvgBp6TTjCN9MpnQaUBjC8yO36DCp11Y8tQGi+1es6hAL8Nm+y1ShWZi2zjkduKxg+L3O92woDP
Lj2of38Ag2Loqng9CqmedeWGInz/ACYqEm5BqNoa2CY+lwf85EjkUMU+BZ8lYvkga4d8GbAZgki2
ZFb3ZAhoFNhDwBPPzKAXoE7dLBAT05FDlOzWZnnTqZ8wBHyOdv2K9GdkQYZjs+kdYBdnH4ezkyNA
1aC4SG4neYhUB2HvescBZpgkf+lACjHyjJ/nGJ9qjjIjL9G0K2BcWrD/bPkJiKegH1FDieaSGX6t
RskMlcnCxmxL5oxxZV3RnwZWnDnZ4dX25CMBlSwpglUK0+3QB8ETR+fXRg6pCS2aX4zeUQ6IpjO0
UaGYBU69Vuw2otCrlFzyWxuHphYxy/aBNLPXdGKfYL9VfAAnACyoaH3krreinjpuPRfg7P/nyDbP
ZYdbv8iJT4a+Lgu2YAPRjhIb99vU/kZJ1oC0NdnBmy85YMAggd2m1bAsv1R4EgoHl+LUvnpaNhgH
VvZh3kKqDfF+7c155AYKw4qphmn6nvCzAuUUZAkeMwE0CYVPzF55WhpqULXOa8ib9a4Z4dbyCE0h
iE46MYkjdIyNNm+uv2jNXF9jdRvBsvPEj5mN3NTZAW2/ilrBrU8KgV5hSrFuxC/nlLi/Y8vLaJSZ
lSieS7n8Dkp2ngDA/m69UFHflQmRfE3/Z5guJ1zkmjptP/IFvE9K7SeuVthcxf8rSWReTlCWtZpF
r/XgZHmTMkJym6fP/xG9afhWxCJQi9rvnrx/0MCGUS02zpihQBXPPtXUo6EJdUT8BbyBCrDBGXeZ
8V/ic0Pw4hUdpru19fCCokbWUl/K7jj+a/isuVCs0hTq7V1ErUnrU0rZaT8fcJFfjk919+Ob08/6
ItMO1TAvOiWDieuJ4gSql9lH4e30td6OIIrLw93dmgRB+RqpXN1lOfLHsePucWThhzUvogSUDQKy
TV0Wi8QeZPT/d1Yn5Qv2rqG9wOTr3aaoKP/T/OjNhjWhK2lEx+jb3P8j4uT5NXrrF3BzRqT4Xf/e
CMd52rHwXo3ldvh/vJEVMGI25Fb5sNmNDCwDPsksZbibeksE8qR8Z+3sH1lqtwwxMq16mTvGsf8B
M96YZlJSaAJzlvrl+hukB3FtGWHWmbVPGsUiFYh8Bvc6moKt7yFCK/nKAljlfhmZYdfA/9+hItIu
dUBtn1+rtcttcRdJDKQkWWJJku8U5FyZ2SGaM/Lmioa8cnJcKKoZX+4X/ploAMqIVZW2QDJ4z9Kr
g4xUUZrwcLPlgw2ZwocZMcD70esM+MKRdxMZvaTTXFUM+jxpq/olQyzTKwMfb6KOnfe/9XLCFVeB
yRCcXVAjwILNz7Aq97vE8bqVb1BF+ypRGkmkUC1jLYuHuFh49D1/R9PA/cTTofID++OVXnQNGgf5
McbJqmzZfUJTOpynYUtXaULNv7Ygdjbp1vlHxVcy5S2r+5tW8ZH5IEw8ZPU95Dcm93x77k2qn7gX
yizOAed6CIYxEFcW99dpno/7qN2zZrm5zA5ayuyJjWQVjg54lYZUhDmOrWpJAAw4FMxcbgL8E/Un
jTe2dZ0Mb7smwBbaOkoeC11hNmIS5/y8Who/hfPbmZgf2zmvYm9Ug5mnq3hm2m4iICsgnxbh9MPV
RyfCFd8alyniDwsqoaU9j2CB1SR4GK+E+ys9kWv2aDE9pby4nqJbXb0MMWmeWtbzrpAwGCWXoyai
PXQWfs04ffsXaTrk1OjDOFPW7ufGR79CZjDZxXHeAyoBpWDo7l5cybj3Ta6TxCisRadLtncIJBmH
RrRoy+Icy11XhwXorYfoK2DX3yCUTWgfpz6jfpVvbPkxJSu6zgnX0JdYbFYhOEY4Q0H0Rm/qPyPR
Wx99QpshVbWOf0Sne90F45dkx2Ki3tsxWYjCE+0aRgEsyveyeodfAr5R13uUzERHg7PkONFvopAl
0uM25iHvU5OBl/TeMQZjfSOIU7ax1A9RO/OE9vDI/vVingtsMudB8UPVZgEKd7laKTO4QskcTvWd
/2c7fqiSnmXFR8semETEkOouv4HY+0Fbr3pmraEOlL+EF+5Hy0x577nrsdSM3TomT6mlUNy7ZXAG
iIT4JGXeq4epAHOzjEGWMuW+jc/ZH7OvkwoyR/jLNDX2MuRCfFnJMAOBcUHPVCEkrB07kNx2XH6P
f6IpFTFNvm9i9Dc8YrLjnziOz8yA083sOnxuyYM4dlzkS3icu6T5QEsnoKiTKXTA6gC0HyToMoTR
AKkUmhNJa8p3TG/1v+UjTV6TapQVnaW2o1Fr++lV11LOz2Lu5uFZ8tJUOh2Npaf7HEkayXoGT3gd
nNIFGZ89bwwqDOgXv3rC7tD4ndYF+JqOWD6PCR/ZI0W90QmOJ66bdp/LSmDp1vgfno9baynjXoHW
F2/9srT3LTklZb9EUfO9Qy2besYjhO5AJeB6j6uFfocMhKF5s0g6EQgNzQi3SViWT0wOblhiIT6G
0xIASTgAQJe1BavnFVFYOiR2DtBd5lH3sjHC1CmAgBGnUwypY3gt3Ni9A99zYOpJtrF46XseLyik
laEZftiRh+Eozi8SD02MyFs/mZlIaSN9t/KCk9ebNagVTx6wFRMxXpq7daR0aQjshocodCArNnU8
LjiIg6MRMjAGz9aQ5l8iqe0EedLxKjiip64wzH8Mc4UYSrD9UvcQmZ0hdf3QBMoZaY/yPfKF6SHc
ottrwWZkaqQGKOKYGMFF2kfQu6xUkJfnjLK8EjLexrycTuK5orFPHzHJaCvhQp+4qrHDAp8TB10j
+Q0lX3xupdr/6iRkgLwWQMLh0MdAuLBVGkuAxnEVexQSmamkigtad9wNaSa7PczrlfFyQP7YKOo/
HKSL8WO10aGGaFauM9Mw7qZB7d9YPb2rf13KexEWadD+W56Lp8wN4OReywU63mTgDxSsgWNNiAsd
PJXA5Lss85lx5zhtd4xAZ/D/ukJq7iSNiEX8oFZ+JHCltRS9akWO2k7FVCdvMuia8JmY/sHzO9MU
cs+LANN62/6wn2W1xwtSV5zxfruatmg/refqbPpvXO2qOGGosIwjCyM5IXNpnB1ifRL2YOivUI1I
Le1xUabrFkfmYzrSEiYKbfP+xgSqcK0c7PNnIs7Toil7VHIv9ulPlnIZvwPv9C9ytJHd5hwpIAeY
Nb65agv83eirFsp7/CuYaTHWzdjS22q8CSXT0g5M6LqglRQpz/Ma2lh8sCg7z/Kp2kxRYyBLmxgN
0K9avhXNVPga9PYmFgp8xYkqVK1Ql7APwZZ3useN0ZxvNbd6LpBC/aB+9BBR/gGGWiFDxtnQttDF
2EOrrNoTq1D3QLkTIxUswG8L7gcjF0LTxxh318I7g6lCUId0Lb4lZeNobRO7rYzymzPfliem4fTl
BbOfpBXncPxHSRzb3zVHQn8hhu7xRJuJZ9HP1TrIa41W8mCo6pQUgv6+kkS94ntdsY0f4CNGOh5i
byTSvYggkYNqbR/uLWdY/ns33wvC3XdqeefygJACwQadNR3wFWSt1P3kSsZYTC61MhFdhJQD3GQO
8WPyrCeH1ETW6joPgYvfjlbBG3JlFgkAKGJeaHQG0fuGLwUY3CAzqFQtzE8V/5QnsUhUX2j6Gliw
7g9OGL/9C41EpJlfD+eSULFKET6aJhgfQNjYf8rwtUWXmS5cufJzV/SVQaJxN2vztSIDbDsi6Ppn
stowZHxYzOTJ/l5zmfBom2WgCoVqArZq+x38coowxsxaPArMkXfiLKUy0Nl7jVZREWD5Lw9MpGKy
TETxUScf782gAFazQAGWjxG3Kv8A0TkJL6JGp3BDmxur+5cecGhHv05OY7+GplGhKSInNNRakwjS
XuzlalDF5JFy9ImCGLH8p4bd9F+R/O0AS/XVUsIM/0uMvnn3L7DZlbwJJbR6k5bcXHKEPqUR8V7b
5kCL2eb/v0nGIHNjwjHkXg7Vqgz25Pp35GXTi1ApHyWRrnXi49B++oXx5J74jAVQJMGiT+FajE5g
VFiUT03bzOgaeN5T3DmuzR3q32jzk8RrHI+Pg7h+zZC5F2tehWAJOwEGZV4tFjudU1npBIOIgZay
oN1fVtsD/DNHC60k2JJfo6AkdkVzjkqB+smcW/HbtzCbp+sq9/Rs1jss0r2h2PkawePItBfD55Pe
Yqy+MngTSE+SdMe0V0BdA9JI60yqe+X+JMGPUNsb5QgSY5Aw/sUAKF+9ImiUOtXFcBGFQ7AQXylB
u/wXEh/1BlkVw657PyA/kD5fKXpOFXtEb9vhZSuLBACix/nMd7CXrT1DXsvYrYKAMGf4QP7w7kGj
7IyAr7jlfTaNW1hJhIprAuSK8M9uG1Fec49NykXnS6wjCm4Y31JHjsysu8b8lGGshq0huT9JRT4U
OdKFGW39bG1BWB4krae/U91WIjua83sKD54ORxHVadvrC1UeiRNAStUrGkARoBlJxzs3fr43aGJP
bwxSP7EeUHY8pVX0wRSkEVSO5ty/kXKEhpa70qTdflDhq9A2TZH6UDCWqDtcQug7H9ZbBnkQBJ1a
M8ln8uD1rGiKxc33iJ5PsgaEXcMp5mASZdALvAgQ27xNNET2LPETkAcK7dtUh3ZB71+6UPe9i8L4
n3F++bTE8B9nywCSNHi3yj6YHo5syG9abPrnGU7P1hlSYCoH4sVJ3jSsdv8T3TRmBkgUnCBBfkiE
QlrnuS65xyJQwa5LxURKzVYybr+g0fty9owssPWNiwezrtyGQHjr3BbOGy5KTtDnu5vSgeyp5aBY
re0T4f9Il5RBJM8N5uHFuobqdOm069PbgL/aYEFdNXrR+HhH4K1TSpEAeQhpvcl8uqsmRAv4X3bN
NeqfWTpiUisMWIdlaPzWMPfe7a0ZbpSyY2TPF6VwKVMYjNXA6JxOVJQetwzuTpH8kDQeq/GnmzOD
0RrbGmkzyGHaeGIYqTJSl64/lxkc2reV30HDv+y9DrLcv4IP6u8Hcuj9kDqe/ZeH0o78LdClFUQB
A9QKpQk0XTzWxm4jPJ0Sn2XPJ2SH58XEvFPnYSYdHw4owIv0YB8Ty2ScJe7U+odyko6WSuH/JAPq
YxEMGhD3wpav2QWFSsuaDyUcihVAlE3+ErLWtEHJGrUvubcMnC+RvnyBJyxI60VDoHczjyK+0c91
WY5N6TzU1vZnqZFirk1xFrtFVuQQW01htq12yOLQmFxiqEwlsxM8s2biG+GIJyqvhOYRzI5vfIU7
OVOoPQSxXuozZ1rst7Hs3OZfRG1TkXK9XfifYmPHTtVSLxT7OlJ7bPa2Hmh7ZOF0m+N5WWWEiFHK
lTl7WPRVKfZCAVKnQqAqeTVC7yXxGV4Kq0MRyjvlpFOcofcujFxxkGddMsdf+m6LTelT/CTwXJ27
qydUZJpSrsP9iTenRZz3u/zlyZG3oG6GLVqG15nsFKwxR2WVFJ/q+cukxuyyZ+QJ1IvieOLRNv4T
Fe0omsUGqD4L4HvWNJNqtrhUbsIq9uNl8jd5G9KjLxekEV3Y2V9Y6yKV7WubO4nS3Az8lJ/R234e
HHR9gHLmX+8acHs/JG78/exq+RIjbSziAyUBkTdHTa6+ZltmBFwTrUvCol04MA+KAfJIkaoBVAEZ
O3+eUNxN9pTYniDI0LTiE/Azv+0d/atLLAthRXDWiW+MlsmgDAbbtzjUMfWpzudTB5lhI57rXHs0
x7bt7qju/0yl4XsM+4q2irnRK0gp1YhSzhh7GWBik1O5pjsaj0OvXucNkNEGqYtpEZSgYClFP0hL
76+keHkMl7i9VQ1mX2vX7qxFGE7Xwr7DOAtAfERD7r6wk2gvNbqBfCcZkq//GW9Vp2zBI4wFHwcb
kziqW9ykcLsHRq748zXb0LxchapmrFBCTFsZcHfsRiBdSTdULandtEQAO9EltRWTabQPJR2b8rGI
AYlCqfReo0y7ovC4bhhCJW69drqcwnU52ACYMzAmuZ8CGv/ue0GtKQJtZB1vj3cjZMqD71UZz5aJ
C+Ct00uJzDtuhA9fthql/pczzXiu3/KBl4220ENe5DLpKdfGPXhwpw5GbGAsmvqCxri0JJTsbz4s
yLwcNg3+JUOyybuZsdV2ufIquGN280PiyxT9Tnd4+G1pZZVsKbIri8ybpaXlo7cShtmk4JotrcMW
QMpHg7ZBwNZAG3NXKsrEJI37rG5RzHUcD10/mfFs1TqaMhHrCL/ZPkcFq3487TLCCroLW/jMB1zj
bfNO6G1op248YsJHHXXrtrdLJKbu/f7pq+CnsLGjM3KHFR8ZToBFvMYZu4M7aNdqSiW+7kcSDK9i
Qdi8OadEUU+8iQKi3P8piLxyZOAJ4Xvjs81DeGCotKPS4Opy9yR788WDuhL9sYdAYv8A90OHK3t1
hHez2vQvmPcm3Z1Ty0DuEeU0rnWcT6k0rZfasBq7sD6gLjEHx3Zgh+fHrVImTzQsaawlhnjNKEKV
V3vrCnq2ZfS+c4A/PkqrB8f3GMK2MJEDKtfoPXtr/UEOz+yqMLU0q7FGKjWoRD1S46AqgjdAOpk8
f0od9QkGV14RFV69iMxRE4c9Jbh6VmDUqxw6wlqLbneZJHfLl7+ldmbviOcty8nLBdti6xvOvRAn
TQJYPk8NhI7ynwcNrSBzot4Qa537rUywMDYrhEihUD18aUdqIBSFWsvoJT5Uaexfwate1siaPGtG
+tngNnliESa2V5mV7LGZRsXwL5/MeV4aqXLDTIFUHlkX5JiRcfKYVMGBgZa4Uy/2QPxwCm6e0WPF
JYXxqauwcPrH4e7i/51kE+I7CtzzzSJZmYV6x6V2Eh5MEeV6daAkSbXL+VZfkskT+nXpKrVGpP+B
udF83DWCX+bfhEzQ5xUiyuyJHtZJ7J/4kI33KzjxLoIRD99yFdirFGnoJYUglvlzGxhSsZ/aAn7G
ipwFNnb1vV+dO7hc35ZDkN9DiWqI1ESl35Md7NoD9+UCgTWyw92cMNER8cGVOpaEAVtGst3pZTQZ
EMskKfNToTboLbXFF1o37XaPiq/gqQC4BDxIY9REn0neG+xT/wZp10/ZpruYNhiVkuZKQoXh3QFP
m3iVAg3tBO7o8zkI04ibFyf0eCQK/LsUD7HEtgCWyfRq37ghvW8qLA/BlS6H6oLOD188P2oGftuc
xdXQjJKGWMmA7jybgmTXXlrzs6F6h1YcMNBBtqtl6jV6p4DXE6JIsf6f0pXSLmrEWHw7xFmWIn7A
30WuENsaB1ph1YNu94TGJNgeD1QF/Mjlfnb9srmwkGOCILkviMifSba7ichLGNDJtmzRyR3VAY1e
Se0xvFKWi1l6ytVeJUnC2R45MRsW1+P9Oz439eC23PnSHRCK7/i2p3e1ae93/3AMY9ng+7pkCYDj
WCUeedFPT1EKBjOCzJKZ8AA5TiXyT/yotAjFsEKQ9qoPEDqSM+1XF6xtIEe2jb6bsE4xNiZqldRS
c/y9zrkMTry1+1fGrENwiFSUYLAihXYB28utbSXK+7o1qpJgWM4HSxayMZ5O7nKmq5C8IY2Oe1d6
kxLFKVR+ea229eDgAqDf+SrNVORWpA0h88OJdHFwZR9vvU+hmv49+AGzm4+HSvYelAfbCnddRTXn
PopDWj8WGMU/303kMgF5qDonB7TwxT0cCc6kxrn3IQ8HRDpprb/tcwqwRZGb6rvGrZp94fNGDvuU
Ip8CknUWnIrjBJccsdImGjYC0kkaEoTtRdwAc8FDSlb0HQ0qfU3NTYsRP5t99YXU/rgKz9SsMaRk
83EvFBiGWLOE/qEUGkZLdgyWWMGbjxBgLnwedqKww4kOyl4buv2l4jSc6u2Dq/aA9Fkt3ZzVAgee
LIUQjSlgqHSBcd4rbOsFm7n6ZwWFOixmx0o4XTbXbJCooPrThQLiYyCSnAZW7D3nnUChCeZFhykE
9L5NlGJfbRI8Rvq50jQTxy4UK3WKJitgthyZgR8Fr8tJ7NZmf+tc76F41n6ERuZrytxcHSmm30Wb
rl7gM5H+vRWaU3ZdVEryBZFquEabHX1TaaOgZAl75cKdm2tDyWC/ZaTzeEd4+VYgQ2PcZzapZoBw
Tk6MDg+TZ7L8rT8yYXRtCsaIWD9jtSqDte+OYRA0/DTPH+BC7Qj18s5GdwY210wKTYkzABFW8QvG
JYs1ateFsIbk8dJMyMndUtOvVanyfY673GvupXlgSAlehc8DtfZYmz6PKopbctrkfSFk6BerT39h
ykzLJAily7oyAdv0y2//k4yGwrFa5oJfCKiWRwUyKAWahjAUwcQg2LE82JiDOWIq4WU17mwpsWxf
aB6TgKAiGSVGMV9chyPrdkLTi1LpkDhkOLJY3jF5CctrYhJ4P47R2h1D2QTSfjfzNmyT0a2tLMHk
0dmXKOhE86zFSct0nHPigZjoAJKiWCemKet1KYH2q1OKGG2bManUtdhjPiS2ockpkhTgIzhaE4e/
wTrMH1cqk9qmvpnJH5vRAoJJUmaw/jWCzWwsnd9BSOW8PYS1BrBbosqjSDxUm/+DSCHUKlqqo7CB
dVv6TgjbYPujEsWd1frNIif8UinQJWLAN3BoJ+iM5APlBnHrBYP1Pk6dthTXMoSNynjHdTIm2n1l
qoOz8Q9Y8Naba6Ij9ENsz6qOOPZL2UueoSHAXipg5cKscUZG52YeYEGpgKZdOkcFBcEeeXMOlUPQ
DnQTQjJ4czZORme4XKoGCJI+YM9AKzmcHeo+PanFDwRDdnM+qg+CWAnjYP4GAQuwK2Ff5R/3Hsak
vUcnNUzS5ZB4ITjU61PrKUvPmIO+IOzzdhBszID4D5GN5HAn7ynzjpyrvuZbOMtLURgqBN+YQXhS
G2kbn9zyeTtQ9kApEQ8lXgznRiB9h9CyCxBGnrdTpd1lqcTT2sTyWuetxLOPg/Q92JBJn9d/rp9v
JzyF2G1L85IfV4y8W9TVIvAxgOBq54/7iM+N+hflv1XCXz34FrdafD5/foUk1oSZMZCWhY8fncX4
MCl/iomSVKT1bQiczWVrDM6rzTmGJJI8eK9KNYR1Et9IODBZRtH8wU0NFWfQAvX2PoKr0zu1oOPo
8bCu/IpDR1ik7qXji3GIxcyNFAfxjHPMNr7Lv9uuNMd9GmEL0gRzYG6eTjA8Ibh0SBL7RDCys9PZ
eRW191shjI9LjC9k/3NLK4DWjJbOGQa4iJxYWknhXl2jxInG1REiX7OfwbkDX+KghzJrqv6A9Z0h
ndODJR62Cmzv2idEz3CkMgmvsmYBxpJa1A1PpeXJHVp7mKyaS4HVHcijydsbIPjrI3cb9WnX8Gg1
aEAz1ryPxOUzNH+vMs2VD/xHvXiQAGdRX8ZFd+aNy18V6bx4E/RQweY5vicfXau+rOyRVPUnfxUH
cUFOxTILWYlOJIMv3MWivd/QeE9TC+GjIjM//K/5vSYqyz4PeQiZDfhMFuku0p6ePh9xPbW0YoSr
8HSkMr+0Nid/93Gb3vHFXJuejqHIlKPymB74RPOIzHY5bJN7mnMG/ksyhk6SSLf/GRr+h9Ph9ZDD
ohiDHTCP9NjSJvmB3yY7LzASyPwANEgprIj3NU2lYHdgPJnkPtQfKP43v2rI1HtxTgefa9OdA3VI
D4bQ+SMc+ZmettgRkeiRWO7s9RQC1KE5yOEXDRYdLLeqezgpcDj1Y0fRW8vQa/iPsoA9xz++KHNF
76DxSSih40XulfpLTWs96tiFJzoOWLPGG1SqS21dOjbMQfdxPaQcWnxIs9o1xIRQC/opU2N4oIe7
qhKu2z0C0FAgVlhkc6mngPRbKI9Pq2ZOLYDV1xChsOFp4OL7Gt066qEEp2/2WHMXILWaV80CuO2y
NMvbDRjKn+Xrd3rn4/aKXyyUX/JUWTsmXibj5hsE//UQW0ilMfEUj1sXc6Q+n6zAIW2B0Ya037G2
Dzrjo2u6EYiSNwBiYrPqxcFIARss+XNZMzxhf0P/nufypjQgHef7PiP0omxjIZCOUuHWWAasMULK
pJioylhf1PgTKqLNOU8EHsu7OQZvTaCqkhA/6bKWnyBhDGPA7hFr7GTkrY7P8WwPMR/OqoklIyVV
CvdOwVa99ztkx727nMkUcigG1av5O86GFSmSQvswoC0zNmMfPQ3TOxaBwKGNQGRNdDYx6AvpanEq
jKkFI27t2DZigYiKY40GsrsQkfFoFEWJPUNF+X5y5fCtFONATOINYorSS0DGu8H9onFdpQ1NrUy9
Z6CLRv9hasH6aQENVxjLQ6NYKMU2OYJ3N2w0MehlsFhXzlTr5Z3KlSiPkT/6lLGZ19k20V4VVWSG
Po/a2rlGHt1uiyGGYMOCz/Iu0cyH8Jzt9ks+kBEaQmreGdu9vnTqDreSMs3HAQcUG1od4XJNGxLy
DxQbDQH5rKqONMA6nowo8IBoXAhZb++wld7Z696dabB0uI2Q3aQL5piuE6TNpJm9oPpIC0wO46/O
ZXC/jbE3x5wpPEG49BLvaDDoUjwcGA5Y6swf7HGBMTsZWAG/U7OcJnS5usBYJ3u2hZLa84QwgftS
mBASCqheFAm8RvuB2i3WIsfLDBlRPDvskno0cpuo3M8ubE9NLjwJrLvsdepKmswx+q1Fhd+4lfqK
FrofSiRlGI3HfzWPbEwoWtIkmmiEuU2zJQuP64qwcpa2wmfRMGUzIWtjhs9TAMds+R2dKL2uLJb1
HZD9gP4wv+dciUUV0TMUZDWk8aY5PQdqROTEYrJ6FJjJ/kULdsi1eGNu2fN6h02NsE1n4+C1AdmM
0N6VEfRfNFVsBO1pJdS3usN+3kVaR9LDDmfM2lEgOiq+7JQvAly1p6dgOc3uqiTLLVdRfQyGudtq
WVQFA/r1KTDAOZxdSGjPY2nNMMldeQZdFUE+wX8I1WjdMQ95ZmfRe3jFATn3qZzVClziq89dV/jZ
daf+tANzUWgsa0WxW2j7262hJQpO3uyVFaXztypJIHd+jv+dKXfWT7K8yJcn27OCaTQKq/P7tQzq
pdjB73bxSqjhIXlVgHUic94A1cCcFY6gLT3m78GqK9IhaPM5dwVs9zg4y4om6fyKwA0b2SZ20Cfn
uaYwV6B4WqGO2VVSDvDzw/4D138oytegIpWvqXeOSDSOla88JdRU4R4hPVv0xh5W3ZcO8TGd7DQO
w5JYgkkKUNkHMG6Xvhp4+mugL7Yuro8RKyAbraX4vv8oz2s3IsH+Irs2GpRLn/ACldtiCPMVcoS/
vb4FTpZJPMNB3OlpobUMlqWDATmhIAVGwX+l1dlNLM9otwc4nNJ3hljX0OlSArrPVW20lC2KNrvX
ZrxGQpV3NVFsk3UW378Q+y3/BSTL0Y+C4MloBahksTW5w8sB2cEWwY3mpl+zp0rpTDduiKXI0I9W
vIG0AQH7Sns1hIK5KLwCNL8E5xUZ0A4VJAjz8eBBs669DwVc3RSVTmpnpcFP8ONyxeU6yhxmxhoU
e6VW/yyfVZFJ4JdpzVVMGGmaJL1R7d3tgfd0QG4Apl3zH0N5YN3MzA6BUhWPss6sLl/VZ5d8io1B
7DYWMHpHBx7HQCruGC10RKHEwHfoxP7oWH6klo0CrgqJaHwfKdKySuZBG8fFRQp7ewUzoGFbA8fM
PQSOHdDwiQkRCDONmhlB5uBtS902zUmBOYqHZoPU2MAMOx+G+JEr2AleKqsnCbWg28Ypmp3ma/qJ
DqIKhEk/rJoEo9wxV3XJQ8oEeT5LvRiGLme+p3/oqKr1exhLWLJG1Aw5U+Qf1D5kP62vimh4vRLR
ntBYCteIDmdcaxcLzlkpuheQDY4F2eLYHq3mu5S9xXkplkzn5o4vEB7NNjqTDEGfVDoQnE/gvjc4
697xyXshGKgriruEVsOpEjvA7ROTegQCJfwIVX5XYRpls7olayuW/TmIJitvDyQ+/rEFBaDrW7oM
jPlSQG1pY0886DUOg623yGvBdB6XqK7VBbirZjalpvd10ltI0JGj0L8+lCoGhQNyHQX5ilYxHk4X
E/uHzQX6oz3lwbQ+XKcjue8hbeWUJAZBgmf8xoPiPenLbV0Z4dzhqRVRDKScwoUjZYMcqB1JgIw4
gKqZfrblSmt2lOWN1u9mdQyAt82vb+bQeciMTyd9Xqzt/qOWavnbwstsedAbz6I08XZritapWqsS
JT1jEKJKR/8soSh2E09scTcZ7rqfLxYzcIzwWxRN4cn16TDuWoh72tHlcIsDWoRvjFi2QbRgQdI7
u6FnfzRHCR7/muDGI3YkLvbaiU9MWD/rrTF1J3fC07tpRzvKtzSQN5ni8f3jLO6xKHwwqfAablyl
SuOZXrg5p+2Tq2Srfl9jyxEwh30LTUsn0RRaHtSJ76DlJs+aMc/CGHXGXcfuJRTMY6G9Nt05inra
jcMxhi/XyXmilNg2YjclB1ZCC/7/umFWljdCQpd2MMxflicAjo3LhKiLOTcFCQPZ10TnfoODAWkl
rzuxLPR6GxRNddWjy52SqtFa6ps9h+bcNLD7trAbH975TNZ/DRFmCdEMEBqfWe1Q93u57X+AwoF2
xw8RzO6TEyp1u0KrDXGKcDwW1PhifNOk6Nu8iNVKcAObGavETw0ahaFHxbaa+vT5wANPevyihUEo
v7QTBRDBRG1uF/yjNY70gUtMxCxpL7LYeZLGpBo0bHR8heBsd6+0zBB52c39RpG0xuxD3uDmJwXf
hHZFGN89mmsggJuNekNoSOGBWIj42746MCNqVaUtpPV+NN3zu4ln1oHzo18jFDpJT9Sc+oYg40Zf
UzoIU+jStmrYETzutPs+6HvYKgZRxlFX498Z8ggZqGHz9amwqXalv2jRiJVbJmoHwuQc36ZvIRT/
9eN9xkSeIsxycJm6RBYpDI0d4HzQ2iyPcsmAjVK26tQDlbvhZn2vBrRf4kA4yXOFgVsgcHDL3rvZ
xughikOc0LBmCmvlO0G/pFow0Pr8Vn/EeoxL9Wv8GAqmmyC4U2+Kl5GQlx1saXRz9ezzYJBPP68v
DRbXxsiyQxXUmO1L9u0Ibl+qsydtqZdkksjMDEjnumOWkgkh4gpDclU3aQTrpoCQR8+4kjyKPmGf
OvBuHIYUqTfj1uVnb3ZJ0dph8KZFREAh7JNhzxGKdVmtOENumriWyU1rFIw3J2DP9dLMUpTB7KRC
qEdfLZpdE1N/VInBIgKslCP7T7leo0hl1Ng9Fmg58ln+HVSB69YzLCYynKhhQREhqHM8l+hpVm14
WrlOcVsrELToNZDGwoKJ5+XB2AMt82ZgIKC2ZMtAdRY5B4n4Pd/L3Yn3jF79OccK/XtteIEFZCkV
KTRwvY36bMJn7rKUD8CunGU5zo/EO8kZ2GF7KCx/lJEpuyaORnMnKr1SM1kqYqOP8vG1ZiMiIQ3c
ohXQ+53vr5GV0tgIbuQqNtoLxItIg8HmwfJjfWCGDdjbivLrDQFc+uLA9EheeSp8GrekveLj7VeU
kf9RNn3scZow6ytz0C7pvj6mG/tGvTTiIm6OjrH1aDqxtQWXckncTkcFG5/cikPfGjgQDE5XE5E5
zSRNhdgp9W4Xig5jWttFt5l/dPY28MbwTsY7PSCUATsYYFhoK12cCx4FIVt5aUqg1NhBy4Ac/N0W
vKC+UsbVIEU1sax4y6hdB0IYmeOvB2aCKUpBqdcOcHKmPv/7fsKKtlFRqRpDMbgxCwg7Q/fXslVl
bnhcW9JG06A+j0uu5mRSorTLmVlgoFvOM+WqsL7UzpDouUh2II8Hb95Q/ajmC7AB++zKxbI5bd89
UMwmYoeSaq6xrDG5K1oTRjQKSWpoMBJRpRx+i6TQc3/gzDrbbR6mSOPF58dOkl5IfM8x+hWaMmAR
/X7xVxBhHXkdPuha0EBrSY/p+K8SBszbiFm0Z2JnMOJaSR/45ih/nh+qcjjFbJdFK9pxop1kLXb0
canlpdI2YDJi7263nXosvDA5U0QJLPBHuw12tGQwrrLaYfV7Kyluge++hzzUBSUPvX0eSOyinkTz
C0wE38kA2NcTlN8XOjoClgxAwizqWls1FN3MM5LTl09JlD7TUQ9qrd97flF7pQGFdfMQAQjeLMm1
Q7waeyuLvT3i4CM3N3G9StIlVDt4BGHva+ivcAxJXtHw4TOzTivdQ0D87+bfWgaroGBzz99+KpPM
hXrSq4bVbUngNE6rYvwz5ePH0XhWQxXolEArad/uo+20/eLJlp2BEVJVsCK1UNwN62GKRSzse4o5
1vY50mCDWMFuYxrTIBbsUZSCtKP5V5K+UTnpYSTNZUpgXiLyV/u4dzOqf0tbfHjjyjv3/Kcr1YI6
2HJgpsehnZ2ukneGWtRZ2kEUNMzlWAa6J+SmI3JQ7PyCJpzxpK3B6djsnIpnoyZa+pDVFiHbEt1f
zTeJ8ZtLTYiBVKy6/3mEEZL4lvb0I38A29ATfQNPFgG+UyEAFjHU0LCJpELPZBhvckBJH4MGRePJ
fWqct/YVxKNznwS7+o9Hx6y3TbbipuYc75YOMJFMfHL2URYCFC6hdNzVVH0t4qXygcigxjbyp0Jt
FswzqFC4njZxsTaWk6QBRTDSqSg8Vg0fBgHEvrZ4ozCIR6+qHM1U2zFnzEj0Y+5MjALKOlZeBpuu
u33va+8JzTxnIoMorwx6sgIRcnvQCHu2U2qdyn+AfxJQq8L4/sB3HszzzQOBdKaT6FNlvo071BK6
kTXn+MA/XQYFMqbnE7C/y/CMcgTMT7hqU+IBtRPIywWqO7BqZtyhmDOtufb6XbTwQxKxd2idcQg4
9xGbbaX39Au8dFN1laAi5O4IrqQTSGJMfzpE+4aGE7gvMTW2bQfMfq9y0+Pul73yZ/d7S3amfLWd
vY4LOFs8AH3UsCswUNsmFeqX6FBuaL9/m3OuO+OtOvdMnn993e6KxdVZZzNDJZm9ZzX++fX1zDUM
1akMgSgwi07hUDPD1nxe4cDEmooRVbkbX7Pg5b4rG8aKj5dMpA+iquxCqTSRM4fsCN2K9GoO6DBE
HpUySqALFXuTR9eE1I8fHCoJohG0hJNfHTYfnJ++tG/9XdOPM11KGzWE0R/n68r4umzzU1fUqeuu
CqpfOLXWE6BUp6+lU+4bFqJYDPjmbk6AGJGja4jhkAAgd4c2WfSdmE33Jo+MS1JIcrz86aeqipEi
TFVE+Ft9pdnZnkl9rRtt1UcFYYrIIIBSNTTPUIN1SaurEW3KBWlrvKHUCHQ+xUv64afQZkOQzds4
wwjAYsO0MyGb7GEiOlXz4qzydKLYIIOr60Ib3CSvA55WZiy5D8Y2zgtII8tNaXvPVB/DLxIAJPaH
tjbMhVOMDBkAn+uZjbW7REceuP99jjR8oUctwxVkNKo/lF/nTNRcYDA0mwMqZoMGzdsOimhzDq5e
vuSu9JrHqyV6/d466GzpxaN+ExmTaee30paSKw9uVuiDHghcn7uN1nMq3Z1caR89CTZFsOgFo9PK
8f8tz7ssTlRKTqwjgECIJxY13yiHiKeiELa9pAEbR+umIac6umRX4RGCT6rC3udGbemkm+hlNE7J
099c0fRNN0ExqF8kevS0D4GQM+zIOcE24MaGMzlK/0FNX7YVWEp4anIEJrLi5evRHGFA5mqYRD+R
i0gnxlXeYsU9V+CpA47y1KQtNEUnQVsQ0XTkmhJCjZZQUBJxq/brftJhVYqoxYTOIbPj24mBoDgU
MT6FwPLfX3JZOQILDoempyXdIs3tsdeYQy48p3zqdt9oZfI3Op1YM9JbTAYQZ1k+0a55MSJceV4P
vAUA8ZWHDCxg3S8iIdCMDtxjDWBV7BXIqmEIhQ+oZT+e1nhMGYPLbSdx7iAVx6XHdDvi0vcn8gfe
QG6DcBzs77ORkQvuY3Qp5wS5K0F6fXy1iU/paWa3QcgUv+qDUDFCVjT/5Y828hc7zFpBV/x/J9rj
XqXELIwqWjGhpHIYfY7Bbs9YsV8ezD7nPRPBY2BmIUMq4eQTPUZLrF7ZMt1Iom2pzFuyaY+cgqFz
3RiD0ZX13/hhY+1YiEEwpKcAWLyNnLv0oKQxmcRqtL1u5DsFXSeje1fEVMR0549tUxIdoiElwKYA
r0mpiKepiVepDL4IoqI4uU09IQTSzyEYXB47e2wjSpItfjukM9oChvFUzXchzCDh7j/NSGOmgtkT
wL1CQ916uhXOAHCnNIxoDkxBjhvdcOBLlLhevCmSNJtW4P2+xURoeEuX3lwH2YrM8ZXxGEXEnKUs
ykVnjmECcTnI7uaKqzzsZQ6SUm8MZTSlSbVtPV13vpnkbxfJ9r3L7EU9lVfd0uQMBtq/Wje2ZTKb
zs0Fn5WPdQBsVXCQtaFbMsh5w2cc9OASmR9IMWUl1e0tjiHqxKLvONPq93cuKe1Amz4qT4FpEIBK
HDjRlb7tQ8XfDUMQ9E1z/Ejr9ULvcO2UEpAHcLmnVgi2LSfwKLTpMn8qTWVLQwtmcZTCKRMNFthH
x00OPhuf90FRDvnWjsWlani8c1TruLKjC6wXSLTQVCPtgX4jBP/2C9CnH/1I9ZP8DTnDQ6fr+eJc
LjSql4ZKaDJMssAfGXtdlZQNljycoj0lNFFoN+vn6AW/exrVggFf0KUndh7kVJGI77q4Dvxtjqkg
VccRgNYSGb8cR1L/Ycs1TRagesMa1gFCxzs2aypGhcowyzwqWuU5ylcXHyWDhClbLmHo3fK3Bnnl
3aTr+FLhSgHekEwhbT2DoTAjBIuy/7oIx3Oa0zoOMiDzAEYyzGLyLSc+KMTzIXa0cpj5dBM+Inb/
jlbN07fTOMDuyKdzj+sDDPEIt2uy2/2vh1uT1ZK8BnIDRV/6QVx+nhnC9gQ/M4vd3N3aJ63hxTI0
0sCV4yBNZpM3lPnRfJK/mi86PsX5IVoi7urk4vD8MEVs5B0MrMXqQ2TJvv7kXrnYbYeoszN9HMp0
g1aEQLaoL64IIKDFLJiF789ofwnWGAWbC8Vm5WL8HWM8ZOYkUml+GW6t7bcVnro35pkVcg96ajHf
H520s9KHXN5Z0RTsqDT4CspM2KEtIgWbBsmzJRdRU4Ai3mnaKK6i+zxL005f+N4ydhoaRIDuNMZn
jluA4xzaLg1gznQtSaqp4/o+ydF9luDJBVpOqPtdTltsoUjNyn04JleQwOO0ixjsyxlSb+kUaC99
bSL42YScu4NUduUVSb3jlbQ7EIwt6MY2qnQNdJ8U55oPdogVs0qCEDNsz8+EiLtfFQHLU4Shg1vf
sZ0FpFEMf+Jbu37k8qiqf6db0abjponE/PF3dOYkYREuFYpYwIQlipaKLsbinlu2w9gUD+kGphHt
YlREXMt+ujwCgK816F6NZeMPyWDp7ZTfFqEttyvBiRR0vdAH5gNPYRRnunqpbGknB2tfqhOIDdQ2
qZDInYr8bUK9mM9BxuxQ8oMeVOS17zFSKHcLVFM8Vn0QY+4Bs2KkAB3toISIfVoyZWIL4cg9pEmY
ch97hZBoMWG6rr7BFVtbYEsdRaAh1K0k7WbmIXtx4BY4QbnWUuWHN/wD0Req+ntplmU2VTWhvCbq
j84O1e/Ko8djOVF/UoBxPc2f5yGLoTXiz6M34P4DhZnb0JSHE3bI4PcHp7qdMeiB61+8PkeM0Puj
J2u/jGGPKX12VIQnZkK+4C28UaS/uzwo6uCiz0NQBek/H+QXzVFau1N9jezxJxME6GaZ46CHf7uG
zfus+EFeUHVtFCiKalzm7/+lw9Z8CxpKR8Z8p3x0XMkAP+wfNjIv32T4VhtXanjGyKkvcXFPLoag
fYP02S6nk76qHk0Zy3u1YNPintJU3oUbVbnEb5MICcYjogsICtjYo/Rid2mRefT+UlRl9w5zP8p5
H7awVsRFg+fVG81Vzf9RnAsgLmkKkcVmt+/xzGF0fztMUNgLThUiZ7jKT/4Qf3iw+1NlFGne7Hr0
eH4sRyoAy4XuZuKYmoQe1j6mMPFbVOY+7PrX9Idy+z0V00nMqyYTaJ2KpgCXrjCwhJW38c8hUqoz
V510/OFoJ/6gZHDSwpqZk8wIdmUHK3XMI0U0Y2W5/hse/LEoEu1Cb1R2SB2DYkJdoajbS58P5I9k
wkcDz5KS3vIrcsnF8a0Wv2t9G0VYwOW0lXtnMvXH4RUz+PgZMN0a1OY471mRAaHRvBQp1+/eRFmZ
TFGZF0/5al5Umxc+wwyFA+1a3JgMubxIarKhXzGjeRkZRQdWh3SvtmlkE1g0Jdxli3NX5tJnQ0gt
Xv6GBuurQmNikbU2FmszAWhDf6mVvASIt3ljlGJELbqJROHTTYq42+EEzwJYHjF8ikPEQuNGYq9g
hx1LKIkoUfwcrSlXavDT/qI4BKchfawVCCFQur+1Z3Dq7sGHNd36jtuwx1TIFlVi244mzuNDtGC5
dcrYbjP9ibny7NN/dsXPhnurmxrlCH/Vb1WGhm0Ay7/NIR+5EOzrA3OzWrLh++4FtTjW6Z4ebDee
THRLib1DQnHlI+/aPzL3XmZSQgR3ZCZLBrIAP/j1b8eaNhBJMq7IKEPmkF30KJI8Qq86J1lfM1Ii
8HoGzBAPP1C0jB/W9qFO7kRueoSnboGwGRJJkVJPmDhKILNDgClH3i7CGhlTp6l74s3cr8uB65Zp
Qt05LfGMfVBXQd4xxUZugqLDiUE7uXIyfYhL4j5qhB4AFIo83ayW5EAFpFoF59u5J409lE8JxPSF
eMIeY8baDK/cf3wCYv+BNUP8tfm2pVy0iKZ5gvLPDCZej9FK0CrlmPpkxmNV/K6r2kksdI5hdfe6
xK5zWp2tqjSNeJc8kIm2pBBCGkzSFe4OynSIa76eV5DQs9eBYdXe26aDc1jk2MpoI63ADEYbMmTj
1IIWHqou6gVgjZKmnA/sO7igZXzYZqRENC4wYai/LYoUH5nHE12QxCMK7MyVQXcsz9JJ5TUy+gsA
ewStQUbswn6x1hWdNJxyx1PmyAKWrBSVncGkf0mo14NeE5gaMM6S8GHG6auj9d6GYUnem1nlqmLi
NY0mpetf4fa1nEgXJfDQUAqc4grbQsiCaqzud7GNJvFb+YAARprtSF/TF2TAW7GsphwWdsUSzvNc
bYyFsMitn8miL43FYBKwY92ngur9EIv2ABIbLXj59UQFceomZx2IvmwstXGd/yIgx8Xn3Nl0PZ4l
yUhwiPMPqX4HDHieJ++EL9GT9fMgKy3ukuwS6U+8k6vWbzUvtuXsDQysIJDF/JCUST3KLy17dqQz
4+fa5IKwnFhoeV8m+bcT8VNfl8Ha3Pw2bysKbql61yphLEozSyb2MLU0nH6arD0nhzhBUX8VmkId
l6+CNwtjScCjZrskyXN6jXL6dzfI6TBvcUlJifWbhrc6Xc9P2OpAufAOwp//TFGcW1v3+LGUxL98
lWEpg8yNoYCrjqHw1PrS0XxmpC4tQ/7+lSGo0TUq51+cHOtRblHWMB81YmSOQygX3PpcPPcD3fst
6Papi9F5mjT7lsUdO6PdEVt2SJPVTiio1YK2akslbcMVNyJu3ItUYa49+lQrQKA8H+PSJga7x6En
O5VvRo6HWcLZcYLtZg2VdUIjpu5k//lZElLSqTFDfySOcgImwYnQ5g5nMN45dTioVeyImYD5EzcC
0x6z+8xjf9DiBeKNSWuGkgl3AU1jVRh0T8t0BorPLJSZX72Ej6d58Z8QcjaCxxpFpjFCBScLBxG9
9a2dn6PhgcN1VDQmYbu2Fh4Romqzj5TYbm/1q9zFbcV9sxVscVavxmVjFO3FdOpxL/LTDB1MYy1D
udbBv9AMjgvJqpZkCPvikrkorEZ3b9qSktKl8ZxQ2LmNZJ6fKbRLMTGl/ldMZlzcBQTcBt097T5Y
mJZ21h2nlVywh3Sa9j/rCKTEfwb2AqXmbXNlByFJJc92wOBg/OlpbusYLSuArXLb9TJQ+XRuYtJ4
tx2K9mFQ0OA+8kBZdsaijRzj9h359czHznft/RJe++ZYy+fg2SxrFRRqhXSgDUzYijU1/8FmUCTU
/o3+yhRo0tYCoIfUvyeV++nuuGN+WzdZDWe97RTDs45YPrLW+hSl1An36Ki2WB9fM0WLkqiQ2yAs
yMG4pZTIkxhWzwVEr0ERlmR9x27AOUsDja8+3zkx3uhCFa5xHyGC6Udoicxagbfo7et9fUe2Ic6P
S6hayUpYYXSd0pAeoneApQ8XzeMvmXPldz7Q65cUoM4XNyhQ47qxdSDJquy8CqOhdyhsKHvbL/vG
TUO5+/wrkvXFvdzOPN5dAj7ZVSCnlBRF4MoaBMO6CjuJcW/sYSCUYWZRfLNK8pgnXuB8T0YmOdJQ
mGu1NwHtYIFZd7pAO8Hh9smpMiZNXfVg8PhfypsypOrRr6mAUAKdQZ4Z6jS12izbk/R5rJ6Ft5GP
HYpBabf5sRyHwd+F+IUp0QTqJb5T6917pvL+xDxoXDdT3eA8h0lpBxWiQE3TAvTov+7yW779SIDf
XzPKbPcGIlDYdcsGxQG864cq9OfYsh0Jc0agfYcWAkHv1c1sRB8n80XkoiYiiwAaFz5oIS7XbTNU
pHSjoOLjKE2G2eECt21MnBaPjG5UDynEsLuFFi8JAlYQIysVQUCF7TwvnWgdyvMUoUu8GkznQPkj
ej2s+wYe1uKQCARPwJn2WG4fE9sVsA8KP7F4OY3Gi+LZYDskqfAyuo7JM1/uwUjwwiidNzsCKXab
Zdbhq0iNIS9RyE5QM5BVLZK9WzjAn7WMzpjzN4HrRxqvHXoZkXt7lMVOg5VuZO9o+FXTkhaL7j/S
yEgSjWfXNaZkZ4up8EXo0KeySjBeYWepVMvFk0/vK/1Ie7pWrZ3r8KqviQ50F2BFEXb1ckhTdmpY
xr1lIO/baN9KjaEOTxK4cGsgHIdqQ2swk4FMtnneIBLFnFG7jG8WhnmsoVRSyBtzd1omAZ9039+U
EZtA0U9W5NUXzgKLVwETNx1+fEFStOuYN7T4LibLtQkif3zb9QZOMPmfQj5BESajFSG2JVTHGB4Y
cWTlNXAgYzdBrOjzmaVH5WtNy+tPUQooA3nsHQ7SOY10X2WtVmIQ/H/aH8AeLsrstarQE3r8jGGp
cXrzc7ByvpC7MXfEgW7UixXti1B7J2xtUy5pKQjNNtUamvmlZI7ptkTwRLGYfk+qwYJ/BshBetHg
yM1zFlkdQvgXPctTUin1ucBwqFxstKPt/Z1PZL3hO8pX04N2PX0Au6RH8atf1tdSgDwSlbxQU+ek
CDr9vnhsrEeVbz+Y6Ly/CRqo8ZvlN+ZqwamSiXQyd96nFQsO5y1rV5nz4Q/eqTokk+mqcK/3TCmb
+SeLIs+SYotjukoHFzLseoVWW/WOukOwXg6hEf/PGEBZ/AE3mTOLbgFmwrCj6ruHMy2cJ13MjqeR
v+Gbmz3ffVWGg6qe+DYk3Cqp9lcVi+/8wYROVgI8LAjcGOz0Jv6ndaBJPBgGR9avmSKza+3/qTEA
6oREpqqAgnq0aAUkjfsudffqmKJDQCQ9OfMuQlKxmz2qnoDXuFxyVCnBNjg3SM56M9TzQvUwcbFe
lz/kpKbSjleMxIZjW25sIprO3sNEPzso5yEuk9uxJejBvc4+UEWWBrMXbCt0VOleXsWkyvvPJAbb
x3V+QILUH7gr/XMfgz8j2lON8WsEkmgfNswFNi9XdO9K+xF/J/yRhR0YseSxYw1X8KX6+wUtbgsd
CLfS7a0PH8jhqUCBWwgWfjeEeEcVwxuvgjHMypgnS0HoJf4tkgUWDSHG+MG+yxrZwr5F1flWpVhS
cytXb64KVyJoZc4bHgE5pMJUGlpHl2M2dc/aroWQ55usEYHC68xuj7QHl60zcHaMzJf4JI4e1S82
JDgY9eZbXdKHlaBdNWRl33nvEjBrVZYxIYdTJ/W9kBp85VcHc8CeCAww6FOh/E1eRDIB2LR1Xxcf
WBuK7RqG47IoQauQqEirhMF/5mZYtYFjsuCNDIbk9N68HBJrKDjgnJw9ORIpAdP77fMfnx8p8r0c
hMwZecVR6s5cR5469Des03HEhFJx9c6AhDA4cAUoaeULX/UGyEK3UehhU/VMwKlUGCdMbxDJCTxp
RJOcC7O+3wy0bY698Y1Fjh1i1+2dkKsmLG+DSnXJY783uCBlJ/zqxVUQBxrh1o2QWTsYKvMQhNHw
0ycUNv/lDpuYCInG3tK/iUQOm1xWTqk5n0p8Yvh0x7tQpKaem1hlOoiXCfteAf15zo6Zp1xhSwNW
aZaDKQM9s8UTIgGfH4rCBolMKym2840yn9jwciMhUSTTKvdK01TdNCuoZglYmYhatwkKKGUUpCsJ
Ws9PAopZoVWC9uycQNNLEML2OVX2widWaysf8B1T7MCuQt6J0fsCKdqiiOQgF6ik4R9R1OoWr+ix
lA4ZajrPuKiiCIL76q3UeTG640ur5xVTRwABK5TwGjbN4j1/h3C/g+k9afvl1FujJhS/3HAtLnOc
Ben0LGAvMNJc1ZDPFk1XVBEYyGsYwJlaj9vr8jpjkYSQ3G2b6scaeAhGQuW90/0rBcLOebuhn4bM
Evec5bnDP69Z4Bi0vTvV/4SLB438jwg3JzrJQ5ZrAqFOyAE52MmjLK3uuz3EzIjZ3eq6PGTKeFtj
wqwWXXlqzzzLEG0Ge7sdzBgC0HpqyYgVxTeXEK+sbliTO/gqGfmqDVm0LTaplEhHiV5a9QdNO0L4
fpvkgV1qqfTxdSiLrzvV4UNcyo2EmKJr9Jin1r65+Yudhb9Kkdwe6TkaRQai9vmHxUVBjXyc5B9L
/lkS3bRbTnqE5S7SnuqsbVpw5T2iy0Nr2xUVb9fGJ7nBAD3fg1fxXmLOZe+s0NdjzLmXy/B9wO2g
nyIAl4uRJJizF11oI2R/VvnnaGaPcBSMqsx3LGL2OV/dBuZBB7YOYeiTYHXSkXDc5xEnDNHoPg5d
dU61RUK4Ok7OgMVkRzXbyqy+yJd3ACp4v58nWlWF/XePVKMJdYRogtIqi3J5vhOni94WIDCVTNSa
D3I2xUERmiw0jeDS6UYjlo2TFqCzfCezVsLSIe+oy0yeRb91DmyCR4QOS401aWUBXldtW9Jwa0wN
v9mPKaI4aOZD2X8pz2jbAHC7IRXAC0Sfkg6L8v8GpTTDJnLrkfV7ZoTeP5KEZhKqoPQxrqBtzNZO
aWNXMmJ0/f3NJu7rnaBpoj8/zviuunLRsxfk/W1olkxTxf7javjo8jOcbdjM9xt7fkwKmZy/SEYO
hXT6QSdhjovVjgAzYH9VOlDc/x6KrKz8YierC9ltPA3AqxXNO4sxgyx0CVdpkRLFYbTi1cjA4M1k
gaf4aCSHFrncajdJ3kvOmf8oPtPT6oRUI/kxVE92FP4ygJnKZC+1Sgn6wkCNtpKh8kXXd217h87z
AOZa+W0UlSZUQUwG4Gs17ZAYMeuYfzRaLXuawzc28qz48QMuI5772cBmHBOQ75qQFygxKyvzlk69
VANH1M0bQ7T7YdbHru4+TdrhjDdraEec0bfi0Vu38pX7MPRn8cS0yiQrPS+19Jnw6LN1Iq+C+0/5
lTS1TnQwcucUKsEAAMA1uIU7N+M+vmzApRku4YaxGoW7nrYusap77G6Oob8Pzmjxh8Pp9LNnJUom
ReGDG+IMGqn/EQAQq1rXYQextswF+nXQIIu6jM/MM/dX6ldH74tWg98kcmLr0qgVvR1v2U1iSoOJ
5oj6Dm1zsMKs163NghVxoSR9D/W8lk4RSoVfz1sCqRi5j2u++GNvtS3LjAZYNrGdv0wfKYiA5F0D
FDUYpaVv74HmKfexffxknFFeUsOyiq8LLX+CE9kmrP4bMGZBmQJMtRuxlxjGutrMpiPFrohT7PNt
T7LRGsgzWSzkTQOT5k12CwsvLNJ54IrEMFwJf9J4W9mpNFYwxH9jyMnKiJM4bIB5rocj5ynbESNM
6WE2+iJVJkuX8/frM6ueVVXWObGaCUQvD89JUmzP+ChqduS7sYP/JcjMVW1IqM/8fYQ92FFVmuCU
4DccB05uwRB3TktzzwjYqhMZQD/Hhd6AVbtWpN5W0TUPFVxAYocLvq2GEBx+tO6XvuOdrH7d2wYH
qmZMQsB5f5T4NATmlbc05in4QNMnzqmrc4Hsef6uRLtxhP2Ywlc98+ndrqqfVlLmRSdlAjP2oZac
hQyzt9ZsvD+tmUjL+YaMsfdDNBTWp2zl4bdCz6/C8eM/e4JYS0OCSyEZCsEHlxRsRgan5By6WFZj
ZA8so47IG+qdc1V7t6U6/1FQsUvwZns4Sjwz48XJc6wDlQe5vR2zwzkUXrjlmHq/rwXqoCJQ9cxk
rpvbZPv44GtMP+bhsCYglixAeDEj/MFlXSybX6cizzj/Z6YqrRtOiCU/TRxOvPmmHjjnkGn4Gp/8
3vfcNjPHJ02oMjrtMJLFCMAVkpPgGieNA6n9+kkpUlmYiAASsJUeG9a1dOIDi/O6J+ZDx/nd5prm
AyY/IN6RArj7CcZ+c/rX/UD3gesSI+Txn3cb3+RGaoaCw/lFacomvWuxzdzo/h1+5nCluk6eOUpL
mbHll962uEB0yd71G17KczIGQDKibwqdGXmmR6yqAX82RGPZkxWgmtfO1O0UvLYBtb8EqLhKyzEH
nBlZJHjd9zXje/Ue8Js9QeaOTFwUdyueqk+Z86fyx5tYs8q/CD+trSrYlkZ4PpQkV+PfDbJDWUD7
6VRTOkxKA1STxI7gqA+chNLZjE/TaqWv/p9Lf50DvUj2bbQBxR/OpBCxNccNtqMn/DmaEPIVEazM
8ccZnK0KnT6hnXlO6iQj2u8ACmMygf0PNxf8XuhR3Z/ovHXbWZKdcppr45RPlJquFcZJW9yTWMoP
u35nKUCmCxiCt6TTCOGabyy/Ma2X59/eey06LckasYIaz7yUg/zKtrZMVTqkLyx54LEMim6iFr3c
NXBJBwIYA6QUVXSpO2WcgQv4u8WcfuVsEa7otf/TPXS0c5c3obpca/Eyks0SHopaIbCZ6L0OypoO
3nTZCWyKTp2N3ULwSmSFYWIkGxa1SwRh7M+UYRALw+Q34mmR1tdix/Ir8s64uHfY91FbUmO3w2pK
wNM7HMVN7mjt9kVv4vFwjlelKyxGGXSPVDLZl5tUebo/qmhfKEIwXRt2MwWJxeJEhatc221CdDYn
vI2tvbLufWFmdw3Kad3VOcabBzaPXXLcjhWJKxHpEkFaGGUriYAw1ighKFUOEi5DEDjY7bCG26Pb
rpXjbckIM/8/dJjJdJl0E/Pga8mqlKhtvCs6VzpcQEJ6oV4Xnl0DU8Ijf6L0ROLKgaYA150I3+X+
sTVp2cre3ttUAAotrhv5vWAs1LJai9iP6sDnuadqJSSvWueo4t2j7E5/M9QCToG5zZnL29sHLVKN
GFRW3jWsAi17oZOng/HKhg0W+eAET5+wbwvQg1zUAFvJW69ctfrKxftRvNaWp1fWTIoLQBGNPFnQ
ZQiwlTb4aThZpAy/zkReZKzMaRKm3Y3p3QRCn9kttqthkTTYr1oifFEajU2WieQ+AdF7y+YODp2J
aJF+NsiP4c4CUp75oOVo/jvmJWB1WBu/kDW4+haemN4L4FE20dpfpiofkFqMgMCuKWatTt7X8gxk
0W1/Vr9cCZf5GH6oelI7OHJx8J65RiYPh0XtlVODdjJcKtNYLqzSBjsX1APwTgrVbeHBW3lQa5Lj
mB2cTgBpaQhCaEDsrRPGhZHXRFXFfbP/Dpoib4Cf1qVHYVNse+coe1DHlh2e3MJf8F35Y1+G2+dY
HAFD7Eqfu3n+abiyKDAN+6ykTAdNDsG25H82JhHrwKZf2n9SfWM0BEA0/l5kUg/L2H/jfv6rJabR
L0x9iwrt7JtzwB2FMJsqsWkkMNZCT/spF5qAECM18nGYNO16DKLq1DiJ2r7GbwFw0GWMW3ts44yz
ExVo6b5ANRKLKXFw8QtumfyAJmdHVSznk1YzuXcqC9A5hj5tZbBGRvwNJ2MiZFUYFoyqgsCmrWJM
1fB4UrgLamP7f0lXUsCFGbJtQfpGUmZjXAabWJVkuokHx8pZ4BHgChTMSHz2od8r3vAHOQxBCAoC
0RM7s+QN3BcA/umz6J/071CVTLScuaLRN2KHUbjr3K9HlJL7TT93YargWmgJpK6SWvgg/EDqgzCu
2H+lHkKiVvp+EWbnJdIPp8DPEy84fdVYd0C+kIdbRAeS1/vNYFH6hSEqvuK5RFu9bnvva8Gd8ZGX
rav9mLmbzR3D1PMdgmEVfoTvdXOF63gLXWlVPUCUun6mSwYfEzgtUxwOTcTC9JcUXx8I6qwzaRjd
RLZlIdB2gnrfvyabqsUcl7IAYNrioTDhrh7dd1vWMgtgqc0wfBuPfvlzu+YJW6PDgv7k/aFJ63AR
EJD+Ya2SO25XsUp6aZkU10La+oo60MjMP6s5gbUVsiMCA9GmCmKqANISbwAu7+RjC17Abb02qQBZ
lnq9K8QmbjQQb/X9UIazjznoBAUZHgoWagDin1tQ7B5hK0yy05Gv+O4NCgbqms2kotx2bD5L6OJB
Y4IKn1JOiztduNSsOhLvvlxD3J0CcR5msA82jL5fqflGrArNKt+AmkEsV1wc+n0OtATg27+6SIFp
oiRjlKYjxQI30cSK9nwXGS/OsOxfK/skgzzRKNvD8plwrLVv1FC42xNHNKI5qmbwlCN1AP9tnQdb
0vQJ+QDcGcGd2nHtXmrnC/jVbcyn5qmBnVKVD0MetkpdgB6QY4Bfw+4zzlbkBXPnUhmLle6Z9mRC
v+Rw/NHff+T1Yl4JV7ql/qqyp2afsVeZlaTvrVfKTKD9kA5/AOSo2c22KjHtUKabybgYeqlWnyOx
ocKSmbiHqTqdAlOihaNLCVp2Mvov26q9MV90l7ze/DdlACTkXx2nChGO6cQ7BonUlHt7i0Yn9jUt
Yyyf+DDQL0pgh9HYGnwgAvmehKSgMJfYkYDsshUtJ+ZdFfef/IbOKrEaTQYgI9vb0KdlvByoJij4
vIudoT8itx+1G/yrF2Ata0uqXm0fcM6WDu2LahJxOWxYcDuLh8HOk4xtvORvo6hA18a7Eym3pe7i
g7TinDiKHaYC1ZUWF1+MzjTSG2GBSw2yAQS+VEfFC50YaNQeuSSQGDUEy4KK77t7XaLf6Bni6jvl
133V86RxSygDUL9kA0Sgkgd/IX1pAitp+T7ej/IYgwJDz/jRSFP8ET2j551qJzKRnRDi4SVEuVZL
F3IzKN/aJDUfTZzHp2OiNz0Lw4/GZjgWUWiYxheHkiiQyRGiB8WLttIRQldUmkieInIjUY3LJCOG
rnoAVIAZkhxcnT+5S1PoTzUaQLsWe/uT/bvg02NkFmLX8Rv37Qej4TIHCZhzZ6hk4PBnpL4nWryh
huZdR8KqTvTEY3ZluaqB9SrIcRyS1qeF6sOzDI9hleCUcBlqVD8QapBsP8nQPA2ysmrtyzIf33Gy
lJm/YQeUbFPc/Ifs9akOq7GtbfbHFhS1QxHizIjBbZQC6Gv/TTwBGGI7TPeJUYmH8R2Euj9990pQ
Ldyc7Kjb01JtcxAIvmfM6gFnRN9FbqRlaDjIiSV/zRKHLtstJCe3YTQ3ktMroK0eCn4nlckyRzNx
oB1igDWAJZ65burRLWehrOeClwo3J/hL756xN7yT1ILt8y3TakdrNTBiXo6eZfS2GPhEtIyIR+5H
nSVSecJC/gVxUD8IvXQAAIQwPfe5bzglZR26Ry1Dfz9V0B9jJv3iTOvAWHTHTRZBnEB4lLaP1aG7
c9hrygjmkJCUPHn7IUH5mGO5Vaf1rZ1UsDbS8A7GKPTSQ9ZwpYxjXne7tYbDhuk5RrD3IgG6DY4E
Qq06DiMX1Q89OCBvmo+zUVVFr5nQGvo78romakhhL1ZR7u4sEobVy9rN9Quv+mWYwj/IU6ozmdiF
oIjNkQ+KuYHFGONYggOog/RD3/PPNbnTIIPfdrBNNgi/gBkWMmZajWTJR1x3iQK3ROaxXO7tbZhy
A1K9pBs7AFSRKKOKNEw8fLZJwuk9vWKFzHGU9Rx6BvHZD98F/L2e8um/7pfXWQ9dYQk40fwBu3e5
Q9wwrxRTtQ7FSTVFN2c+QGDWXF9Jt19SSjratgQt0R1P53Ug1ZCqvxLCF/Zav7iBBGYrvcZWNaUe
dWz8RS3w470tImvAzhwoiaQD6dLhv1PHmQF59z+WtUKw9t42MJ+nt/n34rdTWm2SVAPhls1mhD+I
hwsc8CFkApafcvG8iAUHNBSEL5JWHnGWmA3BXQUjuUagfMb54h1Zzz+G8PrwAnYBlzFGSq0ooveV
zsIDUo/b49TAFKY+9oKFyKvZWcjgz7VPKdy8T59bp4uCu0eNNoeg2WVxWoi1+ZAKrA98kzBbbowW
b8IfUDXcDglXUYiWU4syihf7G8lzBB7RUdzye9spRnfuv9EKkjutCiJzf17be3m1JG1aL5PbS/Id
AY3yL3VSVOtsVM5eUzmaE091SA8qiiKYkTIvMaPKB3g0TjEUIJ5vTcPKUpkmPlVUcPCs3fo7lQYZ
BAlCNw7KuNdAddHariRDuRGAOjfaQRpBsbVingYU3G1OT7QOmDO+Con0kTs28eIg3ZNGMu7+JA+6
JtujQbHbJSxlbLcNgj5Z9h4eDwW4omB7hBjb1XHamas0Z+yFwdf5s2c48gMXyq4Y+TUW+jkNYL1b
UpRm+vP3JGEKzVDM7+z/s5xrn+HPzeLmnG4L+YgvGDMQRWBYuBxas2gGvZ4cL8Kz/js84oqcAsec
QGzWq7BygvXU5pck90J3fiKftQzAQhq249yySeGW0JlqIaFcGqFOvGv6vSZD2XolA5T1FYrZG7lo
rpmyEXZ+Ak/ThQd6gvUoFF+jRrCxU05gRVA3ivpBII74Mq+vXjch2iMYjlX6OE+ARKq0YHJBHE9I
oQu6GZzCfrHfcBPUEkxxUi4j6qIAYbzq+iNBlgIgJnHhToe94jlkYp8RdPXY1J1gmge6CVzgsmbj
pmGDoHGAbXmM7K/J0+IfBbjMxQhyDL1PPOZjuLZKuhIfCNC4mPZTEjw3NMAcmN+kZ5sB5lV9S8R1
FhqRBXTMr/4F96P+rjaJQ/AxiREZxn/jWN2YPkVnWyYQSHaEjgNooNBiKlgZixEbfoleMC1BPdg5
p/MbBD7uTVf2jZ9kgOwN+hqEKXdJTVUolmTpaNc6D4XKY2FRZRFbhMVEr7czZ0m2/SF7MVuKCGmZ
Uzc4WylVGbQuqFvecr+c5jff6Aekn/s5lPRLrNA7aeMmQruHUNwMegPIkmDAYKv5GOBBu2TyUgGY
2vQcP8ZzbenyjRuf+nkdcZyCcYHotyl8yw9mtRqc2+ES9W4p/grRGv5Zz/e1om/yHdxZqk2uvBH0
66DJxvhqWjmtvTK4B6iSqk8gDqW9Wd8hgwALtgqt+EgWCzgJCyBV9D1wtocoLBAYtLF99CsAzdlw
8AYCp/r7gfXXAqcQ5xskMcXM95B02Rs9gR0/6JzRKzJrTrHaYw4MaXDk1lRCae5u1M7upQNZTGmd
WekUZ689YKQ4BniaqbQwHlgcX0IQ2hTOmfa5SzVIW/Elu5WmPHFg3KyXS/MZM9c/IgMgJhRbrDI3
cuCWiNqzIhbiNTYvDLK4TsLzP8Wp1saPzbK4gFOgXt5Y3JFZsVrrrvOIyHbTGWb2/ydj6iNRIznB
CT25tDpLhWbQBDsu8g2OmFzWcYgWtZt2LVKZQnSKSdIWPIFkH4DfyoxeWYafPs9CBAS9cxBSQbRx
prBD59xmpm1KU45JWkFZSGDKxQkGQTk/L46aRomuEkEegSbVWwmASlW60EYyfEeaNExwqhH2jp7G
bXHAYEWl7qrZ2TkFy7xxYrorIjLXTPV2m3WRUz57jpXqPVI7l9/8zCASHxJYBAdFxEdJk+YQzAhc
IhF01/0yZFo7wzsu/aOkCS2vNe1UL+D10KiOnqJoWt9TGnypQO8iVuMX4nVmcN2qIHUIisifNKrq
aghzAfVFyUrBN1vB+qQn0FVaKUTnC6Fn0RIi49HigTgIFISb6D6UysTN5lCCngatOeR+Ai47Q+/A
Y2eu+y4T+cilrPVbC5cDTF13GkNdvoNnGMw0DN5XthdGRHOuW8lH90Bov7xrScp/qt/yOh8Q0TQy
gGY8OafLHdfV6CVUIyPmvxBV7QfkQvNmQgqxDk+13nkMnsZ1dNQmu0AX+kL8hwmFjcG9bK4Ef/y3
JbXpdvTWCSj/hOX7RnAwwiLD3hCzWAWZ8Va6vu+Fy04/nd215+Wpz2rBT8lKZIHL0Rb15yFJXiDw
SJK0YefIhbDuG1V5xo7hGvrWtoeSyzAviW2EkxuETpZ3fwTogsReMonnYeVC8ulL+7FUvG8XAgQf
Zgq4duhSDfs6cpFwK+ViHHyy7iJ6VsrA7DpQWOwwjTyZTPaYE9fd4DVkJ1LKE/1m8Dy2UX7utl38
zrKlC9zZUYeA8LUcnc/oNfyV5apprHARor7pdOhEtqMcZYFILsEm23NwqvCqrC62sTP4vB/YrP7H
DOF4ymsuCiU/E8EggVXEcLK5rwrHVGW0TiftNRUoxhL+cMv2VScwz8jVMJjttWC0S5WkROJVn/Uz
Aip6k/WNI9vKbemf9Tla8NR8OZofzUIta6qKhgglyQmSZG568B9sL5hJhpkR2WkCK8FJ68+ApilU
2DJl2P7JqJPovcMrr30Fw62KnEubYRDHtc2sLWWEPUWKp1yjhQ4X188dECp/9trU5HBuS+kyNG+H
SkAZYgTIcuvNzs6MzGeGOwnXEmOA5t7F96yF6hTTrH/NTmDuLf14Y8i0tKtes+GKUTCOtvEnvQdZ
IZWQH9N1MusmeQwNBz6P/WjpqvK/UDcdHfxeaPDyXutJzT/ol0z6gtnAJpjJZP4DRoxiCshey4Qn
HifTGJr4qh0N5egOWcR7LOCJ3UYrThXpR6dUoHPL1hL1InzEl4w++3QmCdHX8Rwam0oFdlDA9g/l
/xTRQzIlNm6Rrb3TXEcA4sYIJWBYMA5HhkdrLsAWjioWOChaAf+HvdRrq/gZeU8DmdEEv4x8MhFP
mjI1CCR9OwVbvEp2GJS8A+clQnNXur1nwujQZI5+phCZEPyxR196Fw24g/KlOg3Yh/5I7PNAtcko
UkOSTvc4kWBrPbaToY6fcUPD/zWL2V0q5odoomMVKMNSB3C9yArjK22iYKA6wKP1YVEcVbfTVzt+
bV0rCAfRJsd39BFlcZNID+y1SFGRbtFK0f1NBSbhtP1yswFctVWXKUz3jy3gAbvtwdL9B1FK+T67
MFoJXOS7JF0ugZwI8TrTqZd57PO1m2sXbOWd2fwyPbmEnE+ZQz+Of+ktit7HTDMQ1FJPpVQF9dcO
4BqPoGGnoXs8BWUF9AuuImm8SC0P3Tg69QOj3oyYDEJX8EnxPM57mq2GJZLZvCBsT/SM7oEpgKac
zsq33PYdvED2sbNgDktTdKr3nnmLKS20LJ+A7ROhNgl/jwqFCZKkKqYkpZja0VVjYqKX0dRFOuvo
OK428LrtlzpH/ELWPGcstFUFXcI4hPA06Cn1Svu5Vrw02Wd7QOTBTREwuavF17D3r8A0FhvndVtO
yYUgGMIWYwfmSChlC3nX1ckEg4uVfLqMyi1lclDZJmxtsMUhtZFmLtr1lFLk/KTCU/JMAbvw1oG+
RyiFLPSkAr1CmUHrq6hjF9SWl+DPrEq/dTnClQmRRdvCNfYltCawN2zhSaDy+CnJi3ttcFu5EJbY
PQ6ch5iarJB/xkwa6CoWU0EKd2PZ+EcgaQmfxLUVF26Pdlk9V3NnqaY/l1jFA2FnoDf7QDpjsMV1
k3N6SUjpGKd9lLI1TL/0aZPC0E0IOBD5WQO8luLSre2hkq6HTzXfy51/U3fGvwtgklw/7Rh5G13b
zUvvg9c0ZapwdgDbs7JQH12OQHQRcf1ljwwx5pJ6Qszv9asbKIoTElX0tho4IIvIMac5gyNBhXSz
WMBe515B2w/sj2LL7wmNWNLiincOP1Ql37URzyF1U1swuBeFegm6FOvhH+kL4LhrURKVk0Rh2Snh
cIef5IDLG/MCTG9sVY9X1EPpfOPEyPM4gf7hw9a1j9FCKYMufiwubZWAIkoV+q5X94rQsP077cHS
m+jbiCaWKpyVFzXdH/wWK4AoDclpq4bLgv87+6YTR1BpRlm7lvRoIMmFz8FqL5OZUJCElyfzPWVe
sqPL89VU01qtuD2Dy+6hOhNLhNHWVV6z/yCFuwrNSaq8+2QYwmWY4OsoWuJaR4AZWWWf5fQb4dWY
dP0IWG9c5Rt3Nck3iDoCInmgn9pS55VwljiDb8UZQCv/2ADg31+4gaO9BG6SiyRFqYgRvJyJjj0o
CNPBr89SrzigrVDbpNz8BvEIWMxHyfzGAFGEOe2V32clQ92CqqBtUQSj1dEhEMqZO2UV+vYmtcJ1
zrrTYSCWec5R7Bk652++gdVrVHn6T7BIFLfa2BiSCfw9gE7LXGRHMdsH6HolikTImBXt8T/HmBq8
bG0rWUEd0M64XcxfEICimNiSsEBAjr7laMUsiwQV9oq3hPqTtVIoP9nPZU0AhRZhmpNXrqwaSjDz
KsK6JTVZSxwfnS2CLHQboBxHxTNSH+wj4AXU+J9VLgZeJoZDq7nlXjaVpzPoqOLGQbeqyV5kKhy+
oOqhJPYQI0GtKwxmK+P0hzNQAdaXgF97Gl266x8jRSSFUQbSlgrnQ/9/CKr+qcVtw4p09evvdw7r
Mit0yuRv0rK4biNJL8E3jxJ1kQaIE7HY0iVejU5hNa+WdMAfW5BhNz8NAKa+PLno8h/Al/PVW74r
ytkFdTkBbdQynJ5d2rgnPhFnq/IHhPKWd35Msdp2xpLaQsWURCvZ5alPNJYddJ9ylXYo9WuyAB3a
XVii4Do+4DVl47xhNzwTWMZ6Q5tUvzyXatryEbZp4SEUbV8ger4PhZMRxuh+MRj/XjVYWQsR6oTO
JQXC6ln5MtB6+rblcOp2ov0JdDQ/tE3MfxBlpKmjs/91PyvHwCdtraVNFo5X/qJtPCqwuNUdflOV
5f2Yuwq+d9XjRdBbA8IcMkp6KxSN1F+qTmlmkPfdWQPOspNNs05dfFVZBhIlY8uPUOhXqHkj1+B6
+OslKxu3dyXTXUkM3M+CxWXswuZEbgow9bTooycmD87AuahMAoQSHOoXIZ3SAhhRR2SU6N5ysxMV
L0f9d8z8ypi9GIbb6ug0roCPdTpOxbf6wpoOYLlDRUQuyjYJHI8/aH4/eeIPw8Ooe++oBIX3JRif
xd2dtsr8Ocl2YXiQC8S9LmwItuTh5W5YqofZHYFOWlOUB08qnVixHoJ/8BSgwqQGsggA/I3sLAo2
c4fNqBiWJFxrPbkp+dDM0+6QJhmsETAi2+x31wzBMZq6Ftkp2mhSdWoCpKR/ZGEnvbsSsI1z6eqt
kctmUSEpUn0Ot9rMaXh32L5Bj8hTySak4+Yy8JXEpcu4u9AbYRj7d3oLUSUGwJ1Riu0FhkxjrAJW
eha0gRVn/tFsp+ZfgZ5+tcXchbICaGbkV6QmZieKmU/RnZjsiNt3/6M43SFQX1h23wB9cxKZiwv4
uESaxqe8UkYczqIIfmw14Xg90NxZxUVYrXzVaDSm8+OC2oInGFJl+pg9csRMv5L6IK7V8+6zityz
IPXjSYLDJhyYwAkQxFwagSAY3oACWeFN/2pGZPD0WMSk4gQW/KnUjIMVTGa8WMgfXJm424cPI6P4
ARjluBVTW24JT0es9XZQatSQ/ObK58joxL7LbxQSOKIPf+122bg/i6Sc4NNcWW+bNjX3oDEmgeVY
zJc+pOV5oqDhAMpudSL/jCGRVEGsixs2/H6RFgUok/C+tzFfxXNqZC3BwG1JwoX/U1Ei84vvdVBR
qpRWERVOFAkKYQ/PURblcbya2819fucO0+6f0Uu/V3+UMBSWJFJLJ7r3R22JpHpClQWt20opP4l0
SXGXm4Yhj4olXMtT5DqalM4BBzJ7OPlQJMTuBZfNXiLbd+1L8kdReLI9QqPAvl8VdlKwko1zN1uw
m2PEuHOuHXIFEKaJJlWSXt962qua81m5efjg8DoxDZGXWwS6soo6ngeS3oGsHN7QQOV2iGH70jwn
0/spLussOrmNf+MugjxHYlj6ZvJj4D+R8NeUAMV5d0f0U0f/sQ+Bx9E0Uk4xs06tmW2MG3eWoEWQ
fgXJjovmq7mct/AQ7TbFFtkp9W8z9c/w+8PJNnuLFCOpfTMBwAsPXpTjyXBkpGlcww9f1JTH9VrL
OKgBQc8azOEzOsgp0eqRqFUaRjLGkU6DZcNtq+ZSxv6Hj5zQUd0Mnhkrvz6t2AWq9bNnIT6SZQtT
yFFbwEIRT+da/FYrX+Lnk/bj7KoyKDmOw5W8fhvWBhWZTvUggLMZXsRCFr6vU45sE7kLSU2J0H2i
RA7OJ/Xl1lewdyhE3hkP0i2fPdN7vYBIfeuyf+Y9mxtUuQVKyQSXOCr+4SvX0ZY2IwPikDTURXO4
fLgsbxjIHJjjisJcsvst/E+CVwa97h99jO6DeRWZ5iEOgJAhfO17vdldc7BTSGPRKGVJP+/m1J3h
BqL9OrQ/Ayr3zV7Q05c1RwX9afNqi2RrTH/r6X0Q+UqLgW8XJDvCcHfxxQg7siT6bjrK5GRXadlV
5uvED3gW9IC0puPAW1q+PiOgS3ibOSBXXLMfk2gBo7EF+aCwu/Fyu3cjbBdwnHfMpaVwxR3nwUvH
H32slGNqt9SqaRT69ZLhPaddsMt41HXjai6B4aaBMuBbVkDVx0mJ9unp2KDEPvsvMja3BFpA6Nml
O30g/fl+lr0Q95OxgAJmDlfJZE4lKAphcMrV61yqpT5HQUX8+zHdrHINOvzHJHC911s7kA4Hpdjz
YPWqdeRiZV6y77BHe/ZbOFpLV4a/2CkeHf3Vf2xxf0mGKkEdRkMMuSL0kJYHaP12AAhZAdwU/4EA
DKfe4Bwxd7ep/q95CjPuHHSF92qQ2Pw0xkrZ3RmWfSz+ibxKoeekdOSTUukSCkVd/DhpH08PQcN/
KtBCTweitezWiU3vX0gDoIy1fLBzKfq67sZI7gbWkdy+qycZNYpA5hlz/gy0riO3s6sqVnXoubq5
iJMKBCB1jbEwZ4wV1KoNxuqCCa+X/R4hbTigqwB683m9/dm9RqgEZHkRl0dCJLwANIPLLp80neQK
twLwzYLfF2A766GamFOSgveHMu9XQV9pm56HsjI8PdikUmlZ2mQ0dJa4pAhXTh8dH+fEsMOMNRqC
nallstdzHsITRZUdXprfGRHDxxddHqSEuJh7tJknCesfKSe4/CxB9i7XHvuM0N0sNbr+bakdrA6D
wfA3WJEo9PwH5lMInjFRDmu3sRUqrKx7ZHwwHvZF7DOnrdEOdv5/M2t3kwcwVtB15ok1p6YCAJuW
2ab0g/1y/pYxICJViuuBdPXEvMYY3XxWo9jJFk/cpoZWeYSWkoEGWf7e0TsU1i3+760arbA/98EK
xoxrjdMXvJrumG/YPwJK3AhpOqAr2PBJDxd4O/rmFL32LV57TvbMhykJxpIbVYKl9m3ktMhu8dl9
Vr7sXe50co8H4oBp3V2Jd9LYFdk8gT6Wi0kxLu9w8DxZtZ5hlPDuO3WJ11U54FD9Oo2aiFr/tXB1
ZZUPIP3vsNP8MvoR+9KPN3BIWlDWba21ISHGa5uOBMB+LcGoy4BqFFrOQsC4WadWJmVQqv/J/TYJ
4b+NQyc05nWdHBJCOtH+qFjalV7hPiH8yilMGU5duPG1sYGLQGncleK8ftUTjlUPA5WL13mQO1mk
lwAtziRHPqtkPqvKZP4RRbwPanLRzOsGsnc8yjP85+/ntT3R4fbbjxSuYaTlp+7+RoR60YSnmHUh
/JzDx6JMpefNd4bPKE8vowgxPd53zmsBBVFYS27MfeYrdnyF+NFLaOH1Z0gfVPsUGVKMvp0VAJRs
lfmyP/rNb3yn4LXJTPG4NEGdX4F6g2lJsC6WpGlvwo5Z3Ti+kIhcoxC6Ufe+avQXheC5AMAMQjjJ
Lqa+Wk2Xceq2hMqTbpO1kEDSKFtmfj2dXgZT17ngXKe5VLNhdDqnXyEUYglmfGUcOLPCt+dJl+NB
XgcInwDrjyRQg0eIdT+m8sH1jzWJMXJSul4jSEz6IhaUa3RftxsE+9QP16Y2tzPdJhdso+yM/E1c
Kq5tu2T8+FohDLqnD6AnLVK1ukbPkdJNIhvoTEr7TaHj/UqnXjmuGf46TASJFNdaYvfbkzP8qgEq
KhOqKzEbPYOynG8hLxIyVW6ecni4o9SgeIglaoDXAo+yJrMyaJhgbGDrrbRUfxIrkj0yqUMNPy/M
vWx6kWlYBfsU/v9H9v1ZMZ+dr5MlGLaG3DNOqzMcI1vnzQ+xd+sqgLCkA++ybMrSLHYw08H4FxJf
b7o8m6by7ftnHBhR/oDuZwQMMqBO0RKuFrMInSe9stWL6svM8jF8Kjb9Ioc6MYeHdR4Fjh6rBVBG
0TnPRn+CRfKiUb2bg5nE0CPnsQVQFv+T5tfn6dmAgAq3tHbu5c+Z4G4zoXbE8leGKWsaFMHiLHMz
7hOm1dESRoCMI801FmY42IUlSoWDosFycQJMRjXvaQLpL2TWjnRNHXO5vU2G/MOEzgS2LC6quJYU
9PnMwzYEevUtXd8x8eZRpQIgfRnye/Q76nb0clDhSeIcQWQBja58yvbFjL7aWf0xNO4BqW4iPJgg
xtMT00RdLa/xFCapD5GekYb6IlMowUKf4NzZ1JN8k+5hAJpgibrIHbCcD1QqzuOu/e276YO+vuvf
CknDPtMhfGexKro3mKNt2JJ1FZEYC2TmXUfvGbN5Si+EB4SrhMz9J1EwhK+1JQQwzrJlSRceuuGs
9ZNpzYE45xiz6VFZtTqc0jSL+MiaDE1Oq53b5PfaUtSSHNaOwiRl7/THi+LAazgMp471YoK1Qx3Y
PnfS8k0i7/b69pf4W76xfJC4ZXIMrNONx4NFPsTRfiVVT09eR8iJfjCPdDQjkGGspKfkfbE6ThcO
d4/H7OAwaXM3wqbEYVcPrkIO5NeTIETK/1MW4kmUuR5dpgnyOT4ddh4efDJhkzeVY5QWHPjAFMq9
BO0BnlShx775K6W9sCI9B3SkaYrQXPjxNKVfNDsVlAQkTiHaMLW6KFAfAV1WAtNdiZtnzT4zzTKw
f/vc5T7f/eQeL4ygr7YMhOurR12NOJJtxLefZIer9g62UKL8zv3dZ/OhyZsp2sSaI+W1gwQ0DYMo
gGSJT1oYrF/0+grxnYTcv1h2aVkBuIDUjPB9H9XmlzHlCayhNo4AgkrH8CP7q0ziD0Kk2VhjpfzI
d2Sw6K0z73ui70A2+SerGkfk2yB/vQHOPXZmFSuwXZdVNch7Uycev1Pl0Xd0kXa/SG8l6jXUhTaF
jn0zbvpCbahcFNORlDtjVWrGGWyA0S562DKzOrK7w2rPcp5AV1ZF7oXPBlvgtDY2C8szkI6ZdokS
QE9W5G52DE5LRlv1PLGVfEU1nCnkO25x+zYvdlMrUJK99/Y4dy+Huwd5vELVcxrlywzxdDEo9xq5
loJiHsqgdu3Gr5UK/GHCHalQ6TGTDxAHTZ/AZhlftMNf5HXyvRDq+c42hdy6eJRv1KhtftThE17B
HT/BVF97WThlY779zLS6EkonvrWChpbeyVMCwa9cJlLJmEcPWrU8un23Nx7H37XVgHS3wdd6YZvh
X8Z0YaskE0DVvX233h3h4siXB0fNnnioQp49RrHU6FCHEHbcYo8AvwN2xMneiuK622Pa2kAz3owi
X9jDQqHY2nrq3RpAyAqryIJN8zkfIy3wHUUL9Ay4JOwQxLYY82JLy27GRmusynD+DCd4W4w4mSgC
SlRSBjfgp+fwcXZ9qhZzgcgduHDuapsT/gC1RNznCqQAZMjCGAPJ+rHg2Q5UXhejx4aMO94Kj3qf
xdhVJZLMT1/5CgEGtK1A16D6yQZ7cQFTOvxt8MQD/q9Z+vkRBfVePlvhcnkto7QFXuS78k/EPMHO
3Bn8BHEbyW5b8dPg+Ncdepi8ISzNbXwGOLI4p8NTOZd13WEK7LBSnX7Q23q6uZWvhBcL97p2tj8o
A7j6DKWJAFydkjJgUhp+bGYuK3AGM5eZ2GuhoChZAVpJfNGuek1Mx8+wJFVXGxuntwEo53A+OrYR
3faqtMFUbuYhm8DNpJTHphK43RhhI5CbH7z/v8y5pn25nP/ZqR9sseBGOXOgvsaw6xpaKeD5A1Y3
qu+O26mE1MRSTL+Z5SutMCEQLEzybH3aK+jatnxcbK6whjIu6fqR9gZPBhLoWn7h0lWk4My1CiSN
oDglCvDOxBeJS6wsxs8PjwbepEX0bcqmPpdjJpU7XGJOD4ZWDVJPtv+RgEg8+ADjhBKw3qNwNwnR
FydWKiD78QF8JpzXgZr4LaKbB96xAcstoS4bRhO76O7e8iBrcMVjSATS0Pe6/QOyWfYd21/c9Q9X
x7TYtiYUOYgUgHIUeto+x9LXZZFwUZUMHeQv72i4r+Qsq6SNb+S2YbcFedzlEsCvfLJu1yZIzX9j
u5AMHUJMJcZ43/tz5I0YJeedrFW/38IV/vk/bydLLNO2/BTzRJ/niQn4EyLDWM5fVWgpwJWRTEnU
/w+7PI4COLToG17OKJ1e8/pH3wSe4toAOL9P+JCNbNoHmCeFD9PIGjcXJMUa9fJ7zH5DGnqhMjNs
Qtn96Ce32z49Mgt2MG+nQz9wHkvvEVzfEVKZKUlTE9xoAKbqn1zfBE1pM9NbwHYjLeyTyw2atkpf
0ciHWqAXFXSP6xkExVon3+/OSBi99RqyL7pX4uCNmRpR+kkjDoAQxN+jOcLLi1QklY+f2mn8TTm9
8NjaBVoKPIvg30NOkGZ7JGRHOoYXqf8LateVvfUO/oDIfpBGo5JQesUp3bIgjU69+JNx1OMnea5S
AOdK6eAPr5xHAtk0MNI6C8t00GA+LL3FgK70APzP/NO6Q8b4SNiRXVH7Fn+HRY+TbpD0i+igc61a
VuAZ1MGMpIGlPrxvltNDEuRpxurkZUtsrK+TpNSC1C1Q/Xuv4RC6YIEs38zcqfn1DN759eaXuXRf
FYf/Y2YOaFIZguLLzSGRr2wSrB+c/7zo+N6HDJ3yETQpnoAuLsdS80H2oD7KWs4p2MEYHjXotEEu
TVH0P1i/FXnUuLSx567oplGprSIpyfdtABTwij1TLDtdvmETWBuFMz4Co1fBKXoVG4MbWP9XnVvh
N+TdkIpRFf1bnP+PMihSJJQpo3hVppKhWGwe2OeQRPGcRK4j1KFIUkFxuofXtjyudNHsi6fUo7+O
PfUAgzNWAf4GWr3KjnHY+PI7mGefKqQhaCU2q9L3Ot/Q/HIJ8+VbTOQPU33M35ItdXc5Y7E+mD43
DEA0T7zyrsKnySete2RrTqxd6TTxE6MN6K8/zRpnRePCTBw6mP0PC0yotcgtYKHnFy50fadKL/ze
Cu8kuXKA/js8xUEnu3wWUv6vc9g5zTo9idYLTSdnuKzs/0R7kXkk4kSUA9FiFwXI0mevz9SFkGne
oLEMPLRxlT6MvqJFNpsudfIjL1KTCXCCNCYjregy8HPVjSuSTz9Ag/A+j0QRTI9RHyuo8WQgOiEp
LnDvgzA+jhkTnWP4wChWQ2TuKOgi0Wh7NpLSjuR4gmBCf7sIgcfFjABa9Ox6EV2Kzbe9qz3D3JU3
dfasmpjve2L3WuIdrKaOp/+BhKmNkNOg18mT8GUFTf/Wr9PpGgy2AJukVontvu2rsieLBmS4UCpf
cCqNM89MguK9mEfc9REO5EN9qTJwmu7lnLI/GnwRn9A4Qoe//iwDBisAsswgac5H5+iVGjQbPuek
/QL+x/26is+34LzLcPmUhIrUOEwFeOj745iNcCL36uIJSiFuuu2pjHqmj02ouSqKyQxgUzUIFSEA
uiKjOe+aUWX5MTVO43T6qW8jGVQXRg6+vlxHfQpTfqYmC+M2178w+0ohiNUVPELAgagMF8frQPg5
i+yuEUZm2SM077nVmdlfYA/YdQVjogrjS2QGCa3ZqRVyt7NbMkv8s+cwGO2JzL56KWB/QVPLM/l0
8LN2qDFQy+sAfe3pCNTGi3JOQ5IeyZW2iaREWj+5HupHf9JhRpY5VzY7K0Up6PqcdUBazUoq0A1N
AYMlGknnf8w44A3IvZvLJqbdguizu5JB2A5gzxNvtJwA/InL/WY7T+qHpub3wNxSix4MzItHzoY9
wKcNLxrRJDAb9lgn/Dk4uaOjaqaM9Bwik7waYno8HJ+/uWRWJ/ZxkLztxnk7CnP9WDjm4y1YjCUw
0RgZzKCCn1zzdGH3HsLvZpUybFbOUxHVGCSvl/rK5LamHi1MwnUfyU3ld/QeJl1+7TIXjgMvyrsO
+5715M9Wa/CAo7hg/i6bPGumowb562jOimwPVty91jfTW6njl2F39/SrUmj01acQUdHSEAN+3IRe
YL6DCHyxXRPg+K99nKU0EGPgQSvS3TzKUwVe64+kxCDPG8DF4mRqRU5osMFAVzV9mtQexqn5ExnD
RTsm3igkKRbgNM3YqCkucOQpKHidEG/h3Kd+XFJk6CYDpsVaVBwvL2PbdgqKRxqmdfeI4GI0v8X+
O/Fztmuk0MkLMBu2CutnIuJmO+PR50sjVypFwnPIPIuqPiEhli1a/MS1Fshbc+s0upkdXZizhRhL
SLSAn2ZMQAICAr+MyZ6cMRgLjGRdDxIVcDjswePYiLmLb+LwNzG1TitSutKhr6+YC9SXug0o8/m1
iL0bY2k0nkcQWWYrFEyARlfgFWdXYziGCU9uz46RQYye7K7U5tQXzlWc7xKg0XqaypQ4DhWnfTGQ
b7d20Vsi1E+QEZucbj/GdcYfokuxd5Gn+50BKp5mqjMGAwmTph5ob7T0sz5MJmEDbwY1ne6Oj2pN
7TGSxu6zZzIcOIZPfoWwlvUdoeoaEwJ+EpfsGoJIsM/DxJPAd4YwEmDO3LR+LuE/d779sfuBct+R
1njNVxRhNL/7tedESi1kt3e3UNFOPOuynMYCz8lIJFLOHIlG23rMRDzlp1Z4HhjjyapjkRJdw0WY
LU75x/5CtVsrRnccOFDXU4d/YNIpunxjFc6UYjkwBFhfIpJ9zDiKv30lya4TM5RNJntgvIc0w5Ii
aPEuG4DMJyxvApB63nD0vs7o7a/S0IOdtpARE2RRpB0NmUfYUWguJ75TEKBnR2b6OlMa0RJ8Ed0b
hidFDzIpC8A0SsKNTyHa1SSxxOz+h5A8eYwgznk5z3qWRJTX5/Zpdw34BWBS5j7rcplMLbqRjc8O
CGCnXlqiXNdB/1V9XqjFH3VqNh+sv6mSkE5X2U2s/G5Ett753/VgPy5gNBFqpT0NqU79hye2lNhT
e6X0yLk64FZFRmiKwnzku9wLLoKnFx2O8KKFA+axmcSP8uMqHhI9/TwB/qt2Qjh9VI7htIbM1uok
Uxh7palHBupvSdv2V8jv73dsOm31DUJCOnxC/NDsznPjMACGehTiXzSH1iuPn48aoETN4f0i6P1f
HHEKfVa8vRkcx4NIv99oZ1Xyh8q/2rteWd9YIhFZ+BVvL3PFuX9sjjMrsBGPrSxmmpPWlNnE6cM3
U+smGlO/bYFJKt9yZDrEcOh0jqNbd54ei9qoD7i133qPG5tJFXjjwHkUbBXEiptc16WVSWSGgUm0
Q9fu+WtaATce42PIvKOhsjYkAD2diPKkIbubEJPVrpJhkIt4Zsyj917Zos1KmrGIgz5JCmXKqfMx
UfqFxj++s4kLZTDyelafyOwntbAZvFmZ2QVP5BLuasHUW7QZznfhvyK1J4fbBupFeznChE9oww2s
gdQLK+KK0rmZiud25klHPiMz2TX1cu9gmgugtuPquGKlmnOSRZspj9g4sfTTM6LKKRE5/z1aVqbi
UCfMZwm0LCPr5g4GN+F2y7fYkuzmXVqMBBSFjEuZWllvD1dezZM7SrLvjSnNThtWs71RZ7Lpva1K
3aQPVp6LiF5b40Dbsy/3zM0gW4MSY3AlLQxMFBcsEHyIPO8FPYsJPYcrEGch3G9g1fguR44JEh19
Yw0534A7qE5aDOJC3QCHVKfO1orrDPL4R0lTqqeaQm1wz8M/91ALUdW8dQYJE34rmAAFnBJPw+lA
f1hG4PdauahZxGDbMy5xpn+cosQkyFezyaXKv0wdPZYANt+DaUAlUHmHYHkGQh97iwFdwgxNyvtT
n/Y3RsGmWdXNAQVRFY+UI8mdLk8y21j+mWhjqghMrb+xcLvW1dRouGoLsBHSVMouKkrxAHzAdgJk
k7kfeP3IrgiGV23ryG46CaId8LiyhcNqqer9+tP6moiQm0VDIY8xzN/Uqtj7smyLrJ06PO7EAucP
t1RPdYLmFkmU4BM3JLg97FZLhPSEkdIbUNMbSNfV2dws7CtgCAhmwQ8v6ZDRSoHdhkQPQ1yTBlEy
c1H5WlJlQI1i8DTrnq76TaMvkQEKQAWk/8WKo5bATwqOw1gRZxZbSO4buIEczZK1YcDOkrGRRf2h
secCeWTIeek5Pp1FA9jjf2Ck1LPXL9f1YzC90KDMUrYoBeC+NhY8i1iLzWhVl4kMZ+bUs8y3bRRV
XG09w4pNoY/20MV5d8BtH5igSvbL19YWcl4+cIz2APcqGedfIHX1gEbFxW+a4LgUANcRSFEClFZw
qXKrulSHsXRM5kKHr/zlBgZwAdD9EFi2It/r95AY9ZXpjubw05GBgy9jUq22FPSfWIKNznv81U+1
nyq9Jeu6ZY0imjMJx5H5Dqbr/vZvCCxC9pTYkRQxQ/RWIyUtge0kKwD+2q9yAn26ZpuxUi2DC/J5
k0JiXgPRPC4w5YVVaNnaNj/0uEqU9yYXl7kj+A9mfeG4cxy9B7YM71f+hZkK0MKZg8DUJwtB7W9p
lGWynud13aOSGY6/BdvUWudjeGtKp7fl6asFXnejmd/Yd2I423xuk9jl6cheOBlmozojdU3C6i63
oJbxC4pTt2Va8yx7+H/7am7U7D7ft3uAnNRtUfNrjzm8Y9KQ1Pq4+Vc2OQLLhEVqvN0XJc5J05m9
4+vGpAVkE3nEJLvQl+BC6Bn3nn+J1xkifk1D2U7U8T6894KAxEm0kG5GUMFn4v+AhewDelifvnGF
fxf3Ai3b3WQHhkKWTuwG5pS4zp8i+JuqlDbqlv4rdFqI3LVNM1q8z02+6+RFPJXqltqQ3rYC1WWs
yNEJ663KNnRG7KC9S/s291ZEJdKkL32PZNEfZj8RRMdA1x+VylQtiuyI7i9+L+hbXNa0Ftoa0kAA
t8M3s/m1EeqY+CEkLqzfVyshe41s46VGZhqEYMLkKrdWZwNgGjhg8SVWkIabKZXBJIchxwdV7PiI
W5EscGEC8MTDiXtpRFX8jAlecvLWPw4c7+lo/ny+lGEc4lDm6XBQMlc8CkDbTi1YYfla4e6hTQmR
Npf7hB4Eh0w9DCpWcJ3LszaKrn7IF4gqrUNpaKeDjsLIX50hBRBHlf0mxDo7LVZ9x2X8sp+M6evQ
n4Me71StUUFIW55AwpKf/ABgMgm/gBd9R+PfgeNd4JuuJOm3Z3GBdIsVRYVF9tJ0BYB36/x98dVp
cHbAVquR5jffzjP+V03mSCEA9HY446RRCdO47ehS1/Tmtx287w9dWb9Lwd/yFYckho/+epX7IEB6
/91ne1Scbgphek11u1Dbx6U4VZAAKnn/yeZcSic/jDXjhgBPiwdfNvmGi6QNauOk53FNJ67Ka6Ku
VAZzUwDPcKyytcKQE6MQ1+vgx+VtZdjIfqrZufRrshuBFikdFDsq7o31TA11QjeT2naaOpGlHL+4
tfcd0hobzrpJxZO+kPcV2OKrCIWZlFBRDXX/mJCkSQKNWaBLzP6Y0h++QFIh3PKAS3yOE1HfNik+
p0o117yza2CPrbc2dBQtwUWwrRTWDPznVf5TkiSBaYeTnyRzPelcFeeW4IMSvOAit8rUgLI5egwV
BpLpP4fGmFQhmoHA1zzErHptl+gvk9qjOnJb2fOavFiDXIo/jjNuk3KVtffV1Z+BUoY8a+YoNjQZ
lkuBIXmJWKsnB7drJiOVvT4aWMYahHjGCRUuyFmB4PcJ8HcJwlH1s1N25enTCfI4Q1+5Az0YYjuG
YVG1LisLGrLyeM7IsCXnhp25fiK6MlsZnBi3NkrR1Snd/3ILuhrKpgVSAHVXOj6zZD1CiTyNb/Mq
5o/KXbpvMOZ6Hczgy1lNQgdowU6YI7JR098rCJJSt/sWNkZ4ypbQrnd9QaveQ5CSikrKMJp6sYds
BF1j0p7ufk3GqXcVM8nmfkncX1jM3GwTssuLFvzLovXOpdsMDFsZgMQvw58vTC6i0wtStM5CfYSa
FSAMfWo/xWE1m6vu4NNz6xGPi3wp1v8tuqyKOJRcaZXkBg2DzTddR8eOr93RJhwOlKR5g/1YvKIf
gz9Lpr8df9EyJJRKhiIUeIyjD2z9brsxdwJfU/7/NufFT8W0Zc7+HEMxufoutzbylkleghjIWId7
3N6c7CWAArIuFCvFzFV5ZThhhUUpWV0LWMxDvFDbnySJ3hpZhW0tzS9DdFLlqmsQ4dG0HzCh4gjS
ThFQUWmqNmw9XcUT413dxzOihrT9zIHLSAJxQa9bJtalH5UqGDZS00omzuAR4cMSm/dv6M9Yt2eo
kvmeflNnIt/0kXh/fjTlSbEjUlkxfvynxK69uDLMDXitLxp4AYHu6PIANpsMnC/T6zor4KnX2kN/
rFs8T0hpk+uFMGfX9Y4xdAb2uoS7tMVh0vB8tzBM3fToF/ggORrce4QSxqT2dd6DI91Ijnm2CAyE
z7HJQj/vTtcdYVKJ1EAwzFh5ZfZlBaLSJsWYkZw/HqQzef6V5AMISUsO/7fsvzTzODb12L7xSwbo
4yrev/dmyOpT9f8zm9Q5h6y4kBRlhFLLKejYMn40eEGvMsacNDqBVKK1R5ACT9LLNzAbFyym58Xd
OgdvHl5b7WZ5KJ/i7Vht9mNfXF4xVrFqyGCD5ex2xBoXenYvwQSIEATLM0+E2bcZMXjmzqXs46r4
xvkxQOjD9/3lFD1mWeQlD4qkxOWuxVu50pdH/ht3KVhkH6Dop03ON1rGY9vPOB3W6HUda8YgVqGm
cHR2cc1gyZujMTQjqkPNxObv8zo7I75A458GGayne3E85Jrn1sfQHlT1VJKoCY8jgTGIKEpMOiFM
sRpDk4zhfwZdwj20OaOASnb7UJB/e4p6EcXadec4S/N7IJLrFcbFcGqoFhjwA68bOROSev030OZY
s0baYJIUE83nD9+9iI1ScF4wRy1RFnh2E4Fx8apaC5De54xIgK2RxFT6PUYk76p6lnJfxfr3W3ff
nqbgzEAzochi9BimedfcIFM0LHQ6TG5Mt6iRuFiRqdlm3VRPgHEOyHS/zX4qHURBxwU4z4cGijNS
hDkmj1mR64XNNwhQQXwftg95kUfSNcVHIQ+trUkyv//1MaAWn6T7yACLKOPk6Hp9UKOUsBb1mDLA
PdnskzwqBsBgvpOC5aPQWtswp8ulHok4+jMvfvx5ZW1wngcSWRL6g9OdCt4IRgR+yd9UBmqy+G3J
CxAKoi7llRvKm2UR/RIQYBZKcD2vFGyAzIyrhK56gOt3sj51QGqYZ+svrKHyBRv5lrLT+Zl6H3y4
Gma1Xt7bekHNryjOcppVRFjZbDtNcF7L0y6Be+MEI6DfPsIqBM+2ZZkZGXG4lVTMWXySBXhd/NSQ
ldNiZYdof2yqyogIm7ZwBCKEaQ6INajCeVVgDWnVoIom8oxVYTQJ466BhMOm53ILOLXy8EQlJ7MW
fka86T9c/dtUogqSoz1rqKHTDc2djX7C3RyB8YpYvP4geol3ZMx58hcWzwwWtU0AyetUfjPp5sMF
KxoLl2M1OWnTrQ069l0MqHabAwwskgUjxfWUNbOa5jy0C76bfFPYLaKOmotHblnETopww+bfKfCj
9Nf8TtqFZ+OVcfYRbwzcC1KpRQOcdAQGEbREX1WeRKj/rR939+bMnOY9fLf5X/kd1OYDrb3yB5wN
zKMubG8ZALb034CB39zpIhzTZVQK4qpA1y+bEYcgM84ix1TdOJL2+ToP5Yf6G3s+QIzu0QmvOPj5
4pKTW7q5/rniRKSnPgWPLlAwq+IcWqJnFF96D4DV+5o6Bpb4XBLHJxutE7v7SH3o/I2wA54S7+Zy
/SPo8B+4C0eAznJD4wstyQtB1BhijCa6S3rngaBkxGud6p3km2pxs0SLl681VkF1RTZmS6J1mfjc
N4AeSDiqfyIm8ZUd82iuF+a9Hr8WOQpDWjUTgNk/pYBwaG0fuNEVshTXhOg/7QHmy7g2ti+qiWMb
VwMD/y8N+UKZmM6+UBOcJ7+VL8xbv3wyoJVXgwPW6XxtwwCQexbvwoSm4gADJBN3ISCdjdpX2LUO
fYo8ZMZdQBJiF/RXczEnL0sMGZsefkK7tuqm+ansWTPHFLfy2OYOv2e1hw/UkVqWVmAZtQRym5MK
r66IpBxgTDckMxlhNXE/2uqA7jsOozsYHgeVd+6EbN9gi/1et+irycFc8FXzek+Y/JcCdZ49/zak
NsDT0qK/QlYg2WjzG5isJjoWEHYsDXMyqenEYX0a8OHlX936UVJyQ55otuf3QkhRj5HMjbHGK5rM
+K5CQhhW/8QR4rbSZPbSKUWYvY0YoqHalyWmtZ29dSoSLJsfs/2olei9DHgkaQbSOcY2XUcGRcoj
w+q0r0U8+phvdxShv0hZix0kr6S0PipGoxhsNTljKcWCJix8OXwmYEEAjnFyXRyc4Vnk1LZrF9/j
138Ks3aCUFTak1uh6KKxPgVb8HucOPy2EXF/7mW8SSRptYBw0kp8l+8ACDnD0A1Pu05usL26jWMo
KVnLraFPEnghuCixkSdXMW5ISHuvTnxCGPS/Im6LCLd8QLmtCn1oIt9bUnKlNHQZV2pNuFeQ7J2x
WYCMoBAcx68HOw5HYb270y35NmayUT8Xjq9t3Eb2HihLXKPwBxPfkcZ/sWaI8lVSGebBWl2oXSpV
G8rj6sWCV/M8c22iB7HxQH5wPB2YWBLzvYg+LXzkmEk3w+9DUjTiaJyOkze4LtST47YtpikLJB6f
wPRNgHYMDVRn1NS9mZOfQMEW7InDEZCCYa3Z97O5rRAbQDiwPSBmO+iD6PfCW0Z3Zj4eFvgDumH9
/e74WO8ervNprrHPijJ9memB8ldIvxH83rCtMptbQfHzEgFyxPnG7J2nsRUwpsIYg84O0OwUefXQ
6bj++Rhc6eytq0uJn4/mX6vQvUJEY+LzdIj3qE8wMYkZfZGqDYkXmYfbzv3zfHkVCWyT6+lVQ7a1
qdUNZVoNrygUHFsn5DCqW8xpmgzrGLKhDJkkv9T3fprxVz1uvFFVneIAnOS+qYMD29CvQmOVElky
MI0yNx8KgWTeWkeTp7RU6Wtc5t1RG4Q4kO+1/MaFVH7v4FrhiPC+TxcAUGzBfKZT2FFby5Pg8ySJ
FQb/mHdH4/Er7ivLNq/t5AAKRs74wAJDoqhqWlidX2KtALY8Bonpc2sybWFjCtRk+3gWWf3ffg1A
oZ+U8gaYlfH7pWFSOuksCmTF3BLHSVBrQR3u+nSrwnn0Gb2+uPg/yrpl+eoDxOjKakStzqCKXtyB
aQjBtK0zPNWTiedXW4fXmLpt9F30gILfacm4iXo1zHbIF1q8LEqJMj6zEN+afO1XM3MgpXP+KLxi
WjzTQettSG40ST2RIj13iiOsE9mQ5cVOMJVSuNkpcN0Ba8UwYuX+YFpQtWeEbAWtA5RFSEpv/phQ
0laLmBTdNzguS7TrjFhaqRvlFw2W8mAG9XD2hMoseLBoQHfanjImpo6am9WCwzRJ4V631PEAD4mC
FyiA4utaFZAhQ8GKz55zLRgYtK9sLkfJpP3xlXX6O0ihsCITqQ5jSCMq3X3KS/cldSBFK4BV5q/j
YLzEPNNoW4KjnszFETxb6DAmzuCqqMcTT0RBpJZyBW6jCy1DzhkNb/IlV3qK6AeWgS3aS+/xT5Jw
ZpWOoSGBz2WROvox8uEivJtb/f5UfbiwiMqJSpv2UJ41CS5/nCAsOJ17XZ4NC4Xr8J+OVQqQgb1v
a1p0IPcP5u4Ai3zGdgBDTiLZgaLocJFffBUwFjOCPJ5+eadwORvWb2cV35ULKKZmEwbXGDE1eUeb
tdsZ9Oed0Os4wx1LX2ON8sDGthcqZhKlOLJUZP0nixQYizeDoTHVHnOBA3s5KLJK8LZm4eL0dQje
KQ0SYgmIMYgPM/TjPqWeln+2lO5pmtHMB6rtkPQTvpwpQC8hav8e1Gh8A/UmLvwD9WcEzkJpO0wM
lQRGLIf7JPD3p31MvLXvQUiq/XKwYHskiK7Annbo9WVkuyvQ3tZxKIRjnZonEGrGWMeTeFQPNqcq
oSpmA+ejaXv72CkCavwB5h7E5yCb3+746zcuTQY4rZTFwUyeJnPZDp8P4gDCtsgfAS+4CWVBmcb8
UG8dcIudBGwYD3KGjS/HkAX/Kw7oJZ/OeeVJ+kPbMMDuAE9FapLDUIprvWRm3ybeZKUfYZw3onJP
IFcD/2r4K1iZHUi2nl8fZ7qWnv0xaAROqU2P/Vwb/0Pv8j4pUpf/eOj68OUqNgNLRTrjtAxmbd18
jvWLlsaSk1XzWo5U2iszMaJ8NPnXeGE4FDMaRX3ToMFjXEsUfPJwWTql4qgi6eH+KLzNMPUOks5+
fvmITHhSSbnGZvtsjfglh3vyIsWzW9urneOIW6S2Ro3Miro7olJe32B7UthKSJwFqPP71OGdbkJk
HWwtHL1YMz/ucKIefHOWXTIdqTUpec0Bz/zSLCjhcaKHO6f2iAgAhnxoCM7GiT7qgB44BJOGPkXt
OehH7sWAs8+lptG8K3j/HTvuLr1tMZHPqKUJAvWqsMqd5mmmUDphTaSxxEf6nqIzGIpoNV1GumbL
S2MwURPo3kGg2f1hiijHQUjm42jr9imP0DoJuKzGPrVyBEsASEE3HRuAAWGP7J8i9+PucBw/ye2r
ocr1E+CvAOHFsV5sizFlfdsDL2NykNdkRtyqVMg1Eqi+w6qtlwAZx9I/0Kq/7fPFATsWhhCq9wKT
MHTPaNqhrQO184Fh5oN9evF0TIY8ypZpgoKon9y2btY5jrrrWt0JFZsT/ODwbF5rNVHy7M90gG5y
c9G7lIiOSmLt7XJKDtkwIF2Cy4A21fHK5yfFERB6gbGEwXVV/o4Oq4Ou52iDNH2i143bGMTXKxjg
aD8sMI8mb5HDkFvNn6iNPHta3GuOTNcHvQprPTs6w8bn7I+qxhfsPrwOKVxTrtwBWulmcnIDVK6z
KNRjVHwpqeygWBIg1OdPoSGZ8mY218b/jWaL0vOEKP291VKocg3XMK/t2rTKavngWwfloVOYrW6h
GLuc8PdIEq4DQFI9XtIm+t1He9llEC7N/DUGGvJt28d+LB8OucwHdGHznaH8um4eBGnPwm5b1Lvo
uNXGvN8rrgobVHIiTJDsNG1/+JMM8MEXuxAZWj9+zDCaO3xHBp9eSHtuKjxyeid6kX8KQECHnuZN
pdyipszcYkvGzooynrKIdo4A7LZSxEKXrj4vU6LoDFrM2QGzIYnUP/T+DKy4YZX0sFw6+c4Wk4wx
d1EhCE9NsVdR8ZxTgu90GItKnxx4mhh5F28bwc4rB0zBFSoBhP/jGfqbfFy4GKL7AxfnjtNyJPVT
dY3GpWgmVVPaz4Ih70LzpaAC/XPLa4hGGD0wZQxP7gVqETBTJwxpKBjyTuJnCh94ImW/Nn0Ua1O3
iNPVlsltwOjgPZZRxOic64HYKraIX1eZ0s2rweHc7Dj1O1dhRweKYICujrtKdxGQDDEbeGHVafhc
+tMgmHjso8due9X99UHkiAoPawjNNsqCQkZxs1RkY3xVCgfOfJku717daPfa9L+T3ebQ8HkzT6us
bxkIFBlCUjG12xJwVwMauuaf1pcdy78+x82uNmFl83D5vomPzjwXrpVCpn7cdju6KfNKhQPR7TNv
B9Qz+M1l9mSjOfbtyJmuclXqRJFUjzwkLqSxdv5WRdRDaVV0YDJjW2hps8urBE+kJqZmNZZwrP9B
0VVLzlyY7gKJr0DQ963au+2f714QtyPhK5flHIoxhn1jtap/mMV4arKiRvgoE6yUTo2C7aMHWq6c
zNtpVCtnKQiPVdQ6ldX+YvH3qdwh8hiPia7XjuJjvLgHV4Werzg0mpge9sWH3kD/6dktJpfjK7At
gwk91kzX6P8nB/o+UM1M5MZ+IHCO+SjMfHpwFywMoNoDdp9WTLfdcIVvWyOMWJaoN0S38Uf3sKld
uSCbN/1rDgyLh/nFxuehegJKHaDEUM/0toleuVU3w/JQ4BPGIGIvq6Hry1JdZTpavJmYoy42yFoG
cRv+R5vl+mm99rNUSYOGO1YchQh28KFvMfLB2mYlPDbRYwm/vP2gxGyYNEaY2IT5/begApdcyTHP
FJKc2pHQbbj7uXqQmU6XsUcW71shIbUfbcmQTDG6+7kfxHw1yCule9j6uOkQbNlxE5ZigONaTQBb
vRbWLmaSTChUL6Bk1ywER3BlscZ0YODPXmMwNYw62RniMZpQ1xHtbblds2gz7UtqVUa7aTtKL5t5
t9B1/DmKGR5E+7oglWJpZKdTllEn/vm2SF1WrCFzmWI4PL5v3PJb22b9PdduazwuhX4LDdZm4dTd
/7eiLako6Q9cNF6q4WUaDQ+qRqUxQrLMiHCboaVyVGDUWZTfu+tSYJTBt3waw2sVjwniTLErdUpx
q5Mbe33e+h7Sggbz5JkZT8nttqq2EqDk1Qa/r148+3dSeDb6RG1mp9Z4PCizwggCIAC1oJG69V/B
vE3U2CpujDIr1Ie4dqMUDEEhSHlxWFar9miQZogRXD6zFVWKPlfcJjkDTrtiTeq1h56z7ZTban8r
Z4AG7ru80SdDsGhbgHKa7ycd0AufcXOnxq3vsoxUbmB/huYI9tBg151biQIpacF7uhI9rmLgK6q9
m2ISgImsYyTm65ol45oCasQ1vmPDz/fAdnSgYgmygPo8n7cCCkwnrqVXfuDd0pIPQyiyN7FcB/2A
5PLzr+YD8KREGdR+JmPHLj94UHV5Y96f9WuMviMkofxseTdt24TFYTJozu9h172LCBXNY5oy0252
xtMKG9hUHGXF9rMq8Ykq5JgXy3KlKj08hejAf6EaU6Pkxsm35dF8xX7KJoZuOCfvgGLwTmOc1mVO
8rKRRgwGk0EuNK9H+PgyRqvVn4kWNrFrPHipGbhd1gStjIWXucqBN5+5rs9AbvO4J3u+cVGY+q8S
6z6hkDmYJtF6fZXMUE7kmXLCptJw1ZO3iCsdsLs9ipTQn79/+1jX20p0YjH6NbQwHqM9zE0R1E/F
EilT5Bb8cHdNVhInGYlJ3ArNBznBoIQkn08LkVs4H3Vp2DVULQWIEcK6S3Hrq+dDtT3u/HsEgreQ
NM24yVbAs+cFjzIBmL6it0GaRgfNblma1YDkLwWePC8MqcYFqLK8BvA9SQps36jwyYm+bXNwGX6z
E2nFZ4ivuVcTsaDj8wfR4XIe4oB15qZHUVhKhLUfCFNC+NPWKCCii3xi2sdjq5iHWtmvWTQ1OWKu
TuzQ+B0M9O+jhtcPvCOMvGCA2IX1+iOpW9ktqRlR+7cbWLK8vPeoakfc0nwetMS8aVrQuiWWGR81
bMvojWfBPVfrsufNTv5WYcF2BbxTEY/QrmfxhFwrVeBb9mGEsALmbmPCs8KP5AzA3j4hDFP07D/q
HVA6gp9bR9QPQJfX1PPu/3PXsH8LWVfz1G1y1Q44qvs9zt+0ghdb9KS8fSrvhqlxtK+aiym54WFz
LCxG57MOK40WnsDsokafNVVV+spksBoQjybePCwETJWmy8Kwacc36GHx4U06dx53eY1vyJb9AwW3
kcu3cIVYaVxatl4QKqKEHJDa6o0pd1fpJK+0ZUzyY+lPCmRf2Fmsczkp8v4Z+nyMTHzh/jxUeNib
HVlVUkj4SJ/N0g3y2NkEvc8y3K75WcWOtcGWqacy+T+ZhHnFxMhJF3dFxfbI/zRW28tIhusR7NES
/h/cYerHWdWxW7ZlHLp1+U9F3ojdLFkLIc5fttl58FifZiUlU4i8xsvi6VirkK/ySoB3GYMxKWbg
3HhocIzdPw9Abi2g0jWeqb5DkvwBlSEGjwLEJ/s7HPeAhR82O8izsjPcfNhg2Y+TnAfqQrV/2P+Q
s+Swg4LRPC7f0bACKtJ0d0sNL4Hn5tnNlQnqQA+xd1O9PStxuNcoichr7flamaRlSbScJ+Y72S3T
fxTXQVY7PyF5gBHy6Zobf7p7uvKFKhKexQJkm0ZSh8Xf28QOHE2AOdzx0RxXjlB4lckkNL93V6hf
qMzjXM6UgFvQJyhwVtNqayr2TJOCMXhgUpNObXYkjLeNdOP84RRKKlBJ44VAwfzSTsi2oXUL5aNk
09ifVMNMxV5xqiz9fixQtfXCKVlukWvaQSedSWza3ppAXRMn3DgIIjUFffY9aYVmr6qMe4fOZ32P
7+rAEfYVHtoz8dsEGDhdw9PpnyDOEDTtImxM6rRs0VYhVGfOqrpQ8CbzSk8xa6XJwLUCBA/nT7Gc
wR56tCQqTKUWUWFKBxw82PQ523riLH8NJrHPtNf6+XVwwWpMMyzoa367sl5W9frj7lwNQz+Ru080
cwC9qvr/m2saCM+/QRfp0fTZ1ItEHrmBR2sFY4Z7+HQKel7fWe4LQSShEKiwpPNN8lwZZX1NBTtI
he8UdfFKcUgXAaljXqNFaXsTWYVBwdikwaizV9phZWuF7FTj/7d7tFzcR9EiQg53VaxM/d0cJ11z
uEVxP9ISuecvqLOEKdgLtT1lY3QPsSwJehE+rqYe9ZFfh2iTQhir3YDcC1KIBhrX/fFi4f3Bl3qq
xoyRyfkVpmxkFUmquHMVh26KWxZmgFS4pdNSHF9hIH8L4ikp117jNbOS6oolABVDmVoaIVaSgX+c
tK9Byq5TwFkhr3MklCpTV11mLwqbRhe/POlC86DC6EoUzENwJSf2mndAMU6APYt/UQsGONEyP4EG
/GgzxnmjFGOb2ltdVonKNTeTWTWDQcYR94wovpCzXC2gD4sZdJ8UccjafKodFDfc4OMaONi7jW2e
V+yhBLKpup2h2HbzwnLEEuyXs3n2uKSdnItkNtrBxvHAWbcNm6skIetzH96U3tSAMbeZdjRQHKg4
TIxvAjqzdSP1ht3HCjIS38k2zLg3/Y7A70/+JDzOj9aB4QvrjF9bpIijyjIBvfM1ARZ8SUsAuJKa
XZGvKF5lvJGWxLRvjo/9ZW2keE1nvgav8YHYepLg1Q4PfmQ80LcG48SeuttC0eLXQk1T7d3OQZ5N
KlYT/mrWvKuOuLaiQkcJDj7WyLg9YRpmerhnumDBvxrvIU6CelYI8sOeARKf8g5pc9g/UVl7v1VL
u/cI0jk3V0/4SQ+4Cuse0mgCUVIs5Gv8rWH/sBXSHIhBDD328bOC+FKmYZ8i9Am0rYiH5Vbno0e1
DRNUve515sR2zJZ318zMgttJnWbyWaICaEjR6yxuvNMZfPE81jKva77OjErARY+e7W+Q7P9/m1GK
EXvk2w3TSu92BuFQ1wz9+v7elNZxB2QDT3/RvJk65FBEh8CaLsS9obFO1XzVgLtG4EH0syuANahI
aSjcQ+6d521lByaIadDDBp4W3OuMNlOc+XGM5Ew6xOK/O38YAUhW0jnpTBjPoPUMcTDJI5CJ7uHz
vs8CG+uDJe/wY3DboDpLugAfvvpG4eRIUG/qEsz2tQmRM0ZLjpSqqI0XRSXjQii030xJgmxrbJo6
K2QsSnuqvbgtno6YZ+4N87bT7rXX9ddZpMa+3ZOWgNJv1aHh2zBB8sYmjB83XHWjD7k91dYeDxpG
mle9sp00QkY5vqmZpjn3VYGZNd6gWQ/szCpKCfaIzeN1lG8yu5+grMx5eilWEl7dq+HoBQxzeYNV
hmNcdBPabAqJnxsGyf8z+L4OPu7oiB+TZieXpxbFOl8ToKiuytvyDdXr7JBASTSy+D8C+zPWW/24
/uYiemWX0Y801OulvRIur+lzVO1bVZ4xQcMmSqoVvwMBofvr4Ro/UfzYXNN2lvl/+MdhDgYqBfEh
7JjxdOsriFl6AKxx1p3M97F7NQOaRBE4fVUPJUaVQSKtNHdS8vidNcwKKdj8tzCG4aDBPK0B3Qxm
ZlGhnUI3ZhltyhmWP/5EQf5UvvBHQ1ATsqnxpOrQdr9YFABPRS16cK7iFcb/IqI3or8O3dr+T7vz
2XVlz4xvppkQMufJA4hc/9tO6v+ZCu90fPVOs+hht+YMM+hpuR/IY6L7mboByu0kzP7ma6oGjaYV
ouAS22VVScwYf9jeRRVv+nvzeFQZWqb3cj3/a3yH1qnIhsMH282XwsU6UoXm3ym2FSgiQcKHzuT5
B+hYxf7IlRpEZ0wsEZHcgNYjL/QSqm0z3mqhul5+VIDyCibSISEtDUQbWiPP6nDQvg1/IYRaOXy1
otwOnHhsBjbVrVh9vp4rG+9O5MlYjDOW5PK3KXwejHYKsxcDUgVoW9DrPDC37DvidPQHCOuNv4CS
GzYSuGdikyyliC5iZ365ZHs6a49pvsKkBa7/2ck6w3jAlIM5xIGOfLR/GwNhuvozFne8x49sOMRb
D4MORyYn2Xo3B1dlykBqmSFc3oBe78/S/aCanfJYgmHhubUKtSKGbAN/MJ5IPRVndAYutF+9OgF5
OBfEt6sVzLwDBe3efxee+qi4dYZg0aHw/4Cih8lAZBs5ksVx/gYx1kSHggPda+wG0LFtZb3MDVza
fh1KL2qb+Ig/PamuRaZ1DPrx1/HAGZhLnOS3lL0C4QsL+AzS+2c+TuzqEl+eKdXBJqCL+ZqmF0E9
oHZjitJ0l41NJtBLQ1Sg+Ru0/OGflEJsZ1rRKsY/9ZSiYj489bOIyVd7NqMnfUF07U61Kiq6WbFF
X5eJnAO6q14YssJcYylOG5rFRthPfGP/f/CSlqCiZqwwHk6AXZ5phFscl10WFqTzExTIIBw+RDpO
2qc48X1jpOSQS1JUNpmDzEBgKEL1Jcy5szn2B6PtkdLvi//b8bjOiTPExNG/rDy2E2Ep4PD0lfd7
giTzbw4JhPQjXgPY5FhIK6fFbfGchSSOyiL9Y6iH1YS7oDaOtvtKffYJkj0/qNBdBAZ5GLKbETHI
8psNqiSBGYZCps5eB/fefTbdgiUnCBO45BdZqa0i4GUISMweBVUvvZWfK5ehIEnBgtYo2M7jsXFs
LixVUH5c59QQAB3vet67sYNpX+kd887S1L0hPuLYhwq0dbFQ8kTmvJX2M1J5zMhRWc1ZsUEz/gGG
5/qNapbL7PkULx3zLSwodjqzvzTC9ZC3MLvCf4noXs18ZKGRDXSwOtwDdSr7TGa8uVOwkggZb3Cd
JNys3XmRqWrViz1uycqEp1cYK35q5fVy52TAZpCaRS/g+9+8T32wQYde8GeUQyPGOO1jfm2KciTP
oTO7oOTKjm+ber+JAImoF9CHFFqEZPbQ7YiGKgGTa1h6B5uwZztVh/NvrBb5/fYfOU3t21sxkO8p
n9sMgMTih1XVV27jtOXr7oQH5eDkM434J5lwpbpNtg7jIeneIx4edWb5cCH+TDc6EAmPqCIvJzVL
6EZmUcl2+6BF3kYMUFuWbtphLxsV0xdvEZ2AYWF/GjGdirUc/Vx/NZof8RFO/dt06HUPPsToVXXp
yBw6wfH4Y3vpvliCBmMs+UmFW4HPd75jB+E/TDVyicRgGma3Rj8UfAUD45ru+KxJioTsDzt8xA+s
dnlxZgwDk2kuE1cmn0gdjXOvsVSQKt+u0cpZJtAwhXmqaqnTF4NKQfALXsxGbtzdb8XzQH4bVslr
89rhOrK9Vk2lJtrfF8tIjKvIBRnNlDR4B7bfyp5n8hIMgqI8jZsFpJMBLoxuCv6hENSIey2kwEED
erQSZVCrb2kA6F79AYzLyr3WOMLVT0oD2oNNRUKpmBNF37R5uJW80P9J+A+282cqfcEaNdZmcqId
evvkRz5eTL5g0pEJKuBglvyldRfBRZqX6I5JD0sXfWZQpH/TypEAwUVuCxMTkQsRVG7vYrumLo7B
/pxAyi+PKPXxVYrOq0DCtU+QQK2lHJXGjR5x23dJAJYDkx6qOKZOLzREOuLVga4peFm1CuCiOslZ
2Kwr4NuSbzH2xyaN8HhvVQmnDUIsU5Zk3c8XSWLvg5IqI6PdH4FqWpxmpC287BGBpTjBmAfK40sE
8JeuyDAJwdwdKAqSpy6X4LMA6PiTbw9gh3iw2sJEZobByUkvE1FOOoAbjU2kuepRe+vHJYbkkgiO
JgHXhymZ0faVcZEibOyoX8FflAhrPGg4bZIbz0iwEwhQwAviI3AoWDL6K6L2lRP5SSYxoZs2nNZH
vXuqnm8f5zCC1qRtj0PYua3IuvXFznj/VDlLlPgu8NxpE3a1kh2ZooCOaeUbXUNNyyj2yJuXJrnY
2rhRJknH/r1WSl/PQKYggOYkSPQuokY9NOwCji15JApE9BhzpEqUeCAEMUwgW4y+h72FPRf1DeZ3
6uIBEx3jCxBNZo/gSK4orcwKSjF4iaPdm7eapBx5AsYAZ2mV0mftZ5jP23bYZKjwO2EwBQGagei3
UR+QI4pZ6CQODZL7nby1Egi/+EsKnzYZpCgGqaqaw1/nOiTof2b0ny03SmWVx9aPOZ9ih0yC7894
G+irVK8KmvuY44sgCzd87dhEia8mJsQS0PIRxVtb12mXkWunetkX7BwEWE7pX9p7QFgj39/nTtmE
6r2UR0hl0MmxPO0ZxYQwttTXR9lV/7kcrv8HpRNFIAlWl6KwOYhomFnbZ6DUY/+HNQp+xcWx14mH
aIHaJdQIskvLKeSKkSKooQ+s3Z7ydkfYNM9nuKnckzneKoIoby/KYlMx6HoQbZWb2idG+OZCL6UQ
qxXX7Qz4/UPQrQiCZV+I3G+rO0ORYsAZ6zBNO6ciI1UJRCtFHSk4cCiil6JsMNz+xZzck+FXjq10
AYLDdlOiUGIVMyaCRuEW/eSNilrdu1DiDj7SvZZKlue39bR+nDA0SmUpiwzHYxFWSpurNG/bGhf6
1Of/MLfEQP3X5brkbo29rX9M4TVkt2eaAHBDmmbYvqYdtkFux3BBA3552hTqpsasvn5+xkIBHJ0C
ec7tJX+pURwIF0l0O45dY4gecxxgQAVxu6o6MqFksXopaQwfzOGFTu3+GUvZC1Zgjgj0/JJST+J5
0qFsopFhSuNLHZY33L/aAm9pV9fu+oQ31rot/UnSSL7Rih5vK42Zfl8nsIDIbSP+8MRJ8AMeptwb
2AZqgiRKD5UW+mtrboLa8Livppx6US35LwM1Dn/DAQjKxr1kKvX005r9MbKd6IdEaoiHY/J1HcFA
aGZFI0XxYKdaHlDTYOXPDh/B1+6JXvIYzyPTKYWAKmsxsZ2pzD9k931ctb89n1I2RYJNU4TQvdFG
C9RHKtZLn5B2wvtZq4XtkRhBcVqRNtcUYQOZ95ot1HZ+UJD47y9MPlODThTOjMkvDLk2yNjxPOx2
F/SXNQtIpgTh4YUkaGygJ9Z16zvlZCqrrBpRal/z0NBrSt67qhm1Pcu9UfA8ayg9GUnAXUZusXt3
+sLkUee8BEPW41+ma4DKFb+GU9KXJ9NnWR7lPy9IJ/Bbns9TLBsa1C02gp4KFDU1SZEgZxuuDc9M
6sKsCbc74rPYaegG0xRTVkoeDEiYFaBrsLXIwWdij9u0J/pnyWzWfIXiXsWJ/2rqQdoeXJdbfuUe
Q6Rm1NLUAUukwvuF9/PifuFxTWgGuc7VJEGazyfZ4c/Wpa6E/UWXA7e9ZHRl0y+YFrW5H2/Ep3ko
1xHP4Ni0Arb1Ys/w7KaVvjrz4oN+2gj4ocpch/Lcsctb3E5b3HATvkikc5+mi3WPDQVSULh4Oxfw
10HE30Cb6ZhbzmpWvZDBDtqaE+9Qul/5ND5SpZQxLVtr7vJxX6OJR4XVPuh7e3kNHLHOyFRPdoe+
Byeee0n/PNofSIpGeUwGmw/jkKmRVfEAYPe5wSFm/daeFS12cFe0PzJKuN/LhYI9uBX/pQASuAP9
/6PtbQ6liY+s7NGFv5GJKyS91rU2jNWeAP2FR8xWnblkksarCwkdGDgMVjwg4b2ginv1ggcTwBkJ
gq0Ko6Ej/J/Jw7PMqu7rL+0iCpRHcz/vFmjcO1OnLPZIHYZe9llNzdMpMwE5xwqdB78QWIJ7a+iW
vcR4RaaxgkwerS4mKaIP3hU7W4W0sgELT9HhMq6/8wbOJ8aH6G+vZpERoLknEqwjxInu7Nc9YJjg
a1c/jXYhBCohT8sgZT5Ao3q5hMbxSeDGfauonVW1PQ9j3H4qjDjpw7q24qtJT2f7nTL2y+3TsAUc
t9GrELK1AObxjh6/KvXaSYgblGMnm1lJ4pXtpEq7oRP6H26JB+KOlGFMK4OMIoMBVjHyLECiCRuk
+U0he5/cjsXaeiEPGNOxUf64+A1233aVV26Y0QYnDZ9kEJYKX+wnGfwJMruJdV1VBHDPAoZvqCwd
wbXsxRm0Y5Mlfc0dk9QEyoOK76WohqvEIZpN/pWsP76qytrNq4MeAbu/oEZz/p2v4Z/9tP2qHiER
v6pOPywAvpt33PjbeNA8/n+3TJk+fwo2lKiNcZwIuXZrkJf5Yu1Vk1MIKZSffv8b4lHtZv1v8oIH
x5eHyCa9N6AbkM8ERxbmevodEvqFepKrVSZXNDRQq20qAeyEkXU7HyHtmDABGq1KZweqfISVcJnU
FoAwSKi9uEgPG+n5kGy/u/eS8PS/Q0yFsgW3iguhj3AOuD2SKk85HQCw26s3G5AgdOaWKagV+iZU
AXlp+1eeSGZMIpKlSJhQCc+v92h575KljTSnt3g2Z/wYY6CzH9g+iWmQB9OfiV73o8byz8cjGIhY
4LShnvAwywZMzw2/e4Hs7Y1adEnqnp2DVJedc3Jm3e6liSmxoNdrC4FzaDJ44sb/0uXqYeBX4lFV
47/BKSZRifZatyilJeBX9x93kdk9WorQcENlTfZCftYgvM1UCdb7Oh1nGi4kMtg8sFGitQ3yTsEJ
6w5gndjsO5fhsMpm/iZvSBLC6wCdhTnQrKTCdhDwJzh8TsW4vvj2iv7dsuCaXbxP5+OC3mLtWpqj
5ls1gJCc2qOjVBL4Tugxde3FNu1hDicM7TxEtyijmX8nB367Bv8RLBO56Yfi69MbeHdjvq2PGDEI
ofs6sxoiuTFMTz6nr6+aXG/voepzr/9sHpEtoT/9GXpxSTVheANWz/0NvY+oFhMMXd5PX+GHYVXH
GCez/PdRv8NoO3bW9tbNgG+2UCyKwxHP7V35GmKYcoI/+vCtknq9HIuSUNJWoFn5WzWivMEWBD3I
SxPk/tgeQuxUmtmjf+k3D072UUg+8faTBjSNON0nv1k0tJtWthrgc12T6wvef8PMG9D79GcOZCEL
ofA4FMoyXNpbcrTzN9WFWkdsz+juE2QcHRyF7bosbCn4rSJOo7upWZKSzOuuh4oQHeZQiCI1u8wM
v96GLytwSrsY4z9auvKkLSgeWYli7HXiDeTbUjB9+X9RMS0GdTIP6UFkWGrF+zFAVzlxv0thzUMo
8EPEAdzUVdneu88FTnefNyQujt1vwNuPK9RNatQiYcq1BsLWlCDi08SzxoJE/ARs4bFu0fFwHjCb
xN7+oHzxjJ0JTa94A3FfJb2VTREFVf3iXZU+0lapUAWaEqi0j0bLIa9vq8X2AWwdX17/LaycUcoY
5g9RXs3izb+pEU3UKF3bbk6D82hyeY6zPybLTHICcNmaiajeuE4aK0EIeWA4PYO138RLSPSXrcjY
NXbnljCA3SfxquIaJUXxdfWLxxYU1BDIbNEtC48ZZJ6NSxAGK99bwnLrm4yXazQ77Mm6wmRmTm4Z
bvLfyEaHGMnJCQU6l9ZEfOIiW3iFnZ4lSpHCqryPxpduXsCZL38UVXzxTdccRSCs4DWwR+5/OCYM
kQDNc2jvATqqCXnjvvBvVyqqQfZvui3HpV2owoJS+A8mlKOcpHnVSuKF8tGHZkHUqQ8jyzc712QJ
kCMxnFA9EMOdQBAyZcukg+duhjczHHN3BNOgr6Wke0dHF+qNQq57HZS2Oep5tMJI7RNTCehhzcet
q2SgeR7J+eFEcqXwEf72qK//+6OpUYeDjBcZbod0Vh2Uwk+/oLAsiK9QUQvZ/M/uLCF/lzU5qO5T
X0456jGOgOn7OQzX6i3Kgkq07wntdeErdAcWqBzdzQDOmKWqLn++xiDpzJBFH98so/chGZBJr2yN
rvxrnlt+qF+ymaQ7snGlZ1L6/fUM2E/GG1LJpdEL4ecTgig5KUfmSXqTYsIpLBjW/kjZvRWmAftF
on205l7QjSTVBWSOp3o6CYj2lpTvuRZzVYa4zzwZkVnGfqniEWfnnGHmLgI01JUDR6yAhzGMxBtr
4CxcsmcnEOHG1A4J8+kJD7C446w7Kk8WYCuvv6IavsrYqyTiCbzPPwffYHo92DTyJqM8/fDT4Whu
6/jbmwruynpuqfu3zuzEKL2VQ1vLLIxTr3qiaGYWNj3wr3U68a8lQ7w3EKX9nzsguCx6qxUIB1v0
sGuuNdLbTr35JiB0SLCGdqVVqs9Xm8A8EA4aJwuKxyfElKDBK0iWf4BwmxdTINTxH6EqiU8/v3VI
bowrLjX0JoBKepwj+T3iiaaWRNkHFWqfxNFEzfP130UhWpb/fbYuC5tUk1KBMHieCYvq98o9Xnbt
NjwZWpIEPNowshKU1SFZe4cYzvbxvjAtd5aU9+OmeBaudMktk/4GakmKQk53bX/7f0TH7/p5Kh2K
40Tn0nY81RAIC9kaZ7q+6vn5EdDysC1ctKnCZ3OgGA5VkV2RVzfIoUHSc+SbkSEO+JTS35adJ04R
7krkjv8QaHMBWzWTCGQSQML6BkVT11Sax+RcTXbidYR0UPgvkiLz/BqkgZa50AheN2agRzBGVr2P
hOUeUG6b66AFBp9EUujNFvDy4oIhUwqv6iRhVV+3kPNJOn/cTV7weMRvSEXSY/S5C7AjmDc5iQvt
9BGDiuhnwHld+ul8EXERHceMs6EkSuft0eUXSv5KoLUdYtvQzsyUQVPvGV4kuHEvJMLCO8WGyE+q
44/C2w3TGPxgeEZM31mn6emyg7kRQyCojg2du7cV8oKkjJsoNdz5k+TYeia7++6ZAYfxYRRM2uCy
JLKHpDwfUjky/d57iWI/3mcay1LFvZ000vWuOhWroXjwXq0sXgHkcF+K49OA1d7ps07tIE3bCwzu
F+qihLEoMeGnECWANVRquyiY6jmYIvohV9KzGOOtNVx3GW0ZouKSKNoFj9rnD1D4i8smH63LESjL
d4ngDNdf444IeiMcACFEwAnkUiIWy5JbPUcRZ4M2sD0nwkLbnpZAgPOaOieC6uMhKuY8iSle5Nit
krOGCxONl5pGW7941/iujQeFYKu2r/2bsDNM2VsG/KzobmV5I05+LJDoRwSXiz1xoUBj1zkaddsm
6EapgdE3w7owjCiVfrpYbVXyF7k1GJg+MsrZn2usM/Bra99GXSlUVKeW4t59SZcCQ0p0Bln9DukG
XuH5QUyCYu/NgnhwyRPY7WlMHluED4Qb3NTg8fHB4V1U4KKN0+9KJu7sHy8E78ihXos3IkKNgX6x
0mni6I+8iXd95a19LV0Feetot1nKS1OeBr4puQUnOb5B015k2Ry0Z12/HBMtDmNlRCZjzTDI3T24
7JGTHQIx9VEdWEHfOFdhWxxxTwZ8V6h7/yiR43dLOFaevsXtUgiJ7Te4pYpoTe/xuueIkvR4AuuE
+wfDdYWa+8EkeU+gOwYkacTVc99ccDhqZtb/ohJIFfx/z064mfBgK5YupwsKrvPZehO59QkKcjgm
kAEdVs8V6fYx1hRrN4papzaa0HS658I+XSVIJtd3GYJNPRN2XgkdLfxh9uU4l4GYGFGyuJow1Snn
WAYiEKKdyE4JrdNJSEHevKii1GWyGNYP3eYx5WOi5WE3RTggSQN9eX1N1SLrvYFhRKqwS38J3XI7
huqginy6s7KI9emDDlbmC4h17oiYFhNj65WeyBm7PPL9u8hv/tMW6+VBC8p1mqXEfG+XBgEjQ9ZK
SnSazDAhhlgmVIlfWQFnq5d6FuO6CwBY9TDakDpbVGEI+jHwoCF+gE7CuAVLxJH/2Mmz+pnWHTBs
XpG0jaKHBJEYwZJg34wiuGDi+M6evpJhQloyNAsK8aMpVF6S4zobbOGuAU+Ntj3yNzDDugy2W5I8
XcE3eRecxTDdoRtp/rJVxWwQ6srpHJUdC76ud33TY2gDavDSLAqCXbty/RxPAdyVXmtxQhV/cODq
4OCxXSjV3ZXVAecoUBE9l7Trap2Wa27C0l+DjA3iuuQG/Oxs+xza+IONTrieJxwu5zvnpAzg0AdI
l4JM7htoNM8K722wK90ucrFx6sZ7E6EG741MvanVpkxb4GNveDYACzXHOaMAe/wUOEdAW0nfj6B0
DOMEF6wGE8oiFsstAE1kxtk4qcQS4wB4CW5xgWl39ze/pojCd7Rm0so3ZjZ0fvaO1ASyGK+A52cv
oxuPPSOLj5TGcu9nywgYoRVWB/hXMHouM/JjzvJTZOmM/lnWMm1OUnzlsbYpJff2OxBNoxbtBEiD
oCq1u0235yn0rRbMkjG4oOtqqzBJGCI/1wa2vRQGa98KlwN+D3ZNdYFqESdMWpElN6fHr/ExeH4K
VUP3VpfCUnD0+QnVBtNbnie4YeE1IChNz50Xu1+z08vJ+A7ByKVqR79g7sxcUUVWQWnntoUm6Hj4
MDV5dHWcusA4bL4FkrDPfPMbBfy82KlLaniis9CJZU4dAW7NYux+P+JqEU/wVHK9KX6rEFhX9ZIG
ZW5ndUmMeOOekPn+vh1g1caZe4MrI8FYTj15dfJmmJgDo4sz+YCb/0Uqnp+toPujj0nbkwke/D3w
RAb/FEzx+1G6HjTRTVIBXrF8egbo5/a2CgpL/P1Dz2PhvBgso9l5fhhJzMHBJcGAk1t20HPMghWG
iHRpzFWpR4zC0M5PP8exvp1RI3m8IyEBtTl4q8dJSDgZgiNWIO2dYPjjqWgGmki9orv8vPRXLVDL
3piDipc0TAVCjg+4GupmA+bECLbMOzKbcYk/r3Q6cMokh60Xo9KOrbCs1tf1K4nLi7bHxJf+uD85
uoI9pIhGrhamb43gRughAfEqiCatG1TtKE/6eXGoM2hsyDi9l6Lb2smLvfMK8zEW8GOPs4WCEQs2
GAqiqY8utqiwljU3fwnRWQ88EaDdKUp1Y0Z6P4sxr8bDzZf7TLaEllj+5NoUJ8Op0yifu2wGu+sk
NvDnh3CgA7RiievGUpvHGAYzhnGlAsRqEjYd5PQ6iVCOaZmG2/01lqqNT2x+WTIRz8jhLBTwZPoP
1tjhClat6YnJN8Z0B9Ep5KN799iqVdEiEPje5Rt+tx/Ff9N//gMl0Z9Qy/gWpoA9WePMA62nV7D3
e8Ul3WRDbdbxG5CwSHDNkiTXrc+jprzRooWDzWuMienSoB4cBWlkcUvX7XtvXLrRjYvnSo/HqQb7
dL/4Dvf5uCmRQAvYFCld1PD91Nci+GMokWeWfZZ/YvtevvjFMwVPBKgMdBotobjon751becCVYou
skRFMj2/5fjIK32bNQj6hiWuws8Itx85PtBGpcntTUI3WTG0SzQH6+uqMsfTTIWsBakMP2wfScfj
3KqtmOjhBgFfB+EjWUtfqGIhetD0gHNGxy9u2vynRIKiFhv6AAcEw/bHM2jitAs56cSRznw9CucZ
mdAjRflV+L+RBaN9yU9TX79jyQ6I4a+oYkvi/M6SPgf25/A29ng0qNNTEH1QVTJNtHFbL1Dbiowd
n5M6l65uRYLP4oY7ure7UMsHIcnOFHfkK4p6ejMf3VZ2KgM2cAkqk+wOiRB7DDpqYHd2tXUTt0ZG
YZ+FDU22Bf3KYGJu0CzVD6EWaN55x8xb84qYvdXjZ0uhBZWopI6SmMH0ddsbs4sRSfa2c9Tpa3P4
gMVRFklp7aLYcBNDgxLgTF30PcFgBwylaqumaR5iA0292LfimsmbkfieetIFplrGBtZLKXfJZPq0
oUgxLwXH4a+1WPFcQ+Vb9hWOoz3i7gRuKGKYe5jKhwgRZ1FYlt0HtLJ9VwoE/2huBwE2kWgf2dWt
etmXT1efg+6m1Gg/aeX/lkVqF8lZFWhhV1Nw2dCXl9HMEYyiNjC/I/eH0l1/VxkwRL2ieJdnJROv
SfC0MDt3ydNKMZK0vCIk4sIieYDYjUVINfTqj8dTyey0Vf5Tw7Mq+cIcAC6OdRSTEoz5QUOdxkKX
g6i67lTW/umqgyyKYx1Knla3cllzFoa/dz2Dpnpa9dgEmg24XFcrw3htRc+CDUv7PSRM2/4eoDVY
JSaKuCDLcwIXCUsG0SPeBtKV+nIPp8sMDS2anGkaV44VwPr24DoLvYjrWLrK0AmR908PeRu1fcpe
sKPDgJixAxt0WRCAvG4CEo2tLzwjDdvgYb+h+JQCI782s4DrgUqFUH4LXGbhWTu6B69E4y8OhDDr
bx9dPEP/Xqw2OX2STCRCRtUOol5ThwN74kPCSpBWyQc6O0/eLFlC9x4WzMhRF6b9Eug0NC/Uoi0f
A61FsLBidT73lPSNnCSfXh6RgnfppBId4kWlNhX13C6YhZ/Gnu6DXbJ+GO9YHXsHuoC9KRW252dw
ltTx9iWgy/TtxfKfk4CCPOK8gwJ8D/gcpZsgyLx3XTU66fToBdxHHD9dkANoUz/sgtE5JZ6L9oPF
CJCPC5WF1byZA1cCLlV7zJ7f0Zy8mcfA8J4KlEWI8FpM6Ta1PdnK2zAdtChL0+MsjUhLF/BhJnSJ
7LIr+C3yAu5vUhEbu0wqzfq5T+aErlB9b3Tl1vj0wiBbx5SKBfR5CwLIGVHG+lfAbYnqxSkaYIpk
VJbIc4Rkm1YrrTWyY4AVzVIYKf4I50cK2Ikj6PS8x9Qk73lkRpW+O3IFjXX0jzgmZ4rRIFYtUfWt
9hs5xUHnCinuyzYmRmunNKU8kYOOqRLmb/Fo69VRjopcuUmS0myzfFeCKSC/I2tLSQiAGM+LrIWK
Mb4EIufCvJmc7JiAPyECjdFATl/nEJUOuUzCYEPle72MG1T91/Kc2OnMs3XVPrRzR+eLxmGsjrfN
KO7Tzz0JrXrDzyVkUzhDrOFfLqmC0sPxH/alsoE1xgeYHD09euxPD0nrxTtcHGGzjB+CoG9jxtf+
zQ0KHX1361P9dGWdi8U9B5n1sn12r0gZTzN9e1/2XpwCBkwNPwNvWy6cylbMWBgbAy3cRPfR3CXL
mnEBe7r5T//nyN5jNrmFBFNLOA3Q9UD01g/XtoOJra49MybokqEBM9eZcXFe3z37EtRw3xdZ/ryZ
EgHjCdkYGDzRBzVjMWvuKHcs5qNbAH02Nf0UyywtJ3gB5k55PS3VmqtjusAMvmuE8ZizovqqWCC1
P8fIzxQGjpwCmMFEdqtOBVz1JiQ0sAdCw1HEn6mdAwnVhm/7+MXbL4DcY6bPasWDSqM8tbAtYuvQ
mMj2okrTrcryq1xjgomSCQUWpA7wIHaR+ccTq/C2+rgrk17xqhDYK8Jy8F2iyMR05wRWZ690ZDaj
P7qPjXZk45kZEAMaZaTSvSUJKFIovwISabf7pgG1lTTWUXj8Vp6G4MjOPMeSQuWO6di6o3znYoqf
417lZs9PQB/WeEc1O4kNZK8ASfXzfjXcNz8TgsFBYAY2C1KrZnH6XXfjFNJb/Tn7GJlsqpC39Blw
dU2AgzkdBsE3tCQHLQscj8GVJ4M7MyAfio+Oikjmi+ex27V12OAKaDl008jBPgEIkCF45yEsr+rq
JXtTbLLQyOIJs9S8q9/JUMd1hblcyCNyKfdmYjUrYtbKnLwqmqDpCkwTT+8WBtmmZanneqrsF+VT
DzAyVyffIfMTaZQ9fZ76kZGmPauMR7PUQ56yYSr3LiNW3HSNDnKMw9ZtE7ZrG4ppQPmnRtzk749X
t36Boyeu3XoU+0DKfkqki4YhTECSuDNBHQpgYQ60o1mkqM+2KBHK2PtyxUM+a3GLowSxTNDZEyF7
t7qAdpseJTs0Bc9CEDB9NpY+R3HYOuYNNxdf+b9Bftl1T9dViZnpUXSMKaYrRjNNb3eMgQGcmlVx
auEeq+guhuOIWBun8aqZWxApS+CO0L//wmHNHY0F0zcsBgaVbvpaDbWGzqJ1eax8ozrxHZXgXldH
gqtOWYZb8YP2a7puXNx6lRswB5otQB+Al+VCS2UVF/PZOTezsBjQJVvbnUvELL0wqbt4DshtDIWj
q/AnaL2T7Ao9TMfy9Edx8qSvKYVHROPAVz7AL2AQft6uZfz4GDOVSdm3YobYhFGJ2JXJKL28Yye2
IV0OCLoXCfn5dNFjB5exm1PGnjdOtQm4W9wEY27OCJ29FYbtgf76OfAJ3K90ivHpaeck+v3GSJZu
dfMFCd2asH5J0fWTQoNltvMRUuu4t7N7TMo/dtW6q2lou1p5zcvof7fJ/YJ1VqPhNajk1RzY+oZT
XMdP6A9EWq2UjqtTuyqkleYcWrOXQVABFmVRer7wvUKsb0/mRFI0wVSCLzxuMY4UX+7/jRU2eqen
EU1GG8QLaOpxEcxYC28pBB0ZdM+erhj5pTkzQKLxEHERR8IFAUqM2SWMI+nDUO1Lgb3VmGByqW56
dLkc1lHPZschyJr1dbeZ+1wlzKPtN+svB4dpc1bK5nS4n20X1Ko1YB7uLic4pXDjEgi3MZsQv7+R
Www8TKMfJpZaPmFJoKqP91BO4C/AsCEnn2Hyty0Zaeb6nKcpmRQNf1nO49jd/MBxlhzuVAAa24XZ
mXUWe5BplAOXlv5eR6ztoWckmjXEiZeCfnUF3mH2ikYuGp5VuEwxXgnP8khTCAJkcVLuDkYSYVi5
VthT8mhSN4vWdLCHba9XmPMh/vRmrE5cA15KU0Q9y50FvBWaiDSl0Px2ihEu1SuDeTy6UNCRpCv6
1I6Kwj75fQEY6MxEj1prIvJp4C6bqYpzpdOKf6MIzPT/5giGOb81vpmAIFXOIufTuaZFwMvY+MZs
V1+dIrgrk+S2x7QmhEFJLa141r34DDAw5kbrxHark72nrBUY/mTaKRcHgeviS0SxCd42Sd8Av0b5
Y6sFuAOZGxkwrSy2SVXTmgKUWVZXaqLcVmGzvGabgd7uD18cdmgGcAocYW+rlivGWes5QFYAh+Qw
+HHkjhrzldSusrhrZpc6k71VpoofPXEWmBywhVTp3Bgh8Vrj3HjsMrCGyzZC1oALXSCQfXda3EQ0
EE5LtpbhPzCKfkWfd7FsA8sCsD6fPrp7pEL5W2GEeIEEG0b0IXdz73itjRkLHnGvtY683W0wcbmr
VImJoD3g2Qn/SrOB9zaIEJvYetz/DRNvrKpIA4tnP8fXhPFrzsdg6khkCPzQbjkiAPp5ABHjnhzw
yDx4B2hkP/RltyQ9WXOsFrGH6w8eseREaDVmmeB60JBwKPT+uEyUWJQ9gnDeZL3cUlUwEndwdQAM
4H2cZPJBPfwQ9IbkEhYRVH1gITiaYg0FqkGTthDnx0KuXyMyc04q2a8dSZRJuoop3XuczTjkNu7R
RbkbGK9NmzrPhuNkUr0WIxl9ka7K/FfzJaYkoZzQk+y34BiFLyo357e7B1BFO/HTGhO+NoSXZSYX
wM+PLXfCLmvDuZZnj8s1egESzFIgQ/X0fJtG5otNvCSv5OjPnx/4pNWxMxADItf32l4qvJzbNTXB
wmbo4xnijrob/NLGQH0QT2FAhLNzu4ZUdOEKyOuJ5HkjukUFQ1ej5O7qesL8emvaTXukqjLHbuvJ
It4sUyBWZd2wKTaQgzBDg/SA/UIZRi7g7VrCI6ueaJnanCwPdDApU4SWUew5UYEP0vbnRgRXeG/u
fvj4WR1kx3gMEOuf8kp0fZ++fOw0PGzYSQOPyEsptspl3Nb3XpmQZDijtdZzwV6LoTyRpBnF+rHz
PFO7wGc5/JZOJIkdzBKVp/fZklT27po1+dgFGJD8g9vwEG49qKTrrxKchDu7lo0QeYqAiv7IzhjD
m7w6iqBUD0RMKAimGmbbW/kntiSGTKgtMJ2stXIBKNX9Aa/FrZomedwQdnuXI0tReAHfJypvU5N6
51nezHaEPzgtHNJOMEfJfzBPRrkXq4bKh5KUvmj4jcLqdPRr07w9rSejVc6d/v+unI7h45n+b/2r
z2RFCFrdqb2ISa/8ooqP7CDhnePU69iFaNOywBaEv0GLPO1dlQZM6y46tC0d3Jc5C25tD1spCzJ4
LkibhdvKk0fH3huNgPSY5r2zBhDGiXi7ttLasvaXHetEfWAJFvjONMlOmc6wgPINxVx9/j9BnTuU
7C5gerhRtH5V/v5fsSBLyBeueDuT5RS2JVP3qXyeAM5MZqqUNPG2fFW3V9d+GeW/eeOnBaTs7e0N
RJNf8eN3WI4USCVmVxtSFvFfmX6lfl2wvV1fdLfwWJ2lK4vo0qk1YGjK2uo8hUV2qN6pPhG723JF
qpfmSm7dlR906YQuQa/keMEl9VV26CLN5ngw1WdTNwbV78hrxmhvW3GHEBWocKPfT5U06vvSxNTL
B9CKsCLhiiFFs3WJ5DDiO7QMRPXJ5mcdxRuzk58eRfRLW/QVqKM3ZVBzWATFNn89Yi68MNF5z9V0
1gEY8YEofc2j3kMiOhxp6ppmhQJtzHdjSaLjNF+LxX+AJRzf+F554KpZti2Lk4nNu8gqgVprB1Ju
M3Yoa/uodVkA03Dezcz36OhGMPnQ5uABRzUc76v1LTFF6cWFU9C2wn60UZMbAOexdf2W58ipecAG
HXROhmYO/ibIIGjko6+Y7nQgc4xZKSA5zEgzOD6cX62VNIrM4kjPUekgTDV9UkxvRU7udKlZLGsW
j8Zustv7oI0eBE+zB9jIYkHYRYduaSZmnkyOyKmB9zx+EgO1WVwwhRc+bWDnzBiGu6/hr9CUuCwy
/d0qVl+q3BWrNbp3C0zTvUm5oo8D1Tiw1ZTYJW2lXxK+SbumH4SY/LIOs0qliWMRYLaVYw9l71HK
swfxam6M77PL6xqT1ZM3sZQac8xznoWmE5Al6NWOvdNhzJpih+mKMsTyJhNZJ+Uw1IQe2yOVtyll
yJwShO/ewLW1KjRbZGPtwj1EkpW3cjoaSE0pIPmbVaGV80jmzqxsfKRglAOZk2wYcsr5f3OP57Zy
QErBXZcY7V0ypn88ddzbpQT/Z7PJE9zh/91qI7liUNOf32pZQ59MYGuO+qUKjIqj7mV6s46z6t8H
jU8tZ7rLx9wQB0kQloKTQo7CMD3Jss9WJdog8uw7DF/XNRV8id1GQSMrFUpoM6D77fczlOa6vNfJ
e9xB49yTIsWhD0coSmDudRzApxv7onahm/bawtpHCDW8j7mrfT4b5u8Hb7GBCROukCKqHFpsfNx1
VujvvchBxeJzh+/ZikQxvFP5OPwueKpgYKd0UYzUlDQ7xolPSjwhMuYZFFIh/8NqSbfVqvbFJ0F9
WkR1UNyVyw6Tg/hgCLNIK3tPiFcUfkUktXE1fudvqJ78vQcHPlOwTisUq88G7s2JepksV7u3L6cA
TGz60Lfed+zq5sYlwQrg0KCSnL9+zCSFGh80uY4EaxnO9zPMcR3Q1PWPaohraUMTVurCj2pnPg8S
gO1/RAQNW3r+oN+jYStiEsDTmxTx816tfI+hkwuNwjlq/N03odEV/4fAJNNygfbnXa2RH4PIkxPb
Bo9DiC0yfxzp1x0Q/UH6sykszwdSl63g9rwelRHEUZChSl3bCY16iP5TIlPlscQH/cSQRhSoWvxy
1WzIpZrFce7VUeS1OveVloI8QzveLB5LwqVdr+Zuz4zVQ+1/bKJwn1wq14piKCED8jTsCzqIcIsA
XLMnX7OjxKuiuUsYxS/bvMP2G6eWfz1QjEOc7k4dCXml+gm8DDa9CnwLEwl5tZ2/0XqxD0VCad+2
gX6MmrrEcQyK9/xDe2GtKNeYEJN98W/+PAZAoJ10kigd10i6//xC1d9yZwQmAlFvMeJsNDuUC2CM
577D3/XXv5AMcBcpYt6hJfhMgnNOdyczYKYqGqvkp12xUaQvNUzST+R5H+9wlzwZSMYTmU5AANlH
0OdgJoY1lZiLRzCAgo6B6LOa63F73kdxnwPT0eY0YRCh6KY/U7jkgddsMTZz0nIWCDwBjIQE5/lr
KjyVCaE8Phe3ZmWwDy1Y0OTYxH4I5XQq4nNywYJnMMO63DSk5VWngOXO1zrRxx/kGu5jEQfYpBSe
ocdK+nModo4m4gIUS63ia+54c4IDpTfXIU2fvbe4+M7NOcvj/VkjUNu19YY0O6aIrojNvaaCwgq1
NfFK8NOSZ4SNHI6HV3fuEe/xos2X7oxrkDpMxt3C7f+3PYBUNXFqMD0rTtI8hs20DnvHsk+yET1b
p24GN4qrLYsejA5qFLOvDMf6XNNUgg4VBoqMZBAI6xAnnkqRgaUzsNSATk56RTHIXnMNDTfvrHg0
mDUwFgAONzo0k5wuQnkPH/UyJmbfzcX1VwnMM76AgoJlHC+uJ+62C2LZVG6W7XADAg8mkl5eW2lC
UOZAytlblTvZ+ognZ9A2jOTLGQIl9W1zvP2LSCpkZrZ8Agp3+vknXnfYFo7yR2xCuqrHQzwVJQ+X
EAqDrtcXU/OU5oDZRPgsQ8zZI2roEUkpyywGI9JappxUdBK9roo7AhJ+TlUJM9aMXDcORLee869H
oORDF1fpo2Y9YCCyBNM7QZNEPKFblHP0+MqgKS5Hwzy9cA8ordi5I6FSjxB2ArrPqW8dlKKqIRd+
gBqiAe3sT13BLK1v9u9EuCxUTPFKUp1npxOPRriu7DJp18YBV5y1pkDFW8NieDt+8CGysSo2WH55
7xHT8SIdP3UN5B5IQ68OgVM9puh2S+kA/LtEmj94tvJmjptSOt2j3MUcAssc18DoDreUgwfdlif1
9xvZisZzHYbXRIMmIcMiKPA6orFPP0vDZBKvOXmVHuMf7zPGiDNRJ4OHmnfTmNi19hdbIfQ2ByQQ
qOXa46E5hpZpf/jRqMcNTrSFSARC8/SWOm4BGmp3whVRZGIHsCNZgcQak53M+4Hj+A+lMeDp8hfb
Nvd9X4uJ9wL2zTnFO4Ju9YPDkkHZ9fkGQbGNhRCIwaqCY5rUZTrgNH1Q16bEcTYxZNXF2ngLE1P5
7s+EHkKmt0xA975L3eOszaRSpb+aoerSSC4DdNOPz13pgjzvcCX9RFpU2UYXeDZtMrVyyrhk1ttS
mKpvWBUEXzIJepgeiQ1JAiV6Kj800Paz+eEWuz9XRAjHy1U2UQW2mShVWehR46mI+pCQA0kY4n/b
3lj65E3Trlgvirw26MN9oQfQWBE860Gj40wGMzLdZs+YYcdMpvwkDnmiFoYKOVg36YNW970JUXiI
KWSvEAxqZ7TXe8g/6VM/AHaa+S9UTv7Jb1W0wF1WGryDD3GqtOi4ECvn6Phg48gPZXlvTzt9coco
ndEKpApVRkDhzsRj2jaotGuALcxL/ClL+jvJur1ho6cnV9p0ZHXMpdnnlfHVd1pLOjpwh7wJk1+p
BcDVY5VNpBy7IH1E9QfHGiTpHYY4up8RY6Cyl8I8fJ0HCQ49HRMHmay+JiUF6RIUsulpLALxdUiN
Tvi3Hpv5w78ZnFIDIAZlMHuSL8ReWlKmimlZ8l04up1aIdtTHd39HTZigKzQvkANyqaPDeKZtMhg
SfBbawg+Y64T371xME+riuTrSAbtsb0JQF39TYR3D9mY6afDTizZ2+Q+1C7MrD31oLovt6EpbApG
frX2vu8U0WV53vSaR9VDVJR/YNzCVCqg5RVRP9n6En1KzOx99FSTNWsMQnX0vpYV1HQ8Jm8mpvnJ
OEEliXqQEjuYqdA8uP5k+H2tTra82GWx7NzFyPq9VpzkN3PXs83bjGnL56HPCxD/VKhlTpWMu2XN
//RgI0B7UL6VlSqbI6LVOrboCj5dNe7P8acO7DcMG1b5kM/0fL+d5LuNqMG2sERlhTLpfqNbLyG9
ynjPMItpqpLQhSbj1pJeOOeplnbzs1KYLIfrXg0h0laGfxIzaWqeqqi7jFjo/r3BLg93UaB1Dx44
pbQ2WlxJBAgP1lS4PF9UIjJmMoPB+cl1oLRcHAwU9Dn97gnwxB8wP1+jQpy+0O5pRX2ZOVl0vqgx
nS5mrPAC6HiPZ0JgumE2eNYndtYfKZIqpxmTLLOmMXx0Ms71Ny4d7P2jboPrs3WLQyILYcMKmw7z
ONirWaZZJgzWqgPQrjwdHbGfXXruAr9sdRYEbI0LNHhocfz7Mc4CtlaTtDX0y6DaPOUIK+cMObkA
IpRrWqIsfCgJY6mMXhr//IrDGGCcOoV/SOGcOGEA69ynOWCUFs6qe/q47nIEbe8IfQrWQ/ELbCZI
RxyYtk6/7WROR13sNSG/5f2oCNqJ6Ahp9NPHa8mvoPPWFRdwsVRVcT8CiNji0NrQhBD2w40Al3tB
oxiuL2OUjk3bJj4BxFjYRfQCzoEXeyetpDqaH9DL+e0OEFDpXpb/6TIG+EPUz1vaysRbJkYIDrMQ
NhHVn/P+q2tHxcpGmp/cVatiVsdTFVQF2nKM7yCesrsOYbA6Hi3dxHuDOX4PelPh6GXshw5RkY3x
+nrEs4sSme2+gfFQiFm3sYBRPx3FoeGBX+zTH/VDN8wYpLp+fyRsgd312eQ/PS2x1zIHw3XSBhiC
DIb9S6X6Ml0BfpjNEic7exvrScp6HUrho31T340iouHP1G3S7/Rhmuco4ELtrgAL0YmhDblk7CFE
wZA87XuGZLlkpYMuzr1vmQW62V58yP1ok19fqJCDpQyI2I904u6Di8Nrg+pyBp2rhwGjSpQ+M9RR
LFmjrPfWakqmg+ikMQ7MDhPqxVM6gy82Bp1noEcAnfn6GFw+ewD7KgpI16+WCFvHY0pGPulaKNRS
j1UnbHsTYjnSAikAnMvBvxb/PimuMchufCX63BELq+LdhcP7V1/3b5y2hBaCZRg2ujSjykU4rB1z
njMc4YAIGMVxJ1oT5JfXnSahOQ5D/GEjvuCldsZbQlWKHlEL1k1VaC8qW0xPoESpDTM1wFwUsD7l
YogbgnaiMIKk2+sWgsD/S9eaJOOpzvP94M0XNevwMXVAGoS+WxCG0+HiSGRRBrDpsFkP9Pctadzo
yeoFxQZeM+UCMkoUoYWsIj3Gv2TwJK/6GW8NVFi+/W2umFF3S+f78dYQsI2ieDCk/dOJ/Fgebc1p
HOxt5CeUTzE3guaFfgHHCJqL8mWcFU7zXMiQqWyq1XJ/5h95v7SK2cqZJE15Cyqz8zMS9o8LBPHI
nNlr7OQLWnPb2qazkkZ7kqktwaHnabmzAHKKSg7t8EhGm1+8z4YWnw28xSakQcxa73cxdICCoqnC
Q2gGAbU/UxtqhJu3EAyFlWMgPHll/xzWtCRIKWcK9rKo61CIMpOE+pfR3e4+jERnfRdsDn5CEBag
UTm6fhomsKNmtNVXvO/gVPQktJh2ETyPo5NzD9zIRIL5I6Qn6MRT1XbwijizS6qcbhMdGvHYDdJG
1Lf64YPm81CWNERS+QoViuNI9Z61W/S2WiZFv+JM2pR51aduOQCslIlGwpYP1RnrDRdEDF6FzJqC
NbSHxvdy1D9TmWntJ2MyI+qLTRIzz4Nrip3/BouvavkepBDUuG5U9bYs1+nGqpGVZRON+AW15Ms3
SHEWvrhRKFSRGhJ/3RtC7khX7bje8N31JyRem6Lcv81hQK+M1IIu4WGjgtgcQvg+K1WwxA2AqCHf
9pvvuYRsy1Mjc2yhfglimvziD0ogOJ72YOh0USplTttI+Me9kjkbiF5DeLyKnoj2GMpaS7mtKk94
tpLeTCToXUI+4N46VI7phDsCSb2MyY4rKPU9sCM/oBBzdVZlmTGnqtyi5ynkvg4Zhaq4/pt0zo8I
0jdaGlYcopf7S+QyM7TX5RArjXCNNxX+x/5WonIrRlEKggS/SYLkxg82b/GNV7KzVZZ6DQYubXdQ
vBDw3wykK7Y2NHk+QnoaTNt5gQdfliyU44EZlH+ifVt8u8nxvvS2GNeDu5QCfzp4CkUXO1tqYfaP
1H0XZJmfY+IOhJBwOkk+T9vV6VZt2Si4hw/wkvj8K6qiGFr5CDxAKT4t5sZWsYaDwKe3p8ONJEdY
wtOFVKiH87wT7iJOUprD0qD52qhsHtZa6yTUR9B6DsBUCHtCOZbLResgbQSfebeQtsS//CNrI0bC
vFn61g1efJx01MIbOtZfM6bImIAtPT6xuSwlHLUkxuAgMWypkf1TJwhrNFxiFKkirqi8axQjNcwc
6p5reHqCxtrgYE8VyHg3jvCDNMdUplcAhDzNaNWWUdW8RglydcCbhjfz9KobAqScssGRWVaRZF9S
668DT3fIbWj7Fo5m/CrxliRpGVFGGx4kFHWnkSjscofqbx9B0ViFmN2mDlmbu8buD6j3607HKk98
6bdpqKwYJrCRG4ldtsSxUySIjjRXZKr+Ans7DLw+QeLpMHDZFFPVwsgCZ9vsALiEVwKO9whC3KCu
3VvSNYkNaLygtq5DR9wCDcyPzNDy0CLk5T1FkHegndwMszOp9IaU3gTcy2hGqPyVJ2SNfXAYAxTl
grZzJl6INf40XQ2DAI4UdND4WsQk3gklhN8A0uGpeL6bBfS1l095Zk8b4QtuvXxMVUqZg6f83Y34
GilCjUQ15HPhKy/Flq5OUuAkIyce44Ps8Z/Au4wFze3jlThx97lufr3Jn5l1t+6UKRozpX3AZePJ
r1UjjOKnyTLYfeh348ZK4FQ+9AtTQoA3fB+H2zwSowTA184bzve94u9RK+yVgOl6O0EXFr4Q/3FH
1+tBWh8MPLBXfIZVHUkT6qIDwgwAmAWMRi5C/F4vozABTufyVH+e3bDrYR61YssCIMzWqz5ihfMG
PfACBd8/t++qsItGvQJ7daXJf4nR37huPlVv1KNqamimh6MWqnW1JYN3CSS3FGX0E4GmuskXDWjk
erpWtJCRHKZzzcnptp/spf3jF3xi5xcNFyllZA9e/Gr54slWZWz1DKbZ9d1dYB2M7MOCcRXAwHTk
kh8SN6SnZVigpCR/PCmOCzUcihOGQJjNX9rZuuJAZ/ul60pO1hN7YvjNFaC8fioPejdplvTF/PnA
OtV5VxiZEyKd9gT0+wpm59JKI8Ck5fUC3Sv+PRJ6LTxNWAQ3mltCg2rPrtzJNSrAkP510HpeWrzz
In0klTW7/i5IF/nfH1WH5MAOSp8TxNCipO4hFE2JKmRVHQ6CbJ/YO1pHJKaWz2JcMjJHpB1E8ZXJ
Yetm2iOvsIx3H7V2u4i2qYJdkd9zRRQ42Xc/0Om9J3GDxHUOn21G3AH2BORh34t9m/Li3wkznHXw
tKTtyavkfx4ACDmYlqvpwuc8uSEZZJsjohqhJFnkf07U229KDbhfhYZDXeCV9HgFKXWayz4AH4W0
xpmCiRUzEq4MvwmEAXhNFAG2+OW9cDzEdoOqa/lwLn3FPtMA2gxHjpc2n71+kI7Gc7V9m7TCbwJa
/O5G4hUDBHialFneoPFiALSPERWaPJR2EbowWvI7xPtX3dttoKPhEjRSlWDZRNnni3Tt0kFEn2y6
x0Rex5/WPu1z7kS/Zdx1my6QsyjjM0K4i0Ll8Tc4tET3OYrINWy3K3qia5I8tlLlpRC6IZpZ7WNM
rkJ+hJPHX4VDbYRBVfIXTJ/lMSqn43LyE2AD0u2oPV2BRdJ6UZf4WhJ2qPsbP4OLH4XJBpBJhyme
nxp8xlyVVj5zi+V8Q+6aGWHhRX9XWttX8VlN+9CZjsiVLvdY+QFsoCY4TmmDDMV4x9V2xgdBL6h+
ItN5OjF7Y52YScQGdXiKEWlbdK/Ww7wzHeQhPt7XzYp9TL9uH9/xkTDJiFh8ERVACI6ffoQ/C03P
hDCHigJrwPuzvnAga5cqqHSmmSxTXmVJEBEpCLkClIvmMZfeWDJs/0hjUv7eTetA7WZTSeJHQBrW
ls6qiTPAx7cS2hW9ybLba632wIQIdnhPy2hmuR4/2cQo24/idUT1bj8Z9+hbCdwje+t0ZSoT6dFB
AQf5i6+dnJ8pzBFAe/dEbl2fbD9ht24OWheSs5DB0HryVFgnmGFPi4p2X/e7yEJF3JT6dRETJfnu
rk60oKXMEXw8YYpsKtfPyxR2raI+eaavKqbiwW5eshZDPWeYTR/MD9qn41h6wqjhgmC6QCO1OhJU
8HzHQLpQKXLdWwgoMjawa5X4/l/KsemKF33ZIfvKVxEnj9QBlJaFfr8IAHMLTVuKzkX0u5JjOcu7
D1zK4iHQCWy4rbtFpV9yH+u9sDmC9nx1JBnpsF8TVYnhB7N4DD1rymQMla2Uvawhq9EC2fTzUNtb
VR5+i2a8NYiPUxp4BvVVJgekEXP4uMF9M35R0nPb+tozuEBySQaxGUunRALTy3rCfqhJqNlciWWm
DADTEu3Au+lanOyl50mf0EcPONhK+JpG3SteYhj3GZukb9o7Ilf6IXPS/pdFh1oZtvsx/xubYVB0
+ZMLu+cVMBYNit2tGjoTV3CU5a06BVICiiBEqKnTjur8BKjc90tbI8jG3mVAQVS5TlsNIq+PbEHq
ppjd+7WuLKxmDXuA94q/yfNwt1Wct9sjzzEjVgIOTHOh9eOyAb07k0IlU5J79QrP4rDyAIqzRqYj
ozFOKyvnRn4uKlzsxsljd//LaIOKYoJGXC0UjJI7nYt5A2fgPYxB0XrAjV2Me7Kxzxdj9Ix9oW/v
F1QWXkcnuFhKbr805LsspDeJceKghB2/dzsfze0qouXLOu7BPg5rl8YXKvufbWLLCvptuKla+/KC
HtcEMjA1bRWvGlg3RSQNvJByVrSafOmw1Q9b8NPOntTjJdTXtYJu+MuQsIXwihqIBEeCxypn1pvg
zfTNK6YPwQWG+hV4xPacuZ0teizYdRoQEOxsEdwPq8GjuGB9gLUjbu5lZRHfq9u1C5URkzPJQdP9
tRZHLdMKUwbi38N3d31buyu4gq7JJEnRGpaz7v47+t8DxzKt7JuEObaZWoYJFChVk2Lz3jmKTo7x
fawU/0QEWNgcOPqU2qaIfxhULAyufnLRtAY5BfRLvl0gRkolTSgJDRh41MGy9VjdNoEjnp2uQiWp
An71t9RtcF2X5OzaZQIRTVSg1Q7G/S1o1aJf1a1ND5DT+dNWNxUFCARdJjzONHoy8zcFSFBDEntL
WgS8+REM3tCMiHWgdpVzsQXqCcBotOb+ADsdX+pDbj+fW3PFJkte/dnNgpiJg4Xhq5yoFCAS/Cw2
eLeTKKB60W5jOiFyj9cpGdGYNPLBMf/6lhkRBWZqe5Le2RWAYTnyqGeSI/6oQw2rilXpATndnJFQ
m9hN/BOlBYznK/5YY4CLbCtbBpE1q+hfICZy++4MATNmTxUYMY5TJ7mgavTFRqWaEekCH8Et17A1
WFc7CsMcvEx9iOlKuzZQKCblvZl9k/0XULtoj5xiVneJpC8X69/J2x8kVJOcSGoMNv6QnYXEdB5T
1HshnUXXNlxoe8Fi3fY6hBVLm8+Uk3hfqfdUkHPArP3qnbDSuoAyOv/4dxSjCqYZgfyFO7WMTPD5
cHu0Et5cwfju9NPfgi+Lp7mbEITwLpvvnH9u/RHnDcjG4R/4cyarf4QrG5IBRKylbsp7cOdFH3tr
l/hQn8k0+JXOl3k/e79ilUF9pKNhYU3nsN20UCFCSnK3cggzeOa+C7l4KgFGpKzZEy9zk0bgpuac
Q+P3moGS9LJ8Atm+6KTfwnBB6NIJEf1uPTFKYe4fmthB0MdAFC0NsESYQhhMLa3I0E1f2tiRDTxL
Uktl1XuGhNnFxYjK3KOOs5ZQXG4CzGr+4d+Eq/JPBOprtM3e70zxRaz04FRQk3D/NceW2v8PRlD4
6WvnHWcUd5ljB9kEX2oppOpgZiAfvvxcvcethHvJ0W6p5CS37rB8m3SI/m6p3M54LxaLM8dorFyL
7NgTCGzU9lQXnNOejhsbcEOr9q7GRLRhtQ2Pw97G6kzhthJkGOxTDZp9IyYySYp1leF1SQlsebLN
FERHdZJxuYk4eZi9keMvTwdT1zLzDlRkuaD4TdEONwPeYniuutL8xwivSHFWp6i/umj/FCXIE0bu
vuEguOj1qYPCgVl8Mx8zaT7cizu5g9p3DpLtMlkKd6kO7KAUrIQN490SRsA/vxkcsm4ee89IdBtz
zy34dYHeJ0TpmwyPj8CJ7V1m4H8p1/T8kT6/gRLR1vsPUCo90VkF1pmT/p0mDYusdzwGkANE5UKq
QirC8wWHIB3LeWonqb8QFIv30n8hsCNIRXiJoUJ1Q1MVGxXDRdHdYsbniCWDSBR1TgIK65lr3iG8
UJ6rAFP/nH1GQQChncIcCt6af/HoXXliSGl7Xyz5q2jnu9XGvCCSgn1HgtD9839ULRb4xlpoCwag
C5xiMdGNwRldiLnhuM6LUh1oPk4NsQGL3vcRk2ACg3d+njp7RkRlMb9l6wj+viEHd8Fbqh+UPANV
U89KGVVEAWBsflc08nSxIfrBdGY11D+ujeArVnAiDrkly5/Gl9FyM0lc5nN7t+nHodisrtLOPGEM
MsHcdM+VF80O0WIH8TU7xvm9Ret6doV3tibJW0PkbDFkTmdSwiClJ9QX5HeV4UOM1feoTZKXvYgt
yrB8oSNUH9rRGiF1OcBtsrL9JCWrN1YFWO/mRUiSuaiRKP2ZvB7Rl6mEcnsRbrVVa4PxuRK9aopi
qisRKKwHriwZRn2rQnUYbFajqSIDVHW1e5w3bWVSrZEsDvyPqhTQNdiSNYHNhSk9R8aiaAIKyuCd
GPAqw5q9WZpP6wOXfEV5ySHb6dRPO0SlSlVVztydcVNM5SGlW+vDHDjorz3F50gHtd463JYTj5n9
wwJGhj8kh8HVZZlslW/wsfT9lq8Z3J2d0Vf2PXWJBs1q4VU5toM+jl8jXoUBJtCfDQLJCjdqvd3e
e/KZAluAyglMQ6JKt0UWyE79pb3rifZvE7AA/WkuCmctXUeBCOJFEBgRpGB2iXLrewS0N1hE3KrH
2dRhhM5DtRzcMCjhKP3PvO2YobD3OKhv19CjhUHEnezAeLnov74W0JAtOTQ3JTZ8jzDD6Z1owdNd
iMfEHh8PYVHxmBeoHJXjqnJsjs7xY5iAwnExIgu0lQnAlMEq74WDYSKdikVOrHy+sek8iQ+ks3Q7
f/laXfqbBl4N2Cx+TZ/2BdSS5a76f2ViIiPISSci83beXdmdc3YH129EJLcvOMuU2nvWFDItBDmO
iX7plywu0H48HByPR6Mfo8ftxLY+K7jhrrT2wlzCyZFr/SGQKRcBMTfO1huv8AmPZzGKR2lIDkSI
gur/7aAUQQtf4iRuiJ5CVpAUx4u+tkysD+C27xzEe/F/wtheKiJzu6ah0GprlXc0aZC6yFMjtChA
HL7gU79Lz19+AY8TaX4XPJVw1dDl6YEU/Ld7ZCQtTaMqahsZUDteEIrraPzVbsjOqWDcvyDyn8R+
RyPoYlSWN34cgtE8o7nhOGIYtaaZkfK9LCU9i//pc07NB+NdddF0PzoMGX9idczUyhT8t/zAr9oD
fmzHJWDQl1m9FJPdPw7iS5i7apaiz5I7f43UJWT9tkk3UeRlLv7esJWclxXsA7ZDpqU1i9XBnvtz
QWTaR98E2aQAvYY0vnI/HCDcpdiX/RUR8j5FBXB/G2wZLcSAlFVHXvFnl5r1U7du7x8d64ZMHIhI
v9/hbGiI6NDKLR5DsAKmStpEp9vYC7LpC1C1FXDLmkVdZo/SptdzKsqNme5sOH668+R8i3rXtn/0
9lW+eMu6NTfVSOrEM+pHOjkB0Z+4aZec9p7xgauLv048oTLMkHuJRWv2vVUNgGeLytVsRYcyUBYD
cxj3hLJteXyfsotZj5wgCpzpeaZiKVF6L8opwMQKJFOi2maP1zXFFYiBb1vjDzz4Cc0SqKiBb2vw
eJKex8+iMAQfsMtRIBysD+TeCYsfUPfnr+mSafnCRTcv87FAh/wFBUgEY3jTAsil4nL2L8jks8zn
EiLj4+mluc5ZQBL6b4PnT0fgeZQ0wTRmmUgPvogXpmrfPBMyOpi9q+hSSCOpXc1YcbMQxz2E/q5X
yIg+uG63GxOvXwsKj+6dIN7t/84pty2arx7y1nehl+0f3UuX+NJ+NLFpF4qjessC0Y2qu4MCXvjZ
r08c3k/GOPdUiCBsjI4tJun81qaLJYveT1eOHUZml5gzdHUiAUB/O28kyNPJc6tNal8v8jfyCFSx
X5UT6GEF4ELL75WOsrQJ+V2SwvU/erL3EU0ubKKgQfIDhkSoN29NMxZW8YPixeFbEHcQKvRehAbQ
JSO3ZyV4dEm54ZmCADwJj9JzW2274zCcBTqEx/f3vv32CehN96CKrtQpUqug0zgfWCmCBhyiF/42
B3r9Zx/chuz9lLKIwKUSqFCI/qC/1iRmTzznXw5fHTi54bBi3HdUVW+gT4UVrVJbJJvfJzVu835/
dKgTrdJsW+s/BO6HUQs0AwdyuenLx+CU1gaUdeazxMUgWZNf56m+io2jdmkNmZv6HM/AFP6293a5
uvbS4YwtTbkybVf2lkVw2BUFCHgVmP9g4DqnmmO42WQlH1ynhyhdNPqB2rERO7/mWg9+5CQuehN7
TKe6H3+k7Q0A4g+6lVaoVWF1AKwLcXxEV/172mtKX7MfvVLoNU/EBsrkGptqeZ/uXIRFhgFf2/gL
dEy1PZGeezsaHkpl1spfijsnbUzszRQ7KBypk2Voo5uTwEa5GtxstCJj7KldilX1D48P7O2TIVBr
9UeVJVketdelrF8QGsHokLJctwMi+3FxSMGYMylQcOphiqHiyZz1/y1VNoEvtLJxhE3qcLlglRpq
S0nEwU6nO+7TV5sIHQYO2EkrYRBJR1YnF700lorhwt50WUANMitrkPu9KNn0G9TBNPKPItQBEm5y
m1BrfAgDy5uWCTetzvNGsveY87SBmejCcIWnU5DW9Ootf6jWOPR/UiAXi4Bl4ac0pCdx5PhfiumA
paEhCW4h1ceDYtD1nXMT0whgHs/JDzxYYYMaU/3WG/qNsF1GC6UM6S1hKyFXQw+Jd5G2iLh0G4cp
6FgjCAWby46jH+ScQawSeaV3Ap2evRU1qwJwHm8z+bkynfw+xcPL2EgdPZGLhGp4axSvzvTXs7er
q0CglJZn7VsXYhL4nEhkicYOF8ir+noa9nVBPGM1hCU7x262m3U/wkCTaR+0ec8jzFyIlZeUC1sE
YVJqceYoS8hI4DYhQg8+wsK4dhQIVj1PlsgoMXPraTEU5uFiM0QxpjfLswMo35+g08NzfguVExzK
PZGIZhtMDnjlkfgkDTavujFpxWXJZESMPjNobwZEd9ah9WDuhCrtR6sspi/G4HLxdfeObkpa2HWP
Oqod6kGGrT1moEKuZzbE+yfHGcJM11XTsQoEMyNqvRiELxEXtRN/l488T/tokAWvGNHrA6pxugk1
44dDGRZKqgSjD5ERSAqXKrLss92BhjBszoAu0+e7D5Q4qmazXIzo6CYvYpocSe0YpeRrgHnBtNrt
NmdjwI3z7QCtlDSh4/TWKuOEs7Z12RY9ZbRgyuPsK3mhN9098IBOpjNT6mBs02dVYxdU5c50lZ1g
FT0ORFw41VU/ytdLGfiRXvg3fLV8Td5t7oPkfj5X/n5PwvEgjY0DOLs6HZ3ZF7eEvRq9RVD+l9Z+
xRYpVwixbPH3eOneNYrpmAWK8cE6I44KRY935wARySeJYpLDKjaWFi7d2mHhVkXvV4g9sTo5hPrB
ZmUgwF98DmK5boxdCE4PLiC8xk/onGH9sWtgrIuvXHmJnLHVDTYRuVoymjh8NvvgZUlI8zcobImH
hfxGtmz9AjQa05bD81ebwiG5/Jf4I40045leczND/o0MYICxI7a0WdnHhVpU9g1w7lNslr5oRQBg
ssac28N97mCNlcghmJi+QuSI6GRb3IUbLdcbLo4MAk2bXGtiLJznWJw7tsb8CUPhAMyezPcM+4e+
4XTHB2AHY2Ly2ITmW+SGafd9hI+mYmVKlk28wa9jLFaTrVhu263+VRyG8dwHtpGt1gPIQO8FNx0N
A+kMIdTp9DbbdWoMKm5lO90dquWLnLBQjmRdTmPwXqZZTqKEbbp9Guv1zM6uWQRy+YAamxvJ2DpF
E4lsMjqCRug/V+nY1Z9Nuq3y1Z+tL0uVMW2gqUEi04ouwrUV8oa/rXXcBS76xaVXO1esMFEVb6E6
miYhnYp2RY+Ipfh1LxcSqn/yH4cuj2rac209K2mxAGseYnHTYH/E4chyRZovaYUTPa81+d3oPOmD
EdVX5nHRilwVP137yxtr3hwoZBRtUq+PZE/JFNnWWOAwswdJ/eg+Yo3YvnUqrKDDG5CmKCmG+IR8
uLJmsUZ5DNL11nEHS2IOl9VNw9agB/S0LZCT5tsxhr3Z4gjo6n0f5r6Jvbz7wECfxwcPozFlqhWN
SdP2dvQJ9vs6ICeUAa2Af9fjA3A5Xlp5ffX5os+yfICXPy9dHQvhDPPdJPM8Q6rlRb6sg2iRkY9c
r73fO+P+pZfoilWjcWV2dc1x6MzmGYCiyRBo3fHy12+9oFMiMSF1yglfVyTxt4dS4bXHFy4SLtNR
jlgZZWGYZOu5OUJ9voPtGittnU7KpKQ3Lf8UzxLan0YGTttHsWoxHsCxi6dzJJIq2TPeYG+OIyZr
k+PmDAyhVEbXmVrMmwAKldtXhrgHeFFbBC1Jl3tHeeG7zU5g3/jd7NRDrx3JH8ufrRqziCn9SbIM
ji0ss7YnLpJyeIJECUGGSn5ymReKSizC/XXYt8DwM1po+PsHiLJ5eKW/f+kqpGDkTZK8DfW2Q3re
+PPjp9a0XG4LwAahgraI1WysIGMrtgFUdrs554FQoKUM2Fmn6e3jk2VCeuaFuJvl3iHTsegbWTvp
OVD3y/sByaCwRZxg2cC6KIbNPMwHWi+ipFi2DWgt7c9Iimx+At4DvICCqq5ykGQ30dsOM/WCs4kd
bna3jZDQYlJeUzLQyxLzO6KwD4g+XtXntVo8Cul7yRLCvc/FUG4CFahk3mXIomk8wnYDwwc3tvVP
buB2mTA8SJJPGW3V/GsF/1YN7hqBraaVIcchr3Yal9C6IoxpR0sjFaJurv1LJba6xeocyDpWubWr
F1Rjb+R474dMmTcI2d4mRKmBZ2fvXjxEYXHm2JRucp2x72JmO8tr8wLO9IXDqYaCz3pmkvPi7k5l
a+LmAljrLQWTDZ2bgFVro6l6sH25LclEiDRqt5lovfDXwxv36bw2qEfIE5kbIw0ixr7GeLWKLXNJ
j+gDN2LhZua/PEz443Og4BFVTwtpLecGRElD9FshjI+0M6X1skyULGq1Nz7+qkRmz1g2EhBsZfcb
ss2EzzFY3YWzd5if+I7lr4ratD8T35mJ2fJuc3cK97N5+KBB554kCiWCRh0Noercv6CSOS06x8kC
NHkwTwuFaz4kjRfslfvksAHUHNAsz91chXcj2og7vKO/1W70zbWMBDYw8Z4O9i4j/37gyKdVw1fg
/JuoB8ikGBr3L94RQkukT72E0pi29sloKAmBHSDumOCMxEmRFA4rn76j7kajvTSXiBarwXDYxReE
5v04QsnRVQp5Q3E1R2FwxHpcHkLeia2NBzXTko65b40VaPV/CU+YqKjI4qf7XtO/NBAg/4AGQ25t
qGxkkuUiGc5ujjOJQ5xWz8lYqAt/JlNJs7FKmd01SPjHnI3GZi/8BvSxriydboxcQ68wS4wrJlGB
0dGc4wrG1a4clUMGQmJfPy8gs8Hps4R869/HhktzmElrVl8lJCxZRFJOoEK9Px3r+rIhWz52Ko8E
v85lvomOfjjtHvPl9H9ogHvEhTvslpwqtHUV4AjyrCkEmURifZAOV7ILN99+5GV2yCxCc0rEdgzK
GMJKJa8wMFJMukbdtnE+Vv89GedTZ1b7bIiu1YufPdMryIQSKkXyH0SxVhitHOhQq/Gga2cH1MOO
oFoOO+G/PkvP8F5hl3m/OQR++QhlfbNdksTVI6uS14DWTZ/ebelyva6DtNhIV38uV5EgQKT+gU52
8piFIuq0cTcPDS0efzRms4vvHzbBbFsgkUIpfjgwdJ5pQ3pBdbqrK0SS1LW5lS7y3nB4e6nssj1n
BImIClmHfL/1cIqSDiea3rvRxpICXI6ArSznM7sgt7tgIS2ODS006HnvtinbqZyjeeOk/hiHjYRQ
qG8kRZDv3CFcyZj5RvN6oIDt9Kzl3kLai6mafV93oL8oaeexRF8IXnMgTw51iWfg532jaZwxfjV5
O6f2hL7hViCfQ7/45x0gIk/wnBWBekwOSBrc4yCHrDb+cd/1aj6ofagOL+bTGX5HAKw3horPijuu
H9CIwxoIUCUvbN8eUXQSLpC8Ca6AABMev2lkPWyn/YPtp2OCFzotFO2RqxZqVlUBIjQAdhtocJa5
khQFzteQORP7/MfNg7AGYxEVsADdoZeN55K0F6X3lwa1UpKUsoUmTGTjnPNz1W5JqUyly/oQcdH2
ybcEbuL18rTvD6l6KKc4VypcyH0755a8BlE6MBn2H9Ewlxb0sVrWkhk/R3n+Q2M2Ew8OQWduSkow
9pw+eqzWbRleuF/jVcOWH4VVLsaYlVZZNZaqQTKRO/sRBpt6/V8CoEFe9T5iG/hetmMKg1n3WY1K
YlVY5/wXYi/vqGexhzGzE8wnS4G1vhd5ayRk7ZdKcl6n5K1gOGGos8SiMw5XWLF0d38yq7jIqGWy
bKiGB/7wJqH18oWgFIVHd05/dNl1uTH+npRKJPVVeKZhfJbLy5pZk8x26HhJuigQP+GfwnAwrj1G
QlUgTpOsSEi4EzJxt9+DHfiPnAiyojZjHRqaVBDNyPJk2+z5yyO31GOkjTBLxEzjo8bBHii1ja1D
pr4f4pdveamqXyI48Oekap4z+/INCby9fT6CiwWo0lHsB7OFSQWGwfi4zCDQ37xGGYdwUMpW1pV5
qConz4dlzuthZUvy+VqfgKewc/BFZ9qtzffffBAzpnEXiknKtALzSUH65zebyjbBf/gJDUu6V4+u
LVB9b/RAn2hG1VdzRf2yH24QnoswqkfmWL5zu7/pGq+ATL0uaP5R19PXJpsp1LbxQzPcAC7+wC/7
UK/MKOR8bUZRBROGYQLQriizvEKaay8CaofG8uRlRJD9LoZdmcPDeGdLik+gE1W5YZD/OQud7cwH
iSgedvn72Ddee0aUQ6nZHghzN23FeeHeBiqCd+JxgfTOirOfzosIvYWoGvysgP+uFLqKIevOAi/f
rukgQPJuV3vxJ7BNdA6lTLNtBXnuiq+uXl7MAliduCt4WRr2EhR/6/6z8t+AVY8YdOiseXAjC/h5
a+TnL3NTzXRfrPN7PbK7QOWz1HXmCG/PoJWH2vzV6vik4UzS8idBnbvd1EkMdqXmHYhbNyLlTWs8
neQ/kLF88X7QlEwU6GjgbapR9uIV9ZDKTL8bJXmnYtUwEUZtSRTytrrnpKQRUhQor2P8/oMeHw/v
z9UOOrKncR3mdv2hZJwOx7wAGolpHUsQECb+pidYcpHRVB5+ZI+zqX4+jGg8fpJmirDcMhtSB142
CIzUSgF8KCrSrxMXCQSEeIG4ZYyCsN3WpBsYtUubwKfcWgOkwZFdzFYceSC2EGGZjJaPxdCX1vvC
45rEUI+zPU3A/FxTPfmQ9lr7gmMcXBIiD8NgB6HTDdka11v5GHqybNEXIuSTvFl9nsH3irl1eq6A
WWElpUz9oK5c31uqchMWkr1WdXVCXrrsQ43XkQ7Hxi5Rof/F+zbsK9Vr16tLT/+Sni/ezH3jIvKf
u3bhB/53uCuhTP9BVlkSK/C9ciC2LYnfx0wqwAk46WiOde9HhwLj/WB42jjBxMgKx/erPy/WhmZc
i4RvqM+jRsLvwTferfzY88/Zp5DnT5bAsDPRctc9497Lf7RH+AgikPqNh5dcNBPq1NyTGmP4tiiT
zvxkwWz7y2+tMdPSyz/fHxMIuM+V4fnYiho4FcX9lBcvbSDFeEh44f1BHEJ+iz1my+kwXu4rYRyo
QsI74RwMWcz+oLjnln7btnkFMYNVHe+w29rJjs9cc6db6hJhn+q2sxxNMNFc8tVueFzreuupEMXE
oEgCXVEHC5b1ggOGJb9+XuHErlxTk+iC3lvtRb8OQxtisIcXD9ye8Mi9ygkztaDD3TDMgA4y1tOj
YM+U8VI9It74FYfuv0z9QDdLJZaWvTIYyWgX+TXj2jqEYFG3HOEcRiSWmZpLxDf2qSlvHTh6tOuL
DUV1vNoHh02PTXjmphjizmtjcA2RdOEjTpm4ht3IlHsFw5+NezYz9n74c1emDVq1Cpe7GCOup/Ho
zTGph7HT8MWsSsYuaU3IRygbBz+JgCWu/2rJahlWhibznblIN9w9eV84X4sobNc7Pa14qugOOn1p
XMvMG2p95u6bhCkLF3jSmLSHhxoERszwsezG+wMtA1QhWsKZ2da8/GKh8IWOXsZuMxFQIAexPHVP
J1UTyALCVWzDDO5w18BULB50Ex56Hi7FUHPRBWFQgEIKaNVusXcgMUgV62TOTww56X/t5SJ75VKX
VYU+cwCFjVgmJa03T+XLHgXze3WLna5dDOswAtdWDMHcP3U/bibSuGIjU2O8gvSnzIoOLMUZgqxz
+LvMdM2NurahIOqWBkRSc1qfYu6ewZZiqL0rSSFEpVOCis3vOW2PsF5ZJKVGLtP3qONpvoEhOMQ2
9mX1hqxNX/sPVi799hr1Xd2loP4EhUzHgHkJoU/lTgwvhWEuN6X+CfHnZzFI2eX/9AATAE/MHyhG
SKmE7IOZj26aR6BqTbly5PxTJT4DgC9ss1JlbKwuNHcjT7idiheW/HNJmxCwpP1evpIsIulb8Itl
1VkEmc0UP2vzTQzaOtyRDr3WYzVFE/CrHgNKOK027PNjDoq62lW4SFklzw1w9boqqDmPLWsHBsN8
oe496zutDFslhv1ST0885gXiSJo8JFj44vd3piR2xvf26cidBTSs56BvxQijzMN7OSbAD1SqEc70
zJe0g+Z6eZQhNHkwUAwEfZk88+TFReFwZmlteM4a6Sl3BtZeB5nEuS9YAAPtGlrhVHk1DK9XTmPh
+7x3PLBLwNWb2+v2dmnh5uplchyNyFK//oyf3v48miCVfyoRCLNdC14zGlJNXT4PdFvUPfvBBeqQ
RyqxcjGRyW7FQK+j6a8mphO71VEyaG5oE/m0lvY6If5fsB0hw6RXC9z7QwdVP+4htk9tEfnjtEfG
R74hIii+McgBxI6j+yegsq1zK8+0/Alumnwffr1L+UPBmdwlnm+g6PNVpy/8NV+/4Ws6vU+NS+oY
a1Hscaa01Ak3W/wc1/HNFel6BkG27ZNeb3oqYlhPq6bCRmuWWmRtkqA91xWO7H8t5V0MlBzjIkxx
hoxZzjXnziwaQtn37Em2GBtsP0AAesxP5821jGRdh04OaqHnEblmQl8sSMhkIlB1B/gFfRutXBKK
POCLL+Wp43RaVjL1gbCA6JTHBMq4nlBUV+s46VqQ5V3SRnCHnzEP4fRkgeDyDniPTkOGfuer/iQn
4D72JQ3/0km5M8ASc+l7lplJ3JrQCj+EhxqCZBh+RWHq5wBphgInXHq6SNXxqgqWT9624g87l3e4
eNvXeuePquPUsrWbZyQbC+zLsDspu4Hh99WDjNOdSA97isTg1qA9Iy8j/h+T+gHilHXjgUGMP7P8
IqhDbdEn+WYukxn3WocfZH34Zvrm9HSa1xXmozEhYgvtOUwueOPycc5MnwSiOXvzxtGUHJMDycA7
6uYXUSeG7/Qy5MpThuEntfg6IlLEuYK5oGGIxVkxKcFKHn5JBLXznmGv6o9QX3Pm12zbMFaNxHwI
QcjSnEXtslGuyRdGc2Gh61uMO20QBbSFdE7rGJAvzZk3S0qKWRiTSnD/nkpyzQkbMcSgEsSFqjKf
+A6EGmIhy8LBdHUyJFdivvc9fHO9zxq0EEda3dM58iTC2l4Mgor2b36jmw4OYv2leAhlCFG6GgSN
xxeJXrM1PUHg8QrqSsLx6Gbz+7Lpa3wyaqQYmAEtC2L5oCRDUpADJZ+tDa9YjrzYQk5tPM0WQTf2
gkj1ZoLQV30VNqamsf6DIf03UI/0G/R8XLSPNf6KBdnKf/YHv8aAVjrHWAVZKD7XjA1Lqo7M/LGQ
Bd+KFufBA+9t6N2COBvJ7+igJx/O/8JlK1fW9geyDKNfZGsEBoXbbix5xm76oXipU8ogS+RgS/M0
2BB5RKNnUTwNQavn9LLGIqFVzXD2xP+zYwzHISDcHslpvCKGL0TpNlIHlkseJNN3M/WG9bUQGti+
TdqO1ye1XF5QUksL4tG+8swi2ejjLzIVRmJ2eJKq0+zLnYUQeNzEFBQg6ghFdFVd97+bj0w3cxHQ
bKIsY5IELl2afRPBJsPTIW/cLMsnlzYNmlW52NyamIl0b1wzz2QYFkxH1WleKZ088e5DvOTsKLy6
vERWhvKRk8J4uHvsPtMb/RBEdDrfS3p+IIQo9I+gYOw/4txIBENSFOje7PlsWcKdhB2d46/BAvvV
SRMNV/t6C8np1a1g1tf0A+NSHqX5bOUTLWG6m/W0JKU0G9+Q0IKPt9NRENIe2bYU+cn2lV/AAn7V
kqg3zPyaPncCqVllQRxeiz/C68fuKqWYt0F2PFxfIkwODzJRF4NU9rOcPc7JosnQcJiWGTjghYIu
L9XBT2S5CHYe5T3kzPzJiTIHXimIGYhxTQHcT+vUeS1Yt5Pa5AadZqXTIMzu3yYf5DhNlY4+RVJq
CKuuwjYaMe2IuKffCjy6hi86Vc/wFQbILvYxl1OVaYTIcui8JIaXGC0rVXksDEpK0RaDt94Ov0o1
u3vmK+hFvxHIB841tqzLu7foIpKVNFTzXhUkRae2yG9KEvOXre6YN8M1/YVOkYRct/gQqD/X01KG
AxLo/uVEkUWGv1q9+CkZ/SmSOBKk1+iwaRrPSlD+oCuHQmyVlVcka4IvuM4DQP4ZJy5cXxgaNvNY
vubxc2HqmYOUqYW7HE1dgqUXGwRGIQj61+hmyHshc9tXigsyv/YoQTxJk2BRwMNYL/qROrEivq8b
RylqG3dJJIzJr8yxEEwcLVcJlfJjSeq91D1fu404Vbraia1GJLD7DbO5OrLo/oywKQIj8V+YZKAL
tXUEderz6XSULMyMZiSd3MlR+OyJS+4VCeZCvkvDG26G8mzsd0TK18FIszibOu2IdlyDHE5mJKYi
FezfNbDbQPZ96Mw3EHr9RnbxFLYcahsnfLR4UH/MzcZ4KwUFASxpkDB4uSU+cYOPZO1HAGSZx0gf
57chUDxBuN94PFjvW+2rp5aejuRmlGDv9xwc1cVx17ZaGcgX17tlJUpXPIK/xPZCN8Dpc8z2c9W2
tmrnar9yuzYzOgQd7okzKIqw5U5yDaRoSHHRstL4Nc8bvxoVBJ/tspq1akSpn6FbCXIwLoLetG+e
Bhi4mA0igpSmbmOtF8CfoqoIzazARhg94MqH8xu3OwTxDy0j9qVcaznQjwFPMLceF+SKZfEI2y/d
2LdEmFGr9PTcu0xKLGlOnM4iu40mk5ZjdUgABScS7zyqwpwLCGXV4QyCZ/A5QHXXDvBQnuTrlSRM
Pyk1meQQuEItOfZf7fZnZ7Ptn7imuhOZW+CjGjQakMyrNtpxcXHpGIF6JY6BwaEidMbdmTpzpjpv
xPe2kxUSQIBE0e07UpcJo1TBZbR+HmMsPRH5tOZjLE+8zjnjz/t/5QR3JDYadhfPw+cTq2X8+ppz
JgGlz9hyC2sJldJr0juUpC/w9tt5TWQrwiLYAZ0ik0I0qauaKbQxoHGbtsB6nY9dftV18O32bJwt
hMIgKPQ4bV7bmUVACQae6WB9kdK+cwjLkUg1HnfkhB6yscO1gzUD6J5vSUown5OgSFM5navjFztF
P8R1tZ5eT6AoTW8jpKTaf+g8LxbPs+jDQtwajFop+xbWftfz7ECXFQPHVe7ZgroigCKE7xvm/wcO
qK1EZtYyumft6PRvCGk9G0GfVScpMiuEp3kAAXxx5VHW+C+pOrgx2EZDhimF0X3pys67zQFq+QYR
SZdOaA6axz5BFjziPkocHsg8vcwvoP3TmsuXtqkZ4NPFg5ExNd207EuFPm6ul7EvFTixl9NBQ5TD
2jUn+LdlMkaSIn0MV7Lj9lodKkKOwSDobR2H353O+BYqOiiDYsQ9zpilnzNed23/yBsWSnr2DLus
8m3Qtjlpdi/YpaK/2OWrJs8+yTIrsvdkXmCLsokck+rmMhcQGw+vCdpe4d4ByHTY3m7rYtFApT7J
XXk8eSMbvnpXfUlJ4ucmzpdv6yVmEJqU28Cbz3FD9CgWRl3ShYxABK1zkCUWe0cnanCDLUBVaiwH
sp+TXZmOEtJmhXmySOPBRUqyBO4vb16C0a2zVNSYwR4cfJphLUqdqIjHGboCBhTHNtQ9EIw1TOl9
dlbTvNNMNN9QxlPpijyNICFWjxrkwOUmUXo0PNRDKWXQjM/KAbccjmAUDFIB1hkP/dVINowI/jZ8
nO5kg8DTwmqhPt8gYOiHPZ94Inm6odBpYVOTeVy4wxQ4afZaIDhtcZAh0n38MSeJqaX2Qx4XDrWP
Q4eUttB7xeNMzhhHJTRAXwRJSlm/+QQISXlPQuzpYuBv7R9G/UJV1j/znSDwU1vJFiSd9xx1EfhO
0CyEw99+Gv6b57DKH3jimr702klhMM4KX7iXMspBXbRJaRR7DD/LG/rc9jQFPxynJ5krwWR5qHXt
bashO3+6NvJZ74vGcOVfGbi7oTB3yoUtnj0rHcqrBkFuPp5JOBFcwWixJxGf8eldRVgMks+ss1f/
lzlGawphS8Y9ao3pNq4inTU4J3CT4IpaoguvC7vunDY58TNCyIudMxwxBNnn5aB5rMLc5FLAijta
4SKVsUhxNzfuf0/JW/FM40IqhBmhJheS5ffYiJpBWaxQNUjRLJWezbIK1NilmRx1q8CgCZnGqltB
Z/g9bdJUfdvAP9fC0x203Zyg0OQBMUwqDlx7WR78x2BH2N8xQjKQl4TaMW3FjVAcbFHlSeGXRpkw
YTPSK6ejmeiP0Bi7bzag/TSzS7IonNcvnSAfBEb8H0El0OqT5bAw82+ElHKWwxFG209mEwIKeDvs
t++Kt4z+4TsLuCbIzYrvLY9JM2LaxcGIpdv0KRQTPIYt8ZT60/bAQQOwLKuBr7HMRmKHKYwxSV8m
a68iUKe5JYduhrNw4pe8FAmgJPRjnp7mkr0GIBQSGLSCAr3Dm7G2P5ez9Z6LBeRpdZTeean1gVtq
uFngWIm/qbwKRU61T53sz4lQf0SUHypGPbnABpd08S5ztuj2edklUAnoVLpWVxoBOp+V/L1aLbag
M+l6MwbXocRut8CWoMrVRAKCngHZ90xMPkfwQpkaZgyDypWLF5OKCtQmiYf4azEkI4GPibpaYXWd
k2B+wnXuKAqZBGo5W6eQyzk8ShC2BNBVLaiwSf4yoxpFut8OTDmH0z4Q3qVWuhRO1IoOh69ZmIfG
XWeZSY1siv+wPGuA4YrfWcggQWV9FGNbz51Q8bP2NI+Qo0jZ/OQPq8B16xVHN1K9G+P7BXsYmPrd
0JoAd6WTITiEW8jyCPbbtjCHWoRHb/5Ke23ND6zvyMqpdKAzvmauoa9YFCSQ4lRajxbPVb+nqoEy
rSDSPI4Ni6piUJrai6hVlPqbgL5YiUZumEu8F+mt0X2oCeGnXgU0U1fK5dRQ/wPPLXt/iwP50UTf
bZZGBt/chz8r4ddM12MqAZiQ6wIxR78CnizIab2anMYeDswjkrhgkt8qIugyzILXO7/hAT889qfH
SYuypBB0Ve/0XyA8N8mGD+dvTfAW4hyEMwfMIDH23TqY5kEyqB/MW9mH9QnMhhHfL5telKmzKEVh
mMDa2mU+Gx389+jhJHBtrJW4Ze2msocEy7MfoFsDhisLNtcC7CD5p4/l/67TM3y+J4kE7zvofcY1
FYlRlqy7s2nha5LUqzSIwIswQlWPmYuiZDx1rvz7plgZS8vXNe7eTrt4tzL/Lqt9QNocQZMGxAQx
7Zk2NdxGaudfKJbm5Ot8XUn/6QK8LiTLmC/6FSRMedwCn7vvwo1VMyM778Bkq/ce02H/fcu6fmzT
TmneTRjRzID5svXDGPSCxfqGxtDU4u4JFeuSqM9p2NMCqgnhJxJmKeVZKfGIoqdfGgjKntOmRkue
248YQj6xlk3Xo84bIhMTtIcy7mNEkM1vRomho+/CpZ2DmSrzA4I9qxzpoMLvfC2y0H7n4qgsksJi
rHmsONa3qr9sqQskmpsuSixxOrhcLC7ppuswqLtJKyaUYvLFo2t9ZIB/aWq8lNmnwE8Dqy1ol2rH
4MiTuyEkO0AjoN+BwcbwMcsBuUGpmxOFo+xZnfUa58wSav+7jeFdnaRN58LDSRKRSYu0ZGOjSLmS
t5mDo+Ib+c1PdHPGElkjeLVPu7F0gZEF3KylwgXPtM2cI1CgFsJpoPDFFWKX7DnKcOs6wGDtNuiQ
rmlclcLxXYVbTaLFwm2LgzdciD1RGpykW9pvOoc++tCaqsDhastny5n0sp+leGUTzhy9qJoUiRHM
JAUN0XxC+TT0u45XsuoFxs+c7QUM/DYgm//XHRr4TnTjwD1DtBpGp6PHVlajxFVttdOxhxWtgeMm
uZ23YyOZX2EOE6q01yC9lsbpXAewV3evCtsR4yaxZnpD56Mf/2kL1LLVDOv8icoQOMnxTH3C9xmA
quoCKWRiqQk+o+UqigmAV1uY6dtazSdLAJKi5+nWaoGpUGpWLQZmI8+PBAe9yVv0apRG2/hog6Ru
W05qhHf2aYAvNnAvhHZlpZUqCLraMUh85D263jehHX6sEJc5xkJaFtuUMi7F7l4/SMARBe60dwUm
G8s62g7VDFJ5fLcMJfdVl136s6Y1IPYPd1IARmxclqLIaxym/E/vOoPJo8GU3aB7KhwgY3iybhvm
ojmTWhHeyicqUqt5EY3brSJvC4HJK7jUKszHIkdLTp4rcW+aZtAJUzG9xTBjgevCWJ4M8/tyYZEk
9N79/xAOl8Ro/Sbad7sLoZ2UMir5N/YAJmpVVq3M69Gl61cb6iaW4lcn5EBVb1vxPohWe1Dm/VCF
MVJY+ztYSYrlkSJHGFxj+zKp3hfWr1HUiSwBSpGJPkdAERTJnvjh1lJfB894WExoB3TplDRLEN3L
U9mPlu2WtBDJJW6igNli5QL0oU8GGUhkNAkTT3iMOVdTLBViWP+c4YJDlXLfQ7qXiTn+bd7Vx/ku
+3vJ6TIj1sNaSbnIT4LGFstZoEyIsU38NDnwyAInaLdhThtRDZAeWoPmja5uDCtQzVBe0Or8gEXY
n9y6vNKNiD9XKEXMa8awL0KeW+W2sLMbdS+9JUGHpx/HfQy7dmmD1GQ7e0BUrw02Fz4hpg2FstLJ
yew+T8KXWB4qk5QV9FaoNQwjh1lkWOV9BQ2fBndxUGksqxeB1R4p6j1f0SxIDmZnEAQUWJ7PS/si
PEteOfZO+PV4GkWoz+e1PflGWmWNXTCF8ftKhMdtkwFpkolyWL4dOmeMuVqTbknEjuHDKjfyMrR1
7pfBsw5rcDZj+umBFYSU8J7YYtDhcVC5w1yQ0zp6d1sCvjO+QouzKlBciT8evaqiwep89UB+Gy3D
m/BKmxIZMY4ygW8htrPdxmVyGwZwQBC6gaQSK5t2kyYQC2NClijq3fmSyQWooI6jxUSAgz0igqbh
43l3zwUdNDWMJFfIN1F0Sm+n5/uN/xxvkJR+vs+kdTEazk7FGnyGeT0rppITiTjMlp9Wpj9eXpUv
XDXs8pV9tKdGvd79tP/GyroQcIVfAtDqACr8R/W2MTiUmoNCc/XT1JKz/c65BH+gsAkGKmne+zDb
x4QplknSH9DvJxmICG7/Hj1EbGDBhe1vb90zPWinQewDtxxIHiWUkOu2I/0fD274jXvXlvSKUPeQ
0rZfJhdEdxJAKBfYkPXqL08qORAtpRXSFQG6+qNc+7kSKDMwsjtiovtAHQQZR1ArE65jJ9sVz+mL
qTR7L3yWaz5/wr2kPwfSUABc3V4FRNZj+SbP6lGy+g56Mib8js7MdNo/hLkJ/ugOC3Mc+WYG1eeP
XqXG+0k5AWD7PrRX5Xk5ND2ndmeueqH3x44ydat+6cfcQD6t389O+C0CyX1BKEETM2rPLKDGSe0W
/SZp49zMi5zykMsAjDNdTYMXJsNLcuYV8vfy4ZkYPf5aPpySAm0Oy3M4IizFQSjW54ThVofGCPvw
ueWGdcVR9sofcFDJBwsDSPxbarycYgOY0L+2zD20rpLOeZRXfnu/zrT+8XIOKQx672sI8TV3s/yI
hyp/CT777lhYZ6CfknyCzJy8b52+La9p41GxAIu9EnlhIABOxuCuR4Wo2F/CTIIHsH1jexr3eeJV
E2gQG7GlKZkVvj7FoY6sOcLcCGs9azFkU5bv55R+RPeiOGobL9h+ts4GQd795KF7jFBUlrTwx+6F
ZRWcNg39xUJiJDrCXF8/+O3mujWevk1iBajNOGL1lPPGJ93SA0U8ZHfUMPo+031LBi0BXYi1nx7m
iVmaG1KJeF21/0MCuBfR9TBHPNDiiqx2h1O/aZVrgUDzrnW59lHKYFb3Vb5wNphh9aBii+5Pfcma
rGDtK5dbPyqMWCF02vgqfzm2F0ZyN4gqaoz6CvsF/XjuXGZP4AaO2ZKB4fh77624adP2BhJoZm7/
GK+3sK5RKVkoYsBMTxtQ8ub8cEEwbaAftHLgdE3xuLZVBkHpsPTshFuTxl+9H+4G/tiYSf03MIMV
MRsaziSzd5FNgcSlScH34lkv9tG4vlxjYpEco+EiE9Xh/gTVL4KF6ADRKARhsFBntmsK0Bn6n2z4
ZdNF/YbF/OyiB6U5Zm3HigGu2VAQHMin27iuA7iL309bC6hyVfmTjPnZbr7zFmahC45Avd073mdf
c8xLfVz0YnGwB7uIbC5qPwvrtve7ez5fWz375WFTZsEPVuBKHzIFqN/sABbq5jjTeYopo1CrxeWk
inkuTvS4p9uK25OHoD9SV9InExSGSqhFe/cfK/i0ZKblz5lrz9T+jdCDLjSRf6rlfwv7XHuFq9Kt
u9ji2pyGaS69AW/NHgQBPHQSy3y9cd2DL8Zui2ZUj5NN1a5h4rFvf28yDGm3J2ga9K1V/6PzVgUs
LfQQkViN8I/IvfC35nZQABfvjSE7QQMF/ewAp0gRRswlttNxCmxmxGTBwI7Jwn8cJLLqnUx2hhJD
oK3lmeAUtWGJjbHK1jqmcV2wdORdMbKfff/Ee1qWrDcRSTmb+mNYVKzYZtv+ozIQGi61RLcJRQCp
6aAm+Lm7v82POKp5ttXux1gw8sdHgD58mpmsmhrvpVpv0NPHUcxg0mk4jwHxjfHrSxrYaM7hDOM7
NeZ4Oge3BdwnDdCCr10McRvCA+w5DSXfSwPq4OVsXmAe0/2hp9kVbPzcmYDcoLIBI43TlNHw1KMl
mrN0q2oAQVgYE5+tlqa0OMMQT05hRbNwai20vrQmeXwlkA54LKi5HyWbmI3R8YHbKS2PdF8eGoyy
9vrqRPMm52EkDXsQxcwsGteUwjTXueYpfF4BIjMXd3QX6n4EpviLFPdS+OPiuXp/nvFjkiqkves5
aGJBPdgEdOaJ6wzGiBakJac7lNVxqzd/lLiT02TE2XM7Hv3p3e5uuiY74flgCS4DD8nqEYqb5Kp8
nM73qgW2MXT7IcYx5Eg8xSqOyOWcQ0xN5hm3qmNdCLu6Sy21X9b/kMWzZm2Oj99HhuHtvo+Attn/
exIAiKwZS6P7dgbSn6fEFiMBO7cEv5skP8f2+wioFhMzMexUdJUg/d7IqVkcatqkE/7+lCEspPvm
7Z3GlZ7xpxhPEJcd7/GiZVojrDp/XrytdgYIO0ea8BnZwSsC3pZEzEqGC0sBIx4IPRLTdsEYlEsU
KDyDalkLOs832LHOk8eLPYCUIpyzlrz7G6nro7hqK7UhLkcXrjGkH1yzWYWV2CCYeZ3HRoIAY3jU
c1pNea+s1BeLSdtdm4KRIQQ5A4P9GCoiEDp4tKBgpTDl6PDQD0v9s53SPwxLWkE8h3sPB8JOSPLt
lzAbvrK0G4tJ+svN3IL5gMjM8rE/CZk7GXaEHhG7N4tlc2HJQmfGMN+4khFR0JVQrrfYhszq9KAO
A67tZyrx0S5+Cwpl0IRFMmqfSRGkNnfDxz8n+Cn7IF8etH3KGMgw0bK0isaKjWnOOwX9KoULhZ2o
KZkWphOvrU5z2M2hSGwWoOBiR55k21NzeiqIdouV1Aw+xVLvrMUWdKzl/DWcF1WV/CcHP3qZobOU
yau/bu+zR87yOCfzUPujzVInVLRxkpD9mD5kNVwmeqdJofd0Uml5vacgR99qXP6x6FuxT/VnrYjx
vorMkGN9PrLdCHiUdxoQUty/noyVk9tx8KnHCjYlpVeqO3dT0v9XezpjcpanTzg/ESwS0Ao3CyRy
wCvOW1UmNeU+Te4CMfJoVmv72QEjxFaLDmb/RAejzpLGntd+9qZDdf/LxIGh1T0yjbdx7pEEjltI
yzufOkmFHQw1gnFAAFSMxW5VL88N3cuurDxkLgofBtYJR3UjQAUmz0vuS2Y5S5r6AF7xbINoojIJ
L9rxehT2K1cWoZO6Zp9+yZEr7Ddq+4Bj7uRZ9gcJVd0oDahmR4W4Apws0JTGOsVO+mT0peC4BFHN
6E6QI/PJCRajr4V2nmDVUN3r9d6neF9sQ6tk3GZVga4hKkwQDVDZH0LaL60dLJvb/voL/Wkal8pe
/LtW50Jdvn3fbgVnPD8MZF8Z3aKG3AAJGvrjevJQZBPYj7fT1kASoV8f20qro48Imd9NclDZvXqa
URIgzBg82r1h81R9r+mtwNJro6i4Iiddo7if7mnQg0+ale0S3hqTeQkewXiy6NYUT/HNbh+GFn8t
BN32+VNuVhmIsYMqRypJOcMp2XHMtakYO/xsXi3zlFhSqOTdnvoqX6SCeaRHwHry2YGEwaa1FmLY
/u2YFvxBEnaz5ngRYoRXfeF41lRi7uZB4/H3Ex55W+B05oVNgFKfXL28KTVeH6hvo/9Ij0B7+kuu
aPoqH0p8NYe7SMpeqE7e5F7WdCI1QHiLD3n29lAEj1Cs6BfheoNWPgbxSc2aZLCqu3/XFLoCtNsh
obCmR01Ll5cqBXVbj/rIs9bVao8xO3TR5ClpQK5XL2K4LbSW43QTe3UmI+BamnOjkqUwib1VGT8D
JEp8CeAtNqkT9UgponPM9auH4A5bGG+fQNlWoIIAEKxJVmoA9LX6GPh7dUXsxGrqv4H14vaktDPE
3L6tbcowvCQEsvXaYQfnyagJqxW8f1CCJhWGs8mDsXjX5FnhCid2LX1BQN4lTyFY4G5oDQU9bPZn
HogoeAh2onJ7ultblfHwkhsnQfG5BIZzhspJLeCTsdb9iz0SUczDqdnKBad51U2HMCiybUq4py70
nTOaVBn57JVMni19/Z/8TosJixSAlUksPae+Lanv+bXXCy0pQHO7Me8eLfAXbjOjOmbjVexU8Jhf
8K6ahtG60AC7TWldM3HtWhSf77PhWeE2IDltbqS/l2rOFqmo8Sbxegva51IG5ImcmaaYBbV0QmJb
r3ll6y9icfcCLZtQi37trD9QbxD2DCGb0+Uv1HAr17FkTR01FYxWusT9B+Y9AV232wI38oS9PJDK
1E96P4oDfLKZOA2z/9q4Rctibz3bYXORM9jwKRB6EasffQM3zuQ6ujknB9aBxWZayYfervvtIOSh
A+Z5Rb9yztyGY4uXOeKZHI2yracyHxnVgZu+6qX0/DX1OJVSvD8GfaxYr5qQWYvwTGyQcHxpJV4W
hU3L+n1g8YZPNQPkJRLqfms0R3fKwqp2Ubv8Ptn7Kb+b/8jyCAvUeS++s1sb4e+TnqCNL+6e0zEQ
3kAmyGZxDiB+GVgBqF80lb83nT69wxUPH4PbDTnBOX7ikHJnHyAFNobCOwmKLtUa7zZKsH4XBnnl
qAOW6sSeWr24ZEJPoNrt9cCNe+zBH36W7zpXHDi5mHVw5MqryEQSARGPT2qhES+OXHLlnhsXgiMt
LtbHMxO3qYp41zJ4d0KegrH1lppHEQvCsKfvR6OlabBaPN4PsP4eTm6VHPMkDO7unl+ohQAxFQrf
FtsiamjphNzztTSs5HRcSfrxiW85PeYO7QJFaWs8hNCgvT2jJPLIMW22911PF45pUqk3dr5l1Rrj
hS5LRFtbndx2dirkc80H74vDRZOjyYGwZTgAiRVkiTMi3KxpGUANDWuaW5j8/Gih5NxvZQcKg3/q
60RzESPViscGqRnbqdMedp/WzoWyWonUCUyMUePQ1sZx5i/OvOWEaPmWk+nch3XlgZDF+EJs1ev7
CCztekO/l+JTYDuHU93OMWWeW3XMm0dzMP7kaMerSgk5ZnrIpp4GA6UkuGQwJzc8m5Tc9CP9pIps
04qPz7hF8BdtOOzc+7m8Vpay7PP/253EYg6Ew7g23XsdeiwP7ebaCtbfO7+EVOf/HCWjv3cHKxQB
a0g+TKiazw3T2ak/u9C3bi+PaT2f4jNI8xbdrI6pAQVgxDzY053RrWRAAvBidpDfLVeyw45hmmMm
ZK3hLq+sPYg8ft+PUg8fDvoaRhgvsgjcWmtY5lEeqbIwwJ93y9NB94pMe+NenZdBVJb7RrPiyeEZ
mSlRyAGdAD+FvQzFwboUqDQFHhiGe28I+TcVNfz8SYJKOopU5E6R4uc9tkRN8Y/BA8Tn6up9FCNj
p4F8fnCD9ogyyVAXQbnRle22OnOOsqQk6oB22Hp87HxjD+zxkEFeUndfURGGkjGHPoCidt4/UT63
LKSGGQ5RvfNy7Zaxuyad95aqmnfWq97Ss1vGXIRo8a2jjfiI63Vur5AMFJ26jIX0BoCJGw5Ih+2W
+eZX0amjk+Y2fKejzZ+XJ9aKD0SrOrjLYPfRTLVVq1o0jw0M9WDZ7kR43gj3YzwJgaeGuwkbH+8C
nQ32Fe1pITuJQ9HO0tLGSLdFuJeYupTx9hXdf96CQrVOpSzYHmPRmlTzCZ/vX8RNUHazsbW5En9p
ZHOSEAi1vbUfvIeoXUedbyQnSKkfmtPusNX2PkDS+XHrTdeOtISqwkkByDLBbAbgZzElkwyvDmfw
9HatojRPGFrrZKAqEZ2tK6T8W9oeTXrkAZJdj7IE5IyvfVZYrG3NENGy0s08EjaPpvt6zJF1pez1
JF+Gv6E81xQfMz2cM+pyh6oCrmnLM2v4Q9R6tiY7FEHg5s/488EGYKX0tXs49q2HwGZwtXqI4ewq
1mbbxc3/NUEs3ukskbRapJPlvWrsze/F/35Y1BW8rwXByvjJ44h662N0N2WFmq+1+CTekJnNcjQ2
TK39hxDKbSDOb0DF03w2Nff7469UlTaq+Cw0KZtFNduF/1WtRe/0lGhND7nZiDWjdDusqQJPtQew
shFx1eRnljGgwz03dNea3UVGMGeNhE4dhOqtGBj15NNYjl5ZrPu0Xj+TC1QuHf2B0hdEJ+dNVOfJ
Za+YVHy9VXgDsfdDylwjo6SEi8MK9KJgJ0/hgsvdb9h7Px68RDVsAPKAEELmVcctxl5ii5HTjCZy
qmfn3WG78r9bQN34GdiVywJJoKeiDwR+jEbirhpFZQ0LvMdJNe2rBTxxtPQxCTqhwhM3OYp7kwGq
QeuxILU1fnxuQEG6lxthGIB3X5d2YrGTic3tDzPpQASJnoND5nVY3kA5rvfBm8zk94xzjoKbVZ+9
lJmM7cnOGHlx5M3Unyu6ShhSkU6IARUVEbaEB6aVzCKHSTnSks3QiTDORiz+BA5T6Uwkt4l/KVq9
QHKIqkeJM9/cwXnNmVHT9Rms5145Km41lNPvRj7gm+1yEuVRWWoMEN2ywctyEXOwQlu2uepem3Hy
AgSrwlLOjeA9TM4Cg+fRsRtbTtnP2DHTBMk04e8g54PYenBkMj45NS/62GmLQroIE4MJDIlJNf/q
JFvb1xpkdFPDEat73KyWc82J3UB3H5Z2XQ6HKJQlcssC5ihUcK2wH0fkngCaHVRZgIcWhu1g8Elt
qTVlJKTL3xcNBo8uMxCw5zZ62WTy8aL6YpJtGSKFcFZau0EnjIPx3jMmKHfF00/qFaSn7oyvkTnC
aPOZWOOJi4GUnl3WDtCHwD6+g+npZnM7HzeGKVUHbNAPX/Qh3HlKmEgvo2Vvxqe2g0G39YRikCrr
tG6Nd+PQ/F/dEbv3IVLMzoa7gLTaCUQB6oMrvTyNh3a0vyGpSfUyqhcknMhC3vcfecdZZJ7qsSnR
2aSuCXrbsS7iQ65+zjl4QC7NaiHf6PAYCOvpe1txMMVrXQap6hN5JEjJM9ed9wZQzQqDeILxFU6g
Fyn1KF1MJCASVIBSXvYRuULy3kSaMICvYes0r3x+HoEsvYI0ImxRdRV7OnJHIfIkrDNXT4mTGdQG
aBV4pfe7oTHX1VVt+kSIqbY9oji81zRw9VImilAPwjZvN9giWAHTNoVNd5g68XHgEcFh9SAv40BH
CcSv32vsxUDiGKs6w1ws6wnGxRFrlpC4dGpaNYNz32tuGwDg7Ptq2CImAjz87E6aq9/7l/SM6x8H
sVb3DyjD+GkY8Ia5r4os/e3ViNjTNe7O3DDC6nZKmqBvz/6Wy4wujBoyCcORoTeKmPGUQiOI/LIQ
lrSUzCJcFuLEjA9yYdNF1ZbwupiqFgVDEayletuezL9utMxHgr8jyxK2tD8VOwyrKgnA3xBhFxS9
xnNH3auRJ2gYxrFM5C6cFxtWbCrPemPf51jEH/bvUBi2G6AzDveFPyOmEZaU4ueSONvdDG9h3sJa
MOMLLC5nRmd3aO1PgjqBOmyWXgtkUxhfnnQM4s52e3L883Gu+5AVw2bta8L4LGHONfm4mrTUGMHY
aRC7RRUCq/C6+2jhDGB6sAafojzD7xO7MXNjiS35OErxhhKpBYdSmvwX3QiEOEgLQUm9PGkHOu0t
odfUlBJEhR7jgk3Ri6P26OOxeJtInWCnoTM9PXrS8gWt4o4VZ40Q0eko1YGU90GBZULdlUQj2X70
z52JD6jj0kKlv9Hq7sLEDm8NHAbr5un0BoaqSV86+qZV35s04GRji8vAbRnd3XREgkC72ZYplNPB
s7SeRTs2H5V/x1vv1LZ+sLeDIr1coau54HKgqoOoPRh6KwOgM+7/rZ06xXjLe2qlnXHRsZnp/PQE
Rask/lm2AexTNcAPM6rDoRoNGljgCQwiCrdzjJk9kJxd7P7T1ruct2IAoKLdOH04N0+YHf3A4CzW
o4tee9AYBAfT2Fkq/6ferB4CplWjJuy7WHR2b6TfmNzblydZ4wz7XabyJR8ccKn2kKvKZrC4L01Q
3WuC4FVcEYsPdK36kNK1C/NEWFLeyS+UblqtMeqHdVWCx5iPQctF89O/cVm86C3rRMTNP3zNEZOT
Q4Nb9G4tzXtmLCR04qImGicqjn+FpDIZ9yEQVzUdY42oFh9IIdX4pDhViJ6iERHlBV4zLp2CEUGg
ggWtULMljcLvD7PvLZ8iOGSq/yXKtDFzGvxriu6t3oOug3KvsSG/m+mSr8McL3cmyRuZSPKNXMWR
inACpuYVuyw1pbu00XbaUoFCVBMNUCMWnbihR5B/KD+S40HPKDfzXUhvhg6OSknLWlHnMWZl8oX8
lOlOQcawU+Lm7w3cMTg8HeRL6rJDB+Y2NT2d+BJo8GJHt/JrynSBTq80gx9g0Gq0w+Q50zjQLvhZ
ckM84DiD+LOgfNsjf1+zbeXx94VtUdSF5+mUfp7DMDerPAug3i9TEcIx1oVKVLEQnrdi93f2pxJ1
HgEVLa/I86MCpUPzdn+R36iyLWXbpHrbEituFDLib9SzQKqJdSOmkb9hUKGMrVzXHLPYwloxwXgP
hd31vt7+2bkd0Ap630QvtG0eS/I9pNuAwVFdDYMN0/AyzdUXUSXNUD6Hj4a0aqs3Ev8erv8VvAsA
RD6h4lX1xedgVV6YYBIgWqQuylFk1S6wnUKlMiousBN42EvHcAfLWP/zv7rk2foT5qs3wBkEzYCJ
BeTYmZ7U8QjxoJWpcEEvezQ+ricCZyVPVZJLMCC1qncBojlvNm3yiSDxZARFqvTHB7e4jtZhCB/N
kTNrkGPyEDbVeQoXlyFBGHybu4UX/1r9rGJEdWT30O16H4zFYVedSK9RMMQKm4zG0ERwaAKkzkoa
m4Vqh6jWpc3/QJJpPuHllX7goTipkwU72DsSqcy/LIqcb+SMkk5WSWRUR2ujbqiiWZTAZqSI0RHe
j7036FcSVQwk6KNa5ptYbN7dmZxI8zYPUq8jRJd0vCJ/FB/FhaU9KjVUldwgWBTidlkJwPIsLnDV
WCPwOEIBUwx8wl+YFe+seCc/Z842P24IT9e1Q4Nc77nyBqH2sJ15HuKAFvmkhxboLdZD9m842kvw
TKRGi3EKJhInNlKVmBugjLAOWadvsyHbKsQULnN0PsOI55DP7siLjc3ttcDEeUZHRJI0a/i43ocD
eVhLQcpe/dTBEUmJUbWpPkmdKPu6hmYP5zXPHE1WWl25auGOob7AdZ5AP6agyONoufwskA1tBC1a
F/JMOhb83UE4DIBLYQAR5KaxAFyhza4Z5ryINc6S0g28z2fHtWDpp0jRcxe7o41pB4+IWclq3bPu
TWsP2fXysMVbN7K6OlgiHbcniPU8eN4tbroiR++JuI9Lh2oxsoZYGg/0zl0xSnDFUMBkEjKmDkkr
nFEzxMVQPhjnWn+Fv9WfD9jkChv4qUeBUmWGd9nZ0wrU5fTXQlYAgt8KsgfaWgiVk8UXDvraRw78
Ngndvwprs64dAYNner2551dhR131bEvFGjM7hg9G7LrLvNhgvDOz2989hfNUzCu2hMSQgeWcukOh
UZG2A7mgWaqTof0z/51o4+jZupqwfEZwrTxJG8nQnE57Pz/nPrQ5rXgLVMwmBSgW927g4xpZyVlH
kbLkUskzDw4CMBjLREhBag3RFr/ApQv+7dQmQsv/n4oPOAh25vEUJiCCUdE+1nxmK+zIxCaN0fWR
UQIKN7H2ydMSSwDS6Hh93SQH5YppaVmSB3G7gkBSyEVvM37WRo+yy12fkmqzK4mF2ZSeXmHcIMz/
AiQtDXyTDDZBepYcF6SOcpwx+6kxW3f2B3yc9oG0qUWH06J+RnsSy1AnpVF0NpPCFuD/i1MsuMcN
WwAbmoV+sn2+r8JZ/081uDYHN+LtYlxQeTzyYTBn1hHluLB7u4gmSRKJOjY2Iogxng0PG+6uQA8I
xgyraPeenwhfjW9+k9zJ2LQWQDvimlD+19htYXToWcK50Rj7EoG3iOVCizMHAGSt9b1Ap/dZMdeK
h/zWcBG/hv6HQOcXzPOpfpk+a0b8HzXXafWlj9CkTRT8r0YYyrTprUZjxtkZkk2QD5/XMvRKytn/
nMH3hzkSrwOVejPZk3jw0/gv7TCLVW9W6ijxeiVhtS5pvOi6AivcwWlTxtYGsx2scHSwoQ+Vb0hq
0lZYXvur9TBdrETGgulth2BnIev6sy2OC3iEk4Xu/j5Glte3OdXCuleqLDouDyt/AeItoYAc3GC4
odwDhKfA7Nf3U8BPjH0BQRAaIiNcLmghERxJMzrHcw/sN8Clw3WRxwH8ITPJra6af8Y22CQzkm8C
H54Mjq90qlq6s8cSYLUJe6yTYwraPaoEqQ24oYI9LLTDTQ45SGtw/fI+b84VwfD32kFq05UDIESG
53HM0EiH4mzgibxqjWkLdJ/mtwlWdhOkdTVKZUgzwkjWx1ZnioeHhKeTfUN/bNo+aHwqXH0dLy4E
VsNhhvdY1xyzSgeNkTaxqMyBMtDoVn+/PnRln6jj9TGFNkKi50+aBOPIAeAXgBgdJtmPtibjdNmv
20OOSSJlI+0GiJDNlSFejT2OVNIZ6NPQqNU+YMoS4kdm6s0EX6URSFoqvp1hXcaHOJYcQp/jZzxo
K8e4EfIe/kQ60jJnMfRfZGnMtRI/ZMztvLD0Rj5XeQVkaHfEpNLnV8LauW3fdjLgIflWP40XqGfR
GnRHj3E+fDunx+nkiBVBwLZ9P0jtqs/go2FUoY0V9rpEJKhbxuRInazFlneE6Uw8ldbuF5asbDGg
OKTTRlqVwfzUmxbbbIO6QJj70uhpHUlA/xBfGZZhTQCMoQ3IUuyGC0SLNBkWZGrnamreCxLQrf+S
iX+EXTpqMATj1Xhfqwe/D1woJi+e4NGHcMwzViEilN4WBI+7c3gz9DxLl+H1qDnwExxsOPTbyNVT
led5aCRc2ZRjUf5dfwx5axhW8elO8DVDE5FSnu+kV519K7mS+j5dvnSsTQIQ1azJKT87YhoJPXKl
O7E3bBNLyG5NaSE5N1l85lEoBYUGfyc4dJ1vfHGBJLamDAV5biWD6wxLCbuOD3Z6lQ+Gkj1ep8W5
kZ64P0b2aITRlawOgom9k91WzWvXxIcgpYA//adBJg/9f+w/mWcE3GQPXp3uwrVgc0sJvVxI1Cqm
WNxsOMgHUbOQaBhpVVgwcz8pffUyZpTtaX6vDddd+3w7qmS/ig1O+D4EB4MnIbSO1XzpjcsICKbj
GeMhp9cbKyDg5LOhIka4vzW0C/Td7FZl2fLpt1Or0Fj355nmq1tWsaEkelYXvVPUphZvTn7Bwuee
wmab9csqdSaVpZ4tnH7dq8TcSyfpK/LfpqKulqWf7CAC8Tk//nCIHJ40cnbLG/7qA7unKyg9TXPw
t86azF6P+5gnf7CtX7asuHcy/bxc+goh7f90AMOwCE9uSXea7VqyzdaJk3R5evn2AdevqNPUMLMb
aURe9X+h7/hxZ2CBYmcdP2bAVqE5IzpNergPAQyC7SnVEOUOXxFgKZPdxUu4CVPZaOsVPTQ/yomN
vOpeVoL7HKFHuG7Ey/ZU7xfTNhuxMxfOpT9DaSco6KVbYbJKJZ+ylje0mHiEqgmEKMxjhpgLbh4/
a90MKxhxFuUo4KTfxau/+7/EGP2cJFCmOCg+1i6UFjZnDwhLcn3I7ysn6vuY57EvQ08G930c9IVs
z01TevUvTaPB2IOohMOGJnIYxMx99ebULXVTCwCHhlPcL2rz2mYHhhHhMgZKo633MXfmt5TnmhkW
6Bd9I8l/l12wcFho0WVM1G8qYOpe7gTaZ+/yI2y4YrMDQJbJkge7862jeJsSYPM75fTuKg6jwAOw
ngukRqGg7Lz3IPIuWyuU7wJY+msZ1kkLmObZ/4DbAdGYSyPQY2VozAkLoCbCEZi9ug3aDoFC6N7M
OzP0L2aKZvGTMU8Y3hX5qkx9nRq3P4nwcdFSJZMYFXOOHc8F2QtAhpMgpHUAcb15qwDA61C95uFF
BvJG6ikw3U/YV9uUf8hM3U7e6R3W4mvHmQHpmmY/nwc8gYDq1hSAvSIVgF/Dqvq5Oz0aHOkjF0BJ
DrSBm5bKJw47qFUXuIcRWGe1BxGf1WgktVy9Yyh+Y4dWa5nsBCnlCiBl3+drf3YtTO/GKzP7TWEE
YdQZcsQd+t+H1lByWqwyyV1XmHgZf779qkd6T+1+oFuQ2Nu06+bprQdIHXQEsKz8Dt66++npdia4
O0+HKNo7augnSglhT4awtQyBP43qiW5CJ37tfEkPcfe/X3J+8fFuplTcs//QzHeiKKiDaY1Ycolg
0d9WYCt8m31mxe/aN51oPF90pp1WT6RpIYd/knVKWy8tEYGkOSPlaQ1YOvco5hOYK0/RJlxNEL2T
VFk1eV86c3IX/Tj05z0djmWE8/vV52j6C+kWpqWFLfsArj6TJ5+XskLRh4SeYQckHhSSlAk/WC/d
XZyvSCxFAipcMlbPD27mOfSZHhh5E97cIVgztAk5jvpRefhjhadeLGvQQnwI8GvmLBKsqU4ODQUv
Ygm4e5F+ILGujOt8GzWOzOp4hbdmY21Q72MvsOj+D3MOn4IYuG61n09s8Y8BS6OMOOuwsvZwq0ww
Cq7RE0+I1Q3/e5RvLvDunbAvD+w1iEWCUc5E6K3tn1W1IZ/ecW1d8C+k7CBCXwynbQyJNTwNaiRf
qHWWHfP7qkdl9RfrQzuPEC0Ha8ZAdDa+UgWQe7O8kHcgY1nZqNvGP0/qOhdMO/mjpkDnJgYTofo5
bZR5kCh9GM7/JLIHqSw/g+BP9uG1t59RBDqHzgIxitmVpcEjW7A8hGliiijGD1v1V6yDmJxtuqKE
xc0hYrZqazd6PESPvDPcv+u8xmspe4o6QDCqZSmgLTH5gUhT90CqXw9zlsnCmXmM9+WMXmxtUM5c
QG8d82O6rhzCt6Qd4i25d9tvAbtvt1ZLyNg/Z62Wlf2gQEeJWwQNGXuSzhdFCXVhcDBubI/iQi3r
RPMoTkxVZhBlEdbxXZVvzCwcemqQNV2SSB1NqzfZpCT+ZSok3oqHBhUBKcKYpJirdeyPDAtuHgox
pkeuH3E9wcz9iVtw4U6ETths8Bs/sRRFIMY2qApTjpYF8Hq6UZOJe0VjnhD8Q+AfrZD3nn1fzFca
VrIGV8k23yulx+ePXpbkuiJ7sZGiUfLgbW2wYxqRTyBfgYQuCrEWhDHpqZkYT5i6LeATGG+kk1Rc
hL/NWoXv2cWT5CtOTdXbRlQO8qT2TRUp1BKo1S0Ji/p/px9QXtDRMYCuP07mZ9c/AxXfnEzwbIR9
QwS6dxyECrLDIkkwl6yL/D2rWtlPiLgExmOrleGRij4Df/i4yJ6zOe0f5IdRcQdu0ZFTFVP1KJBy
R9RznGnwhubze0VhGZDjIFk5Nz8eibbcHB1GIZofstvm5NFZheH/PoaUl6h8Fjd4pWMTXmDivetn
eBm41E7qzbNqAmKLu/nSWsBmkEzXEn4Z7zGtIyJcBPtXe7chJp8lhcJfyCVd630E6J/KwuyD08Ew
6LhkBeVZDrryyXUjVBDSxXsJQIBuZ0ng9TYLossMyUp90ji2Fn6OlLs50n6Ogg+xBR28+9ueYphY
Zq23yZNBCcmpyF9beOAaic/G+KvXNPOZVkv/cDRqLSSE08gdTHCwIK4xLSGqL9L1iuXV7942eY3m
Ycj2aydigKzfRg9ylL5xluyfGjSZKx0Y0Bp8OkV1SXdrEr1J7pDq40lDzH91SMtvy7mkc2aqDf6G
jMUfRo3QpDqfMS8RCMwhZDu3gLjejFTaLDaYpCWVAdZl8QtlrriOGAf+HL7JJ1Eg6NsmqK1r6mAW
tRdFfJR7Xur16RbL9GOxWZzPdIRod+2fvjV78RNC9+Nk0QMRnXSMC2dULJX3/UoZm/84X6p6iEMw
DLarJ4cmkvze0h97mcpw+B/aa4xcvSMwTg5ndSaoNRy4BVYTBncJe86Oh5OnD+rBrwYCoq3xmI7u
SQAmQ/1M/PyjMkudEtl3P1LdFprIV3cvX+EbfYUIwZYS2J4R3+OLXfIszzk+SKk4l0jq1ywoNvkR
SuF981mrVT24Ow0aa4ytI0z23O+Hb6gm7knhIw8fydh60ihcoLmcsMyb+chekhf/r+s/9Kx7iLSN
6+u3waJexRFR+VyEBrUMTe3UTzAVLzTOs1/Is6Kd25+E0/mWQrFDF0z03FOjtsUIXDXMHAPRvoFe
58b2iudUS4UgZfxfUOM8j4vmJLmlnS5XMA+MurkedNvo95m6bGPCB6rf+7tey0e1/zCLeJm8aHWl
wNizXjQ9/ADbw6GHat4qgLSdAQLGAdvhsessGrk0wzDZSUx1TIU9VJ2D3ukSPyG3b+8wDXGrYHGK
dY0mUsdH9UF5BSSfMcYRbmJG1b5LbvE66tp0gyQPAoDMyivCIdgO6h8ClGH7QWHgvAoVOMwvysRy
G4FVr6rOr3f+5F3nWobE5YgTOxakxxp44dR1+XKtNa9p+JvMvKLZ8QWYeAuSDfc0r5U+qhpQkf/P
R/GPFUOMxH1cz3c9QYBV8SQTHAYbGlo8meVsQ+h/6kxUunfTIH8IOluNKK2vm15Gu4Qihj8k6F2f
LhdmOV297F8SupBlzwJkbRR/NBYbJg+uX+Jg8D0KaufasEA9YzfZ7Di4xPvT/vTsXZDkaVTfxfXO
VvKij2bjAOTrx6CNZOlIPL0F4c6P6Ro7/imlDNIVJLbLXk6TfjBZHCheDQBaK+hYtUslsamxFRPm
zmy6ncFKCLxHKapNkPnX00vuH/4zV9OjMwL+Q1MamDjjrppY+D/YRW8fTZ21ys51CiI7Sy+nRBT3
V/FgMq/wDXqvy05MmohIBdHP6s5qDWMf0RWHWc8YRWEBDpoS9tG1bR6m3FcJoA8TdNfF1s4rlkcK
42EVOSPGOhRqe8sifWEihdnFnQTldTvBpbKWlIEZIhNAseg+T/Mdut8uZR9mG5W3Vg+cUHEW1WtB
VnyQzDzXnbVkXzyxLNxZsGInCeKkhw5RdiF+SmCsZXS34QHEXMFVOG8z+wgFGf0vlmsQXZhfswjO
9sROAwI2+U4e1WytORM8eH3s7eezrxUp08UlHbak89A0V7qckwXthBM7WOSLbIejbfDq8e2jrQpe
OSX6HcxP4UqgESan9iVCShN3m+GetPWdL8kf5Iob5q5c8JIPVTESnViZUAOAG+MLhk9Wu3z3o3TJ
NCXGst1eIorNZZE90XOlHgJ7Dow9LRuZycHRJUKAFux17mPES2Qr8oRL7ARaYPhOAt9trL7XufcO
WU7l37H3mNPpez03q0SzX17eESoJSqDhHcUTyJ0OI00+pTqGm7g8sj+BDEdrezhVNgaseCUhMdDt
vOlvLu9VrxMeOdY3gJ1XDuqFMp/YzROLiVx2pC0xb7QtGD/KZLXpi926SsGGv175uBC362GiVffB
IbeUSZ9ILzaAWQpgEw9H6ytwUR+e0YET+Jh94+xnRazwxEB7sHDSzgxrUC/2sVIyTX+lOdrYV7KW
Lj/yTiUm1mPMZWthcowjPKKzvbYuL/lGoJiYHOVdzD5p0pSSVmJTGCqIc+79Pl6EI1m3Prl95EZY
sseyvqWZCxHaRS25aq1tuq0kb2Dx/LrR0kVlHUyDPXvOTOW0vHVgCYc7WNZFztCCPPpnwNy/DP/X
zmCkRbEkA+GZD5UuuaMrjnNOVEgGuJ8HvXZIWTIm+IMuRn5QwjkRoqcmXKxl5njJCO2VXDnmi5J6
+X/GWboaeCD/GTtYOk+bH6uxpPtaco2D+lbtzY6zbl+WGAy8e4PeAmOvyGXbPvNXqoGfxePnJn6i
LbUzqO4PwrgkSqGWPDQwyyU8GPoi1um5sfN3my3UVYf0eylp6pKR+o0KUDeT//pZ/I7vpYEZBfh/
122xMYpucrpmbuvOETB8fxCbZg5ko+CVSB5EytUBKfXSefcA3n63SGc6DyzqmEjM0GQgi2LlZCQw
6SGabkHXKKYk9aFIrdAv7t1NlHNYGn43nnu3tJs3BijgW2r5CK/HC+gnmnjtju8vbdo5twfCct9R
LORm6Qct5W06E9NU4790X8EACNLGl398bpfoKQEAFxXsrCFSvwgOFAadQ91+I2cJIon+YG229bKA
aICrg1hNpyS3dIOvc3aO0gHB3YnzzVh2KWacfdZeQHgrGubofGFbbsepxkZnx/9GM1dkKBB9mz5z
zrin/xX6wfwfyUFYHT+bZNzyi+4bIt+RKPn95nXv6ucu6KvsMHayRM9cH99ViMQPVZWZvUi809Qw
ZR/5A4fSivrvgrs5VTuH5L4bWRMgXPsMU+eycm/h2G7uBoHkYa+hffCllXYW98nV37wpoDWjWf3b
j0EGlT36ZvNfTVw23diZ79N1boXXYGmpl8dhYDajE3RuDdhxstD402Us+AFOQvLE9W3FnqaugRhK
VXveypdCfBeay4hblZDvZaLDMcFk7hjkYx4lO653aznhIDAkcQCq+Vm6jviyUjZdXXhUp9q4+YMc
dnTcLTMknedO0E8Iz87ZANKFVfAOFjX2AmXzHslrJMgZDfxUQ1BaCO9H2jg/l7DLZz9+vxfWZXux
/ZJ7BpzfVeHmj6FB7oT3D+P0QSEb4BYn0lty8O9JtxJuNCzv45WtPj6jvDMrZPP6XnL7oEMtxtRn
kWHYv6ChA9m/MXKWg7furWO0IO8kIkyipStwP/cV/iBUlJmbsDQZ2UQTzzHuIZQ4YnzXZZnYzXX6
YhCVdEYAcdfOjsxKrxPpWVgejwTNMFW2lOtePzdmaUpws9xTrfqGG1Pcuq0lAJhgKDvQTdkAFNG7
uGbys8P6R/eySw3MC2FIA1gfEyFaBJth6DmuRDo7DFhVLHj/9Og4p5i0pYLmSiGl3lVNYnuT/2SK
lEe8FOiGxiZ7Id44HYpE2AuWfx44EF3rSlwtVvmjEdq9SM3qWSz6kfAxgLkH9iLow3pVRzFobeB4
TOWOB6Q3d9s1ozn/j3jVeSCQY0x9ww5dxJuHww73pU8ENPHyj7zrm4QWCVRNxmF1+3272MgzZ4gb
WL46vVe2oKhaWRF2ICLs/x/HhUQOmT4LiGTjGDfOKB5aBcoXSTQKFKGSFYYcm9O6F8+vLzrX3Xdk
AKakA+5z89uX1EuvreNNgoKfLb7/Tfn18guRDuMo6RLnPl74N+5xQRzQfPAU0sqYoqZ7aujCdq5f
KHjNqMpd8ng+yX5/1Vv0RcAv+dGb5fz5f1OsPBL+pM0WuaYPKBDqx1mMCtFgMoQKxkV+1n5Wn776
3lsqTU8WqXGwc8bLnP2/gENy/0HyDIRcLNtt8Mu33M9zJnKqc2ySZHMFcHSdvC1FgKJR4myXmjNg
+ZEho+GZvjnuLQ2GoUBTxRnp7pmXfTMZv56L793P5uBvpo/vf3tLtYlxYyLqKbW9R2w7Xo/dtaDg
8EfvQCIV3Kg4naESMh2/XqkSyIPFQhOeu8VLPhtY1KEM+Ur10s9fqpug0s0IlpTQfDSzLtHWttfF
m/k1fOvizjrrs0xsICfBOvt60LrVZdPcdFdZ3ozpR1WTSbnJF93q2I9gPdz1QSXmKufPjDNCyfVo
Ed7o+9aCXwM73Q+3JI8CVpDZmzvkZzAXDOCVIGQ+U75vYCL5xRQ0m/MEt19JZQVQ1D89vQCkB1re
Zws06QSyepJZOjfo8v8jj632w9dPi2AG/jAfsPUezn4yfBisOuZwfUMyzixhzgEN79cfu9Lhktpx
DXvsxA18/w9cJvyCpwms26gYOf6LQ/AHm4SsAlIQW0GAFHW7o1gBoM6jwyZLtIJCUxCuRabX77+T
9Tpew/GRd/g6H/TLiSF7yT00AErbulPpS7DJVYxX836AteoiGguOeMVXSCKhioeBGzAdtb80g0pl
glWG0xAAxkZ/G68WDFA3y93oxn1baEDlDvmhT5E1cxDBqfEwbSK7FQh9Jwv4w6NeYvdMXtURyEIZ
vnAfVPaPHE0X4OFie9wfrfgvd7/4nfk70jgRFHDFiSCFJyUQxRVmvOK2KUdDwdJwcJ93Sm93zWSy
DWd9dWG+NjdPbQqfJmjqCC4V1dSYk1Jh+iv6hqdr+5z7Efj3ITTHFJvkAXqVGEMlAK1pNKsaFxTS
P1hs+xlWUYDsvc3HFxfaJOuXd3zUrgpeIuQKSziOsi5scbip7WqxeqJGzQCMTXoEI8fHmO8OmhQv
Nr0shXehGOkC5ZSr0VXfxUdKBR8YMI2qmKRx/jgr9o2/F8W2Yvds6yO5MfB0lAKlGxJh8ROzsxyQ
gg1vUYYrre/FUn2AHS50UIYQ8I65vAlUDMqMalPx3M+LCn91XftVDnRV67yG3O5cw6cN9NDczLrP
9hQvcZKRcXIU3qSstEf9p73oMhOGU5o9J4Jr1gvHQnTcdfZKWQaOFcYX/RFLLwi4QKU/2D6w1dQB
rPghjQb6JARQvCmH1MujqZl5ty1QBBvxGGgobZq0k7iskmBj6oa9uO90X2O/jWJNCl/XuJu4tbng
qeF3lt1cXHqeACnvm/fEDEx0UyuIp+c4MNDg2M4ezlIEwz3FROuUGti2McGrjy/uA/xbCxmL+dYb
GYYh+gn7oWB2W7Ibj9MLjPEJyztJPo23ex2nZ6NQVqwjYf9QsLLVzlosbaB9qRmhrzcsdbcnedtx
J61wHeUh537d6ckhIiSpd6s4oqlRCxQMlBWNQ5ZGkzrVyvNiSyXCP1eroOw7kf273z/2ZaxmrOVy
KJXQ/DtcRhtTUaQW0pI8o9n63shgqJ9kLYC0c/aKuPkXhdmtcdewGLjOrER/nifIw//2V673YuKK
V7HT/RhHULx4SfU139b1yYQCXqcUZlMDQ8JcSukQy/JrcmUk7Yg2jwJTx+TtwVWekLmoBqnyLoXh
hIE+qA2vnq9pVeXtow3499NcD2RhWn9lyJsqqZ2eFGx0iwYjWg03IpY1jl+Q5LlwZ2yGD/XejmyN
e2Yq/4+1nhcTevgA8NgbZnF6TGk1mSLxECzE47UCmE2RV6SeHZjk26IbbRbUlmfDRus8sWzCLRVB
CpMhFg0xFLUGwMuTnwhT+reD2VtaK/h0IiRLKvB2ETygyRhHieTbpJ0K7Yzo4DclTuoICC7S3iUL
vNh13YYOmTnI1Qcizm1mkaRNU2QpyNYQ78P3rHODZHMBEniMfYkGKG/h4OG/p6QvCiTOX+jxLaEM
vVzgK+7W57rj3TtjacxXYW4OK/hHUipnyxsDcHI5lDTZcC7XqSyV7h+KHTRxZebQvcIeBs+M3yk+
dK5ool9oHT6fiNbjrEc9qLqFK+DtkoRNI6L5qT4DgtK/wDfQIX2UogfxYWm8OzBIX/PkUN+YIVuL
rxbD6dnAeoqRRTWKXbn8cIzCyFSpC9zK2vvWCQYqpHva87wYKPbHNMjTYNhKm+LGrlCgKU0AmrQz
qWOGNmuh5xkGLoA93KfhXJtgx9Vq3nqQZE2VnHALOJFX0jElAKFjinjCQcnz5B31kw7IivImneC7
Pg2j+QCYUDO8jvOOgZjWEgQMHV/PnuFPEcbewq6T2LbrHJ/dy2rSCH4mqnhOVq8An4ZKbkRoHE1x
bxIIhQjqVmxC1xp6ABB+Vo1ERhg6hDbCHyoN6wm4LeXFgGUtTrsSY8PJFqY6+06/6WA0DjbRGujO
+vL0A0GmKkKvaNOiF6PaFIslHGr3OeBmDSOsmSuqSGHPLJH6K8pwtFYHoClpzvFrj+y+/Bko5k0a
tvhFFTb7HjMQofsk6nGMrjAl3U1ERmg/LqcfA3pTrK6x9UhZsoY/lLxAW+xg2M/zFoCv8n2CNEuL
PTbeP8k4UwlPkC+G7SA47F8KXKbJSZXHTvGYLsuAxjDPwIm1VHzgnZaxXXDZnADkyuPI/WcjtZvO
FGEXrq26coVWGv+sNupALYb7vjLBy7YrVfmLUT+SoDmMeFjwKJzgl9z8BJYyDfvcZvfNhTvVOCkP
lVVwAqX3skgf1Are8BVedbVyVmnQ00DTdSHjMMm4Fn2NnlAKQlWfjzqFzskWa8AbvCeP0iUPp2yn
lvr2ZeVkfhaCbRmWiCum1ZRxX9Ny7yvHaOC+vSs42atLtpFCX71VGAW+vL9etcPWcrxgA7rHhVbV
v7XsWyADfBpJiapDJRsdbL3vhIOPV4TQkXPiN+38lcaMjWzjenAQ+tNJVVG1wIK717FqkCxjJXgd
7CChftc3DjuT0VdTLtUiZayb3OYT4pEv+FY/7YEuFd6e4ctDxCbwfOsUncnthSm3ZrULvy9sCwkX
kaV8LtvFpsbSfn46neeKSo116stE0uDsPeWQhQiXnL8SHreRmR0IVOPBsd2SHiP76PB76BRBl3CY
yAx3XWlgEIXdyJco0zJ5WJuJ4WoLw2LPZ1U3/K49Hel68i+EvVif09uUCmxpWfU9l5yAUGPRu2vW
Yi7jHYdFad6F/FTlcPsBVy8FpmZk0eQQj5UdTYxrUk4xXgVjh3JDmI4s5howRB2FEWnqGxNb4CoG
1/Aq8BVi/F/Fr3DooVwwqRLSK/umF7td+Y5M0bfQWJ4uv+0M4/qXou+n6bZumX46fkt28mWz5VYe
uW2vxqmb03R8aAidetF/v57VEFzZ/F04lyc1m+ULVPEcA3kB0oSRW5AC5OfpHutJ/bgk2mi+Pwip
Yduh44F40LZbxMkPYdwCUcle/+yQ4gP7jeqALvuvPsLnnqGIgmtfQUQcVFL3zsEed0dsJR9yD09N
xMsdLsIramuGU6A7wN/xoRjFR5MpO5+wQcVDmFPLgh6B8mEtGQf2d43NKSG1cMy97fMo7UIxnTfO
OcrejBX/gMeSMjrVXZNTwCGh9938tqjwERXJcetM5a1KqbaMEutzbGCe37DX3I9TRm0xaZXhmsj/
M1fmGx7SbNRlEIRI6IST3Qzw/aH9uVwQMUzESaOOXqSY3pDS2+SXT1Pj8lHbqCH918D774fKVHqG
fuou6CMKbjOMS2PeqRCwtZdI5+yI026fEw2uyFZH+RY+x/GWmMQ1zAgSQFdbIaqDaA/yK5+dRlv/
nIS54uduugwN6/jsZVJZ/rlPw8T7LbCjRrcu5JPGG1rOVZMU0t5oZOU7M/lgK0rIl8Ar9LKSqow6
TTTzGf5v695fQCCgX97UJyHmHbV+R/c0i6kfS8sDsLGAnDYc6MKosryttgcTLpK2tU5GpM2yuFnf
ff0o8XFI6w9lnM6G9sXRIU7OetQ+Ze080Zo7TfYmWxo7DFwwLgMw4rubQH126D/RE00MGXIQW9rl
7L5B5rDtsjWzuygMIrjRribVaS+Gnn4JIaWzLBnd98WKzvhdwsKiI/UX8AcOqKRGleZmjOANs1qG
huosVIC7cffTI9tCrcYNgYVuhvfBHOf+rJE+Sem0E4P2Yk4GtKAltcw2ocZEbTh0VNKnpEqDnVLg
m4uhfuHDsOJO/yqtro7w5dxUhZwGSPYLelPMICYDy6bAlcLxz3lu0G+zpJBgzAvhyqhO8O8O9ZSK
AdPpz3+QKk92Ny+qsHkVYT1AsFg5DOLt2U0z5K2u8r3FmIcNd4pmnXP9tyVHFDtYki9gQCNV8oOw
qdRYZB3FSxAQeZh2CUreDObKwDnSDmLLuAvmfQg6HtQOL1PeG7zEgEGCp+YBB8IoqeOMjZSuJM33
IQqW7pYOr7R9lVXdcIVbrxHf/8yufjXPSkWjwp8se3vsai7/EcSANyyATSn2m3rVnThgBIO+AwCa
59MqpQ9+4fQT7/eHNla6Ms/oUde+tVycZpaS5SZCP1tB6zKqGyRD4D+ykA7SBRuEpCFFhIAeblGD
80o8HdYLo0FzAErM4tg4FEgWM4agSxIJmN1dLvSM33+/BZPHSTZ0nz8Sc0y/QDt7SYAS74w/D6rw
5RO4qiCPqPXRgmiZxCyVBujg9gXElGCT6FWjtU3SKx99Qz9SIWvMFrjnIKy4HRhxbZbopHh5mlrm
5lDEx1RzHlF5J7o4v6Qv63hy35zuJmAXMMbAkeemesKC9H+dqba4P4Vx4RqsZNdWiFoypyZVYbc7
qg3En6nn9RCUX+oAcfFZI4gRdNRef/0IMlpi1dy8ER6QTs//ZzaXMj//8ZxUDIGz4RmrxDvztNEw
5XGt3fxXE8QQvE/eWWq3Of+GMNygYAOKWLI/yCDb3+m4NMT2LwsVNqonNtLz7O+JLEA689pDgCW6
FUgsjBPIPf+chL90MJGeEvrYeTPSkK9fEpao9Y9A0dGW+kh7hRGWDH3ZGkAEIGRHYb9KKE13udiQ
QE4RJzv3dHrbmqKp7nozYppuvwfoNW6tervabd2dKEXPwv/lvofsT/d5f5JR9ZvZ0uRm78OElPt+
1fEE5nn3Ch1yBUYlZwDEtVbwpnjjMt+zZB/VQeT/Agy6maMGpapYpLpKMsa6ZBoECrdRrqP5wH80
hrFZnoyTX4L1F86Mj3N8q+pbEagLDJwYBfe9bSVGq071s8Qy8m5uTncWRVrurdGMeDMpHSvAVY9T
jnRIg2N5QJcRnL8E5McskpvkrdaDygHEhU2aB5JFAKg4yn40oN5CQ6NXgN1DFhwhRf/bMDF1ii8x
PIW7LtTX11HCryBhIXFL13EUW9rl8toka4VLN6+Y+euN014+H+5yhszJGRriRPn4Yaq57sXJoTW7
kjWBRDF5uXQF4pvLzGfFYW2gWMiMkSskELjmlz0auamQTcMX0RN/Sg/UrVG2+SRcpUH5F/En4Epx
uU3HvdbETke8YnzTlo7bugLxHOgXVospOiW1NWKUm1ICoCkCQdO3k/5y0V2zZ44XrwsABLFj+Sie
ijH0CmhC7sXkayboV6Oysd0S67CqhdmU+vft3sGB+CEb6d3mGbaEfGnkghePy+xvDthiDgZ67qTX
wkWYPNmdsbd37Aheb/BxjGCSlkfgIRCcsuZjdN4MI2PMeXFwcfUfcz6mVMyEH0IrpEJVRjuLuUqu
Kf1ymAT3txC5p49bZHGHKiczRT2pXapt/tZiyqal9DKHjiKhV6yf2bc4P41DbzpGw69ZKZXRLJ/4
sZYtTmKLPjFm+Of/xNBKRcuwBtiGYgIRMuqx7VqMQ5RXIlUMne7z8+n5trXRLCM5e8ihYTVr/WaK
IcNP3ESI83kSgHFlEGG1VM8iFzFtrmasl5f9tBSHNFjQCqLA7vrbphNK5eoRD/RdTw6wmXHtiSQy
v1gyXN0d5IuB14iPgvGyyFScdPCqdqzqRJ8nPQRDlc4tmXwwhzadZ10qtt2e0FqWX5n//Va3XQxo
ZZ6IarRxW16RZWqLC66/PiDM59fPTM1dKFmnoQMiWgemVM8J7tCqY5VNpkJCCTNetsrmgB/QJpjY
FA+mu9yrPQxna5Ven4nRr61N+nOGLWjO/UAt9lo9O5nVujctMsfx+Q7+7SyIYUsrUKQkQVo/8qhG
xPgbbBJ22MZd4SiPMGwIVw4zguyxk9DLxiwI5h97D/cHIzi5jqaut47jIFZWfQu7oKwk70itzfb5
/1Rwza4xLTv/wd1K2tQroUebvfxWzqAprb8AQDkvbQqlJ4mGqzmY/uh8Gh0QMKxNNl3PH5cxpMgQ
mcBB/PLCGdDDrsIJCDbu4G7vdg89ifnHkK6rB5PWGtv/FT57VAbFU2FlJMzEcjJ6xER+jVPtfe9X
ZIxnLZGB3ogpjUKsmdhcn9TJlaQCPnk9WdkpJishi++7/rVPh2CnQn6gVlQbxfGyPSNgz4ZOR1KE
auEz60sdGeaiTskfGpCcf4EbtmTsem/zsO2pnQQIer1RVZngQ+SCceW7i94t6IrcuU10fyPpnefK
tmPFXVoKlPr4QOw5LVbYRJFU4wKr7v/6pi3mg+GxFAFJznUxBLNkvy7TWrkpiDCLwL+qG6O9z5g/
qj2q0qXkuc8qf9PsmFOJZUSQaNNqTLIxK6XAFaB/PXmSkMm+o/wgTXc4cyzhfP6S5xfHzIGGGeF5
PoK0/MprLiXfCzd4uMF4YNgyFJ0marFFVffeGN7b2O/PyOMUykNhxMe1O7XaT1M0v4WGmMpl7Db0
UFyT7Ha7gwfncot6iyWtefR305nNjvePMhqWkhNqD+VOkE7zor6ZOrTdPzxwpZ/yNMePWZ+cv/jI
u7BXRZerEdyLOUmosA8iH5cVLUfOoVgjQOOtNtYfC4jqwkO79IvLCayf7/AMXuR2Ur/kZSZ6x+bN
5BRgb/OR+Q6NUrC9+tH/vkv97PdFRLIkJPVm3TIfCkTUYbsik1GIDnVnHpFxGMxC/OtZqYPOqHEu
uwWHTgqy8jFCivae2WVyWC+4q4jDTGAHsAQQwOIe8ESpe627GUCYYUzOobTTUl9lYxqEfeIwfZhH
zZ1ZhOeUTp/3HEzkxoRWt6F/FMjQXCKqwF/mG97Asv/wCvmyRTOlMywZGl01qLSaon0F6IsZruax
gomLCxD86BWs+56I0OwFQ302Fst0iy9ZgJH93YGAgHm4lr6Emm0esS4DM/BT7qx8DMSDqmODqyke
rbXX640qwDSzQnBYZtt7t89tXst3TEHbSmkSjTB7GS6CpEZC5CUuhhbJiGo7UmvaqozlhsWcFw1+
0Da5LIyOwcoOBwpdD6INeWCVQ27xnpWxdAPcP6+F6DFrCSCaUOTKkmeQVTvnO0ws4Ij9iFHVhNTe
6UKUPewl3VrNmq35iOKpxPfaCitf3yGC/8qQUucUmUQfAlarppyzE4f0k7GHtx/sU1hss14VWbgK
atbtTo808XbpbGwSYgMGb5LT6MqOIPc9NCnSa65z4uE98v1Pj6wCe+B+WsLBCtIAsPL98WUGxrC6
R1vUQNW6+8tsMTTuFOh4b6g76JMSE8I+xP/PYyv87fNj8TyUbqKDR+IwZwgfElm0UV3a0fYIP2nT
FHjzekNZh3Pko58g7ZvknBFw2qiDqCRNNmG1IEfNyUS9eB3OhoS7M5q9LTsOc4OumOfxYSCUercR
+TONf4vvFLTYNC1uGQPNw1PBtw5XCQHTxX4rLO7Um4E/6apKzN+wOUS/OCimOOaQyNAzOCM85Wdn
kCBU4FV48xa/UmoD/RWCWYlCishChY3oCiTJPqefHW27XDXW+yOYK+eVhLlIr7WUE5ImWoNRdMIG
j4K88SmvSZQnquz0s5f0wXXEdWPgoNzh4k7AdkT+z5nE9R1JxxA6pNJKUIWzQBa7Cpcco1G68NVB
jdGCP2Og+vRUopGH+KUyRVpvSLjWtzIXWhSVYijDwYJwlshoJEWeyI0DuSFX0MKhz02MpVV1vuml
fgZqSQDqG0AE7uQupaasN6KkzMeLybcT3xE5UeRPKoF9dge3kr+wzHMzCZW1tvIB71xV7iGQpx50
mI3LK9noGq8ShLDa5HkPoeEAWZtHiKJ8PHAz5OZNcV3B7BNpKlW1pcIWphtyaVzPHt+8uRetkmVT
AAPwA8RoTOxFgKeIhXWIZzNj3hvKtonlBOuy67fIuuRKEEqoe9RRNjyta45Gbn3NX5ulFHtRdg2J
IWoYJ3U4oP/mQs5BVVKOPd//G+gOA0tusU0KQHau6JNuwAlu95+FfS2RylpioEfu3uVYzQcX0DaF
7u2ef3EqxuvP4AgpqlAQg1XbG1Z9aEsuQbw3OwR5N2frYF1UdbVvu12mtxJ4/2YnYeweHoFUy4ws
u4B3w6OtNZE/RKMWxO40obDrwBvPJXQAPaQyrWjzl27QbrCKvipk9mGygIgcjp7ktHXK4+qewr99
3lWlJ3S7sS1dHviNb/jWQSbm+ZckT3LWyPWCQtCSsT7WOBzv2/csQKa6OOTIaSPE+YIlky8fwJ3N
iT9/k91QQiePZpwCnhxMYF+JHWa2a1rdrFLE5oSQbQ5V0darct1jmAlT8aaGg2a9+xuBHg/iny8H
DH9+fRlsiF8xrS6Te9VSAjYgrqbAki/EtOGTfx/FsTwDoDP7bhhGc6WY18wkZb9Ceg9HgDU+7maG
mmEeFgGKA6tDEQbplt+KKNEeCh1sKdxKoXqpPuuc1Uj1TjyW2GJ0iU01PxiX5U6tGEagtha1PP1H
5+MGMDw67ZULbvHt8Ms7rXS7SLy2Do8FnMv3clM318taWMNV/N4+KBJ+YqIT4nhDxoHF+9CH3Fb0
RtL5bueEIwmOW5lHW0DOGVzNKwbYYpptCx6D8XX9QG6aQ4WdFkcuGdtn+Ei6vU4jhPfkZMNZkpAi
N8+EORkmjrPNYxdr8PH69kA6jcDSPq1vsm8M+AMd2NXQq3wLVOW0xXP13KVyIpyKGj63nwx8qwuU
jW2ST3IzYbtUOB+6J5P+Pm/c5u7GyQK8x5l0D6J4KY+CYQactP45K3aMIxaBcYkMnAiLx26dQlD+
94es3mqcfayCgq2ZUNINFKoKByy3qO8HmkDcVzuDa+ltc3DpMmyEOrrtmPcb9p4+MFNDy33E3x9z
lIhi7gDt7D9BISWZlkwPC9USroYdpJdpkHJGa73T44nTtkFSA3VnMd9wzKW/MAp8AJzXSm6tKRrK
OlaEgRhImbzBwo04WRwIZdBAnXgil2aqVUIiqP3kB6o3IwvKzL/lFnxsWE7uFjNvbp5xbmexCFMK
UwEYNipsUuwez8XqgvGvxcxftCHi1W695cgjwYljcjRmDLRD2LexVbiZ9D3b+srPvhCA7NDcQsF1
hc9tWa4CdAIBtVakBM+38YAT3Eji8Z0Dfy4h3K8wbAExbegbVrYbKrYagw0t58TBWu/A5Qizyf+2
cA+zByqZPWr70+5qTxE644xcrBs4StyJtKN0HHW4ygmHpLAQDtaFRwD4q14ez0Iioj2AheCcqLfI
esBVgtPq/2SRVFHEgqkFymTWfspOZGgTocIXbsUdxTUpJW8ERYVgEiV3wELWJlyF9jhgkPqy8LD0
TSsaIs6U/2LFTjcJosds+4h7t+OUsPved4M3V1Wis2f26Nxf80Q0GT6IPufIXbS5otsEx8M5t5Vf
n7G7h0vVwTFWc0PcJIBT8wVZFxpf7aq3s8Xqst/1ApXfdya3wB+PcimPBI+52bZw2CBmIG4cU1vT
uba34Y+zk5kC3mTyn/y1teaF/DmJq94C6fBpY6aYEqiwHOI9Fk6cOHIFKVMAeCywgascm2c5zuQV
eJhnNr8WEozK/RXJyMX9wWArgzstA+NSZcpW+ruqD9LzqsryNdMHeIjNIHFYeuD1tIdsmXRSnJzQ
ImEdoNjwcvn+SY18fiUoxe4LkHuUi5yAvey7qBdwkHQkRm7XNbaLLEcUROwiZzlLy6hZzZSkxGPD
Cg3NrOm+qUUt+H07bP++rHAVsyhexw04Zd/t4OZgLQI2RuYVWVJ0YkLXPEKMb1drQqZaABZM5VFk
2ZWKGT3rr6OtdYnkEGIepbWYxVFvIVkpWGiEATEOLyERPxhzY8sK8NO+cqdpcdph9rdbTusMMJKC
UbFBN3N3bBOgu3WO18iG6G4XwK5OJUtNpvIFocluYfV7o4/2dS4uV747kRKDSfoOnWdbrDZhMeza
spVBQklz0RkjTD6mKEEQ7tMISyNmoRoGcoRLUpIVBmEtrTnNO3OfncpWtohP/hK6yajeF1HwKIWf
A1lpkmhZg0WAlsWo0M0mFgYpRaiNVsx4dQqemGz+rOVVbq9v5mc4qA3C6WcMPTC4iJ0Ypbug3MuU
tF6JWsbQFtb+K7YX5Jqtqi8DHYNUVGR+jQ6ukFyeeaBs7L0uKrudafhtzxqUelDjgwMQOJH3Rw4a
p0o8u1WqN0NzzXyHk66YWTEIoqhlUa0a4yDkuo80FShXOlF8hlxENEmQmJXLjP6cD6Z03j5dDVtt
jiNfzDpHAl5llcRMU1NaQEQ0j1NGog7qJWz9utqkNU8037IlH1D4mkGLv95K1rOZ8M1niv1sqyZw
CcPdgWX9vCKJViKpZB+DrtCqzAY4zDbgvA1NrCiMcgpbI+efZee5YDgfvVIyxHGwzKTr6FZSTm8u
u9dDjiWnZ4GIpNPz2pMkte3H4jJysMWbApgKP47RBzToBQOfT/m/9K0pcsWGlNgQwk7/8ZSGji8q
+uLuoZr/jxJzMDqAeg6EL0mDWfcDiI6+wCrFg3c4IasC4mFQhpT7zWMVQjoEiAkMUVJTIq1Lp6nG
3izfuQ9HPX6AYP72t/a2Qbj43mBeFixd3GgdMrrCTTO3lwkFBamTP9mEjs8wlqm7kMDbjEFuBCxW
OJlrxV78Ccv6EAHGKo6sy0FYzjT5Gxz9S1fgzA8Vdyj4NHH2fzO0RfuKXWN7ALKqZBWd+JxB6y0z
n2W2dDw6yJOr1GT1NL+LAa1mU+R3tv4VJBltOa2qrlPC57vJ+A/+YneemKjMzXTR2gxChRY7YQHT
s36O0Jicidzw9qiM3oaSpZMUa7KVGAtPsNozX7kchP8NBiHfzFyYd+NNeLd7ayVIv1AxDw5//If0
iFnJ/VQ/MECNRY6F9KcdmXmZAvblkUerklsDOXBQ90T8E/QDfaQxCVCRQeTbxZGPUNszjZ/elgAc
Mb4W/Mpx9NKCtztyYSeutwxnYZxn4cWMxezbma3M3sXV3iGhj4amgkHvhfcO5bUWDiYvy5C25Cfh
cqBT6T/TMIUYedc+zFKzwpKL84Rueywbu8YSkMISiRD/j0Vdnnf7pcDVINPYLwxrSklQtm8wvbTC
mRz4j5WAr66kS7V3dhhport+lzlHhHW3yb7ihkS/OAUZZ1KbWfQ1JH5D65oIU/Ax1YUrx9vwccyi
UbnhhygTPioT69wlQ1rW21p/DEpjpUtwJcw1TQP2+SHLG5bmz/6Z3oK4w8Kh9QUkfLeUQJs23YKS
U4UdfFTFemtOOmRBJ5FbhcDAR16nPgCse4bQuk+L7tsjR0feupO4veDNBve/iHPORJ04ruETcN7F
3GGBNfjWSUY5IaqDE+eFrKf6T5ZBWDrxIbRMcYSKr0jcYtXroIb+OGb5VyMuvFYCJUUgodRVO5vG
zqJxG8z1wvNBKQ4PAkF/rcTrRLLn/+l8chCfnUnkPlVa3R9ly4zg5Vrhh92uZYtKZSic3TiatBck
I8aYAj/lU2Gl+q0ei/c8Mkci8SHfrcG2gr7lf6NPxRYK3mo166mZ7rce+l+ElGRO5OxCWZ7FifUI
3OqJR7PWMrMqmgaeRrUJCmbs+6QZPatk38Ra8GvVMvhhqZd2PkPJWl5AQZgrCjrzKXirDhtzBzkr
jSec7v2vO+3r5AkLsqo/aPt0otJxl0oYlcdRNzviI/0pMYGjwc82Dvmiax1FublBSqz/FeW+tbvh
J5JoxkIfAaFTbGC2/i5Kzm4D1/+tUusGwVjuvwfTwm14JlRX16dXEv9dmtxMG8HeppwNJiw0jK8l
jVBtn4Utrmzfhqdh0XxeyLLMVHUUQwqIxe3sX3AtdJ28Zq7r0820yheCbUoY4HtAFhiEOAv3LOXo
plil5zbqytmt4iUuZb5NO2U19rD2iJCch+qYueaTQh9vjop5dy79LZvWjU4fCyJI96Nu3gPXFAg/
5hBV+cuWIu+/VpzOogkCMkF0PqweN1iPG8ytgTwebqA9ELsuwv+lqFMIxBXwPQBMIbHkrfIzVT9/
t8gjbhjN3QtFvKZ76ulM0WMDmFb/zXXVjdSSaOwxpATB6W3gyBJ+/smzwG9J7SOaOJ6P5PKtbH5f
PGJM2ZezGlR0XTt4d9V04Pu3gDaI3sU8zpp37T2bGhu9ROMDTYxD37e7wpKvBT4XQe/r/8Zo+kVI
vEsIDFAPLA7IKIpDdJxiCe4SLDWgOLXmjQSskyW6vcJYCTbu+WZ0J3mtHi10sLJgZ8qj4GEKeSa3
wPxoP8diCQSvJKUO9jiT4WAHeghU065ioiMb26rMa2D8qftgASed+0Art0CIWrnAXC2zJRWwzwV5
Lc2a26n7YNTsqrCkwH9/uNRwswjbJ3r2Xkkp9ps1FAdi8UCqQEgy6FLhDOWLL3jwxVHeIGlBCFq/
iG/syVOb7WyDs4eB04o83ZL51UY2kzdQIHmhYPQV8p4r70e0jzQBCxjPdJHZqOTxnfnQojXpy67u
APge7dy/BcASjuF2jZvpYANCalvKot1mCz2llnxq8rxVz2z3l5Td+IS/Y9QoBGrSKrKO3txEXmg8
24UXjTzntFBj26xpm1E99unkhPTOOano2vApO23M9FlPB+3zt6GKmy5dkEdzklfUn/wRrw9iuWoj
3rdbKEEny7615cL+rrNa7p4WIMRYBjV7M3uuN0rxDWhtBihsvBfADaErgFjilJisOR05WLVmVmjl
AVqYv0UsKfoN6uF72rl6UI22OQ4ezBmN2ArB/ERaJ8SMLUBVaMZho4wqiagopEb0E+kCX4Q1ZmzG
0T7tuuHSHX5ems3+VPxyfK387wmGUf653nHkjoUwv2kq5+i0bLwNbxq0qIYQfH+gcWpSG4nmevdV
ueIA0J4qoitXpAVomsez01D1sK+6pdt0NaBWqQ3PrxGfIsYMcxMpNgTmEPUP5ErzMSls6oq71AIn
ke+SNd5djgGnUG8ArQ4cxl9/z+Y3AV9tiRxJa2rscZ5tX3k2OTkakQKJiAvlOZdJvLeczfGsHxxy
oIANIWyfRNvaqVvBVEcQBnX2Hl9naDyNjex5E6lMk7sE8zdZDnxf2C2cqIN0yPeqaEYOns90PFvL
b3pWJyeBbYszONa3KbYwLKCCYHp8BupycIzbS46OXGzZkkYc0E4xAta8BdAcAI2cusEHssAui76X
5V7hTHpvyYnLGe78E7A9SwqoStj8a0VitetbRxTS455Pejm3sn2MdEO9O1AWD/4MSaY38bqV2iXL
9z45feKB/UuqjJfb2QDZOEqpTWbjZs3Y/YmtuaIDrus/NFObuvFehtK+Jlkpn0QEAqm9T709KXeA
+2wJb6boW6DHgBg3d4o+qwKLxhc4enJDROrBe3W3XLu/SPqpFGsb5HvjQ42oD77y2TJu1tAPWTG/
/yoG8MTygZpf7HeKomydOC9/Mnfu8/GiY7eCV+4JLB1JVGEJGeFvn/RPntg9SA2u85aEDdcp+Pyi
Fh8TwjcDu+FqECm31vm0O9AdzvaCRysrGt+3DK8ywCCtk4d5e8EP3dZPmIqN8q2x//HrIGawUY6+
MuWlQtuW+KQ7Ii8PwmjF5UZJTbO2IJCWnjkmdlGD8dG3kenbnqAhNasdE7pQubMoEbG3GBwNOpD+
BCTlk9AUNE3fERy3e4nO0Ixh2kZLU42C22v3LUkP8K4Ox54/S4PxdxwqAbvrA5flP/lP2ULePepm
+Lky0/3pJy3GkyClvb7gWYYiYxsguRozYY+MAgGD9A3zxjrv/eS3aGrfj26LbUGo6cZd6Vb8X8gY
JICqjL64ARUpLqXW+6cfZM0nRv/2uQbInD8k1TeiIoBKADcxFhSCCFzRVHJ68rwP9+8WP78YDYoD
mzxnBMrTx89u5UuawL1Bm3MKNDgHrqY7Hg/cJZR7x50b6Dc4CPYu/MdibEqGpXw+YobGvYWGaUQ3
ej2wkAZPQmX6htZJrKujCopIkYvRvMT+KKvv314hUtLQJjCEoB9rmGrtrX+nzW671gmAGaa4USlF
wo0nDcbsqVHnpuOvuJKMWUowZ95tEILL5Ye/BYvL/0BLVLwHzxB/CLsDMfXYgIHcHhFTSfui3+xz
j0yfrtPZ426aeCRCH3cgOrRqQmsdyX2SPTyrP3L2gzG1f6zlwul34HOGtPIJRoU55B+PQ6rCQjFg
MsreyM4qK4KM/fQ8bZM4VHn8FxWLIkt90cjIfE2wWBBGjV4qxcwJOf9xYxhQR/LBENYiNSvdDHc5
TyB/HMY9hUaTX47zCqUBElza4NJI734IFJPHpdHFpY6FvPrTIPDo9VRSCRa6BuKGm21u0t3XYQzG
Sn0Kl5IZ/CrQZXXeTr3CKRt+PG9sIXH8W16PAalxcW3hA0BgKq4Hx0B6shSPlV/S40RqBR5Z7cGs
JSQcFuT0jPM1DImq6T1peY3/PVzmzP/+/Q0z/AnpwlsvhLZcqUmNbBD53znM+D/urGubrTa1H9g6
NteUJVmPc0Li7/9sYylZzbP2+vGTix247NvR8C5GZ90Demz6tuRGSH3Df4K+2kQRHfkCT/ygFQc8
Szzjzqwcsa+XFIKG7l812SJCyUVQrXeTk9eHiYo013DNpWuI7rUSjqHZ5IdJelirPDmeR0IlZdUV
sdAZznesvHjRwIjx+QzHanJu0KHWRL58RxI5Tnt98WApZXDJLmQLhrtQLnMSr5z/GPIbXsrhXOtl
iKLMAhG675qkVyLL8MHT6qkunFqIwS9llC4wlucCS1IggbFkucOHKeZBcGQ/IwcR/SlaTALnPqYp
3Pdy+MJXw4Q5PP4hsZ9h6UiOzzWVuQJTSoZxI33/+k081oI3lSzLu+vngw5CabK/gO487LpKupBo
TzY8PrJqm4xwpgf1L1shSBY/MD5yk2ACGYJBnp9OdtGi4laz9fA8N076E7cmA8gtaQIndZMIolwm
D3PM+iVVQ6dRTd0gY4+cmQoNUiKgLXE9EWmXDrR+8giTsjPTfU4E+E58r7WFGgk9aWOekXvfk1AJ
swPpe7VkDTjY6beZuLhP8VnbC7BvsrZ0OLIt+/ntLOLE3Fm+BkVEUlwjE2xJcVIzV6Uh/ouJPxr8
dS/YQBJEzM03vqxqgyyP+9OTimYXM3Ep9O8wntLFTCPUPQwhR4XEQJnzkIksO8P0ro8YMO3PPVSc
BwOALZ8lD9VHyETeOq+MVfR/7cMHk5e9KlHlBnY6sWYF+gmZzJ/OnJJIeEJCTfqbW0HTLtdhVnYB
viCYb71JZTgV3GA4giUZfC9YvsQ5ZvS7Tl64qi/45RMg29xuj6tMRPWkUlngPPPuDJoRYyUpcj0X
J6axglz7Mu5e/7XwkiNJjmJMivmVB+Ivr7vfRClaffONIq8pTRbd3Pxx6kiUMhkNQpz8sfJycGFa
tTN0WtN9Gg3AeYXmO3IpH/R0HFJFiPIeKIuu5VhDIs2iY9Zt5qh5GPkSSJttr9OuI/av9Hh9kjml
dg5nhHyCVDQjPufNatdac9CX9XllDyW17cphKjgNRAods0pjAPxTlBeypLqxYS+yCzy7Y4lLSZzS
aoLGKBKavcaOroRYxpo/YhsfO6FkCf2xsVcr8PkC7Ex0GL97zr3UXYoX19xb/3q9KPbhmfe7uJiz
ZNFV1pMcvl43dSLACOpDNh1TVyLGgv7vDrIyy83TfaWvQ2Pk24Vx+ImPuyz6NWt8wkEFsN8kDIeX
HpZzD+KNCbsbLO3/mNkT6xra0ahseKjZTfe9Acgvjjt0Moil7+w7TF53H8tbjby/Q4rBTXlgCI5I
e53oOSA/llqr3Dw36uO2Nzp5wsoWmgGUAIjHf498XBSGBEX/C57Sr3QgahRFtV/dS6ItZzeNjBsW
aOteC+551xzII6c/v1Jw03qDHfr92afVS0XLmTFp82Oqlo8L5E2+2l/rx8eRwJVZYvFgqEEC5vWu
m5BEfcHAAgpc2QIZH3ZWFhhFY43/ogmDQ9YMkf5PDt7G9EKyGEI69MolTMi0YY7zFmNivQRpBwLa
Jnozd2UhlV43I6pOE254Gb09U9M1dPSkUVUKFsG3KpQOGy3arYfr62bHZ6q9S1Vho/gi3idtJn+W
aq4lLUGtuRuvasx6E1Or8BentKb2vxKPwBAQ/uE4F1IBVcL5ayctOb6Rp14mHiPos8RQQaVMZD81
V1ByUjkXtKaRzvcITjaVYLQGaedBo4W6oPf7uo/f1YIYAgJ6zrIXfHpKjcwp03ofPh3ubOsKZlHT
hUQVIaLYD/+opWJAJ+YoXcOglYFqxwrYifAo6k15xaB5qgQMvzA1pNtuiITZ72q8p+z1v4x1xEC/
Y7ELvt3sAmS7QEVN6S1w6p89cRwqOeGhdG1FW1BANRoLQJYbcLERASWfrQGLWHtS89YuzWLUfs0c
fKNMOYTzoMtc/AW/AJ2d8FmAIJ6DhQJfwqoV3RbdDIUrIa+9ajl4ghm/I52RTtsOXlkMl2QYvkEP
aWwaBYONV+iZgETqcr9169S0GnkXihjSnD5iV6ygqxE4rvbbaY0DSya8kVWOYL76vwwTHFDctVib
KWWDVCHRD2y1KSFZ1iR/wGg+mQvx3YILzr9xf1J8Yn/p24hzwC63IR1y9GM+GCmTlpRY/5mZsY8o
485O1R+GLn94gIGYTYTtw11zGXegnMPK8suQpa0IM8fcDA68WicsZwq9MwDp6DZKRmzuUehnuIzT
5dnzD1rmC6C4cWS2JQdU8WyTzBnYSLeSC66j44+fQnqula1X9x1FNtOCyfXUH/g5uOb4rwR1T4He
4Sjujel5BCe7c2ewk5GZ3iRPnp3cMljX8bEPKWQYgAyYoFzuWQOkm6jN9nm5E/3zJ09Nfyrvkrcx
l/2XpPTNPoMmgh2UT9yRET1oEe2clBsRSolwFYTMGfj75XG+1RLqW3Xp8883wvipbzQqDIBwH+1J
lTslImYKdCrPD5nr4yPlYIG5t+9VUnn3i0WSixMKeNESmXIfpoK1hkyNjhSms31mK92AvEvpmGn4
u/DPwnPNWV8X0vW4Tj17GXtlyeedP1Y4uNJc6gLhiyWlDaQ2h74UeH145Uk6/vV+3cBZ2zCQ+51x
7xafcGqejdLrYre4DaM4IxHNkvZjRJ/1cKOSHQfBsCu0pWAFRdskvI2KvMbfeZjKJjd47VkNb9u3
WwW7yHlUNZWUlyD54wjaZs4y3JMCZhCCIWXGPyVv2kEudW5fe7GDmCKwNOWlxXD8A4H+CgcoItY4
9v8hFw6+tDT63MaPJ42yFOzzQwuBPs4b2Wr0k5wmbKSS1qdL9VY6yPqPsG4IBlD7K3uppvu2avOA
9kp1By1CAUZHIL2yzeCF/HprV68ZJjm0/VpE+pM11qRsiFLkzNl50AJOlZQdpwzoaqBJayjPSsUU
0F2F57K2nzzjEboNYI+9Yx3Eh5bhuN/C4qgSc+cCYUEPyWeBl5SMG+LslnMbDUkS0FIJsqYzZkmq
AoTEioQ5mu4hViQxoIrM5/WFwDFBevr4fZpWq4DvRFWDLidB5WW9glTwvD4MgAvBZldbq1FOBspr
TZIUUyzJhJbxBL9sABQZEXvuqqWOTWf1zhnQ9WY9Er97YUTWxFaXDW2ydNVPpTkWr7LEZBzjtFww
zGfUFAxq3fDeti3ihg7PGZAfNnPMa2kQzeph3QCSRiuZDuw/Tm+kGGLS3UkszUW09tQMA73GLzPQ
oY/Qg1/4I6RZhkv4/+neDnhZIUKBUt7KQNURX6GwxyHuslyt4NtiXkhflE4Cf1ose40XSttyiI6y
SaACAY0TzrggnQ8ipqH7cP3SgVpvAtmtfGJhIcoOjFKa7hSfVauftRXFmo7Oi62yjQMAjaOD14yO
NMd00LeTfAawxyZ2c5WktBw0zzvQuPQL+WpiCyBDApT7Pqynsm8A1howlNFdUqM+a49tWAWqsI6u
bI74WBKEMJUyK1A6KzMOucKMtYJMaZxR0q7VEQJMN5T7G3ebhYorW6ld9o/4ZrWNkhEvDmYwcSwP
M3jFlZe0rbCxOC2xhqD3s5pEvtiHZ+92hekmI6AfhqIvUs5w2XhrEUo2qlwH4Dc1y2uIYA3dYGx3
hDBRpBhOZMR0+quvwwBaQ15jOkPmN0gaIH5UAhRP3uX9AQq8Y+mUxUqCaNk9hj9LbtNPFuLfzXXj
48qs8ofWPAQbKs+XNpNY9fhwaRAJsLLRVWwOnPP12ycHM12vVio96ehqGRoRBs+uPWDCm1ZdSbJE
qfP4H+YP952AaVoepmTwtqL+HMAyTHd9zi82+/bh5LYefaUGikv/tPUEU7f8OB8AB8r+9XB9qo8I
QjQD0qoIARO+fvfChhuS4tfY/b0wripBDQzSTuq0tsT+50Psj0rkGWZTRroypIDQn8RiZelm1IoO
BAXqzhdulDGGBTX8Cy2aT/535OX46cUOXi9lZvSAi09ZE7bwRCHqG0tn2Hsna7OYflunmg2TrVDM
rpCmhvVulClEsh0MEWyLDv1VHnPdp8WDi2PX9M0c5eus9ACOVlnOrGZzATQOkRnfehr9OUoaqYZZ
s8g29saitoHKeozGsbaIPuN0cFjKaIHAX0+SfeiVLYq/bjBd1FwG2Qh3/Zb+otRajVhoqk+MUdo8
IC/SmUsneuPpa9uHyNvmAmA/ipPzqo69DZ+iraHhivp754pXm0Q5MzwA0HOPi0CHJzkePYOoQCSn
AmFMd66igqEvalmK2ht/XDgbd3gJmQiy/R/dq3qM+XnLpZXicbr9micqKskjHGxkPsuVL0Wx7L3r
kdlWC5Qd0xKFrFlJIsTh/yjBir3OMFQt73oLAXuoKgdZTu63EYAEcaJCrj1s1v+hFQ94waIr+NPY
crQkhb0NgPhy1FT6zP8HtmXSYqxbEbRs+2+5sSxgllNpjZ6bS/SUCOvyGbR8pfzvvaYJiwoq9PNY
cdj7q9mw1W43LwHHT1vF6UgRT9l9j+aBW06ATbrJEnSnow+3jz7eiO0Y/h31v8rIvhD5GlGaUbG1
+ZtgiDoQvpIuwlmCWdB59gF7shtfzre2PBbNgokF0eH0lX/EmKYsQKQkVIhQI0keaq7YnNzn7Zyf
eB5mFnUjvO36W/KVP8U3z2cfZJGHz1T3ZDraKYzEqE8orw/s3uLwvOmv7K/SAutJo7/1UxuIqwIS
MgFHGcKGutgn/xJ7Iyy6zMN8ovZWIIHQkdXaQN4iGWMWQdWPDex9rQbasKSOJBkDPsZL2wS6CWyo
8JbgTtVlThGWKSbzrycvtB2LnliQ4VeDCvkPkLzxSXssQATIvTOi90BJrq2EzZDWO105miJw5pOe
fTpwLks4FshiBtMS6APxWtWNdMRRRAXE82CXWkJEvQWpMl9Hmqf9eY9fB75Oy8XcOp/7ixzX/5fK
vlMKqQJzHi5cXZNKJzCxpmnGstYsSDgm2JrII+vzMBbIEoIrmkQSt0t8mvv48og3AfK/3cD9Jthy
FevqDVU6sl2XxlPTJ2U/2MA9GyPO+O78dKl0yZrlrDT9ljJwIqLajeByAhham/z07fIjvQdwy9n0
wvxwSCq7hqilzg9ckBeVj6qt+rlttuSBnA8eD+5o+OaVFv5JzlZOcVEFjm/PUBYtXcxGyfnXO2L0
0sUk7JPL1CNW/I9Z8zchT14oITqwbsLJ5Y+BVyJz/FnEjVAI7WNc7ELBU+hSga105bqYuxZyViTf
c0aHAFl9k5HkN0OBFw76AeOOcvGJkNJ/I/R+fUjHTd6M01F0QxMCIP5+UYVbqE41j6IIicaJkr8Z
Ovk3b0z6zD1i3lO+otED7jt+5bkTQwePDd1OQa/u2oe1jERO647J1EWg0ZsXjGm7BboOaJ+nW9wq
fyGPKCX2VCuLEJNVCW6zQap+CpRGtJRcQMXYZ0MGhIw505V5QmQbCUvM5txs72ltOnp3QPFrd+Nv
WuAiL9su4iw8L0t31zq7YCxV3wqn+sgg8AkmM/bF/xOOY46TSIGrayHpAEbp0zvRmhLpmHLSLmnu
k2JOANRMdLD3rUO0Ud4Jxk8E2wOKCqzwGzm5J+qbwVrUeJhfs+ByMAoWPOv32ECnxj76Vmt/1O8V
QZyNbZj7ybOEyWK7W/CJCarGIxEjiL7rZB+P1Kzb2VV2Gp5KqyKiOOxRwDAl9IBjZ0k5ZLAc7mqX
0q+pB+EjvWv0XWg5D9T3DDPkl06jX5u26kQcHNVWOaukwPbdcVHYnTC0/GkA07ooNzdtRWtgaOYQ
8UB6gksSYbauGJ6I5DAMWwn3TjdKoty8STM5aKflIg6B+JIrW0UpryaiERLgC4cMTuLOaXm/2AQq
mjt6+7c0YFIw+4KxwbPg1fWod5524BrSJebhQC88RK5aRGYkkU71hfllofX9+7lfi+ahlvIdukwc
kEN5UpLPg+z2GmhS0CnC9W0SBOm2aUzEqGP3zz9TqjWAVcgWkR7FiSM2rlnete6WDSMgiNNBtnaG
P9io54USyV/hn4AMtKqP09kz2lU8p1JSHIC5SK4pqwVy5UWpWrjlXdoLaqO92FNeP7KCVV9lTE/+
+Wj7L4yqO/7NOjacvM4Jqa70KAgW6y7SLbMHdeC8HdIsfde3IcxCbOMr3ShR0jia2MKtvGPtRdkG
J7z60s8AYReiGRRFNmU2UyZtJsLuBknHZJ1Q81N8saW6CnonclIzbJSZzDVuyC4u4W4RnABwTDSA
G+iBDJJeDLPdBBY2AQttrFpslkgXbZVb1Ugqim3NgeSZXxKRpOUDQwdNpX/yku/+tvWoT3oaKD/I
helRU5nkKCp4NoN1J5DSvhjlw3EpX0o9/DZk2LaPLPHs9id+zBfWVChvogGxdKoe9vTVzPQ2LpeN
WyEqwPfn9OSAyMAiosUU6QHpU1A0unwiv1gOE8BKr5HyUJkUWoEC9JBY6wBD2M/OGP71TzFCcx9k
MCd/h4gBRHftqo3VCaYLPPSH/IvLm94ep45Km4fb4HVuvpi1a+Ak1CGBETuliaDvUhnHanGcyECN
i3FN79il4BeFauwojYuP2xZThLOAmopgWwbrxHpRaWhYK6ftV8X4u+vRFnv1zHp6GXBaqmvkDQot
4hA2k2u4P+DqJ+OPvGspt2Jqy6VAWF3yFs7qDguVfRr9xBGZZE5PrBKoK7q+zEuoOvk8s7eHrAZF
9pv3OWyLUvgJP2xLIshcE0ywqGGegItAAzBvvtS5UnIQ+sfpFpBtgwTyFGat0D4mJODLSOdFfczV
MwCOMhHLRBj7yB/PsTeM0eS3LjNFpGCx4fVbvjxgoEkZS2+n9VGhGusywCMz0kiNPqXJhk1OMTdZ
P5VPrEtRkEQEr4xKSsuxozpEKiCc1hDT1HWH3IsWejK3LBIlUOn3xhvAsPHCwGZBR3nMCzysjtie
L9ssGzUkwkTHDKoGtjuvkvucv2STqVdG5n+AFy7HbrL3rsNY4JOhWuwh87PqwUQao6xOAAw7qloQ
/bnPA/YPdahsOrkvG3osnh7EfuJFE+mENr2O+HL+yU6Jr9x8UqI37/9uMIZJ7nLd0mbwQU+1IHF0
FUeXhSYLcyxqUFocCqJqX+QDx+jtm2dhZnZOFjZTAShEdIIL/Ud1d69YZKkynaK/QxqHScER3m5x
0ddk9QHGMfOPfD0f94kVeHcIeIDONGRueZ86Ck8la1UTgPCbiZK3W+Cg6U7Tp1U8JYkjhMOfDnmq
Y+QWauHWbya2WaAHlS3RLL636jL66t3JMBJAcbMayBGAv3vI0Dpug5kjDXdndAcM9c5YR4yfOqJq
JEQ00/mQFc648NQVImYZCRPFUNZNwZfPXFdtIpMJjQawo0eavxbRd4wKYCb6crOqzo1SOkHfyMwu
NrldDY9Vnb11S9+s3aYCk4e2eG5DOar1XKm+SFFPu9D99C9ZOsOFMhmLyM3gox8iFQlNFqI8Amzi
53o4LF0shHl5TddGaPBbqK8m8/0q8JtjwegVvnH6wbrVRZgcTGd1WTskw70EBt4jGNz1KdkwaTvM
rACIIg4e5QlUVPGYSXszeLWHkFxTnv8NN4xwwvByA1Xp7SToc//KAI/DEjof70e7CRXquV71L9P5
+dGMagSyU0rcxMkHwVGPwZ3NwKCFJ+06qUVIc4zQAVbIFLhiPgzsvSa/9+xaCcD5oxv2ciqKswsr
LcCRn81TmPQVH3Ri2AM/4fu5cFzM1r+O3DVjy1azMvtvshJXi+hKviBPXpiPBAJy5WqDLNlzK2fU
sxjVt7BUdiRzrwqD2MIom5un0GBf5YmELuTrm/XBTQ8qcNm3NVepGDpO1O0sHvCtDkHGupxXPUPI
AkJLmXIYXl3qvHIr21KAD8yawjlry8u7ktG3/N4e2aEhUCkwW+Pr4H0I/HNdObUj8uBSVfmgKurj
PoDiJqUbYl6bhMFlq5OnDMB1+KGd/HK7TiKtjOVJA9JseCy0i1LS++jI8Z+Qm+5i4vhWZrMz2Ta3
FCY5rvPP3ssboKJXiNVFAo4YKUe1i3rZLuEvMk16VbrNWk1HT37+MdVrmMAzu5F0hKLw6VMeHLWl
aPuHvg2S2yyV7Uwqrn9DqtA1vDUTG34ECOA+7Xxqfd9ZsJPj5RR/hhZQSgImNqWKL50MHLh3c6r+
/tWHkm5kvgawR74C2I9FrpEceJXXq5Rvb449emKGPCffmxX8Y8WW5qEocFwC90714SJ0W06XEbk+
Et0uaPKi0GiBjkn37YieGma5T58ImHoPaQkyB6qlqEaFEKJ8wmTlPOUC89fVebsSfPJrt247OMpo
ZKW2Y/XBpoFJyuWiBpP+yARYcRYOSz28mVyvByywFRhDn2+s6Xxj2fQvIu/mosnHn86AdD7kfM3D
dnGAL9VKmDzFy7R281kk4jIgFV1neeoEZ21JuXI0P3Dhntx6xrUsVjap/EnzFq/0MnKlJ0HEGFyV
w293VyDtoxjCUAeEh3gCPnnH789WNOXeMcL2Wh4VDWzAPAYtebiRN/1YH563stxHBUWE6kC96eW5
/0GayS8tJbkCMJYa3sXXLQNwqz9o8i3PyoQTpw7ZSj7wGFePzPcYW/o9VD+5nBtL8MWmQ4++mLpl
ux7fWI9RIPFkiH0ARV9qh3APw6UtXK6UP6i0I2oNqKtUsMqlOZ+xMhxD6pmO+JYFsFdv8gf7pTrW
T+gAF3cYqrMkQ5oc+Ipgv+RfWrtw0r9w5Ai9B4dKKmWls/fRm1qSpQ638pEFF9ByrM8THVIzOWGm
HEesSRelcNa2eY1vvmVaHaAGllLPMQQQF7swjfO3hNug0fKEDj01wesjX5FF/ih8NUcHqe7IhKl5
bSFXval7jFsMJXpmtfFzkeBSwWrsfUyltbUmn/1VjmAgPwqL2wStQwMBNSRu4SmJgM6f49ehnklh
5tMUsWwTzXR1z/WSkupZyiceNJ5bg6k0Mc+RauJuha3q7xH/eV9aIBano7MFu21EWWAyhHcdMb7T
NPaflQKzamYh25+XkoCBaJ/m5PVSSS9TAvxQCaFVMPzXkZAZ8Q19bZHuXou9QGMZYnzDQscjALD9
0kv/2MuvsqL0be1yixNkloEPjZo2N4pdIhf5gtpt95uwIApFEuzhw5IsnTM+vM3fEOWWKkQXDKtd
2Wh5W9i7HCywEJrpUmpTzhEARJH/hHGnjztQnroj6hZPjjlRCgd6yfnxcFhpJw9eEsoW6W0MLNIc
qU+XY49PyGBqbM7HPBPH2uxtL540VfzQXtv1Ndnk7c6JQQYuiTBtVdjYmwmpR1m6+NQT92/OkkBK
GxedBysAgZkq+6pbK/MrR0zzLrE2tdjO14xfVbp9XdHp3UcLy0YKHFi4xvxXJEeChRh4yCI1ne4g
Iy2frTbY4SqM5RakOb58oq75kGxtmAL7Rps2BiGrOCZYXyfVCbH5dviPVfHKXFyYhZg3E4GEGSYa
klWO/KqMwvXWNBk8uvNzWqFl0EUzR+nAVf/fQcQnvobFrJOaENHiipZ+a4uDrRibfY0xx+QCdHXv
yFLhfPtUEjqxanEQX+9rA7lzwS3Viksmif1bBmWKJ6td0RtTWkXmSQLOVEsU1x4633bjoBA7Q6mo
BGao4O8SAru3Fztn8L7VKyaNCpEru9+qNkAkiW/w5QPINHcfAkeKqOweCckzQA4RQGFy9DppXc/5
L8LzD/kjFI4G27PcyeRA/+yMJELmoHHmgggIBS8UzGlnep4kJT1BOCebYl00xVEB8oTDW6/MGB5L
VWNNd4lNL8XzY5gb23s3V6LGjsmz9hInB9JO+4vtHJP29IqPK6gVXaRvCk+X7EF5uhSAU+L7rvQP
4QAULX4iwxw4ELb6EuGItxIbpveTh5qnamTPuzkQiN66H2KbQp6s9GSUbdrJlS3lYK4WBEPsMWcV
E8IQNpqRN77mXKefO52PGDlihuEBk7xJNpEwvStu00ZvEWTIWs/a4I3EIN1cDgb2pF6FWWr+LLL7
sCQhAD//cjxNxvR4UDSyzp9Pi9opYa2VJsnjSEjLw4h4wT01TqmhdpUjm8nqK8xS92oF6+BGnONY
YshqgimgVKloYmhhUI0H9gMEUa6Rnf1tG5kQHoeYSjw1VS6rjTY8Wfums3J5qz+cvmZVhmnzq7OQ
BMMCS3EphQhuhOiDij0f1yMA5lRIDaL3Uz5QUxwoN4M2kJBS/2x+BCFqOO7WOkwgFQoAbsyfmYoI
XPQGreuY0H75i5DWADZdFbhkGKhK7oh7i9GzIQFoIhNvF5z9z29ElsVQNyo9Hm9WIiMPkpf7Bmxg
3Yn7Mbw/MelQj0jnbf1LbzOj7yqrQop6Edslf/67mcm4QCPSF+icJZJkaA0ejxlJGpvnDyVuHxq3
jjw8rL0jYIsDT4XL3Ot1yxsBy0AaVvgw3Ytr8CUlLk5OwmByLGnBtER2yxBLAIKAKvvIO9VSA/nh
OhTEUwG53Du9PfI/N6GTNIQtV2qtlgpS3zy0kKdwScjMffmL5JOKNvLVQJglFp/vPk6l8Pz5BWN9
vsRYMKxcyM45UwmOsUUXOq5ZuFQ42WX5f100W+WRxPnGKn7ds7VpBpXBwtY0u9Pkj5kVOEJlN+qm
LBaJaupMs/SYMAMJUlUDDFCOT9mkX2r82pBYJtROO8RYe7/DyrGbtaZ3lAOCBYYntNDVsa2TeLCF
zsVrsnqliMz8bKBcgVhcLVyPL7zNrpHMuBaPsGvteB9dC/v1kiVpyhuOfeih3XT9txXc/yFXL7nk
dZ2PaiAy3M8tBBsvcrOGSdJeQnaZryf9mQld7Bk2gjzqtn37qoIGRIk0U58V+Ny8kDm2TKq4jRll
E0jU4t1jlJ9A/QD2kN1R0EqoSPMP+A6JwNvgaU75JkjXFzzgcKzhl8GWwgNgX5DIcx84BXwc5DeA
Zf3/lKMXDC1WcnBMPdrtnl7ctrN7D33+CfHE8LHsJDXoQbRmwychdbc43JgXCVRwrR4aJmpzA9CX
svI88XmcmAS+yr22c8MGmOWurgT2mgeJp7tv85ZpmwJh7biCwiW11CisH43ebWLmsqHPDbr/ZCPH
7ndEhtKy7oJGDgwrDQJAnOJ3IrakIe5BBHUlWiBxps7yNDwzVe4lKdteLN2dKTNaPBZFKvJqM0t5
vQx8f7msCvDj0lYlNotzUQT4zKCl9xksedDCIdnBP52cpQCiufYeb6iolk8StfrXc6/8ta30nGMM
WrRQ9WAwyM8T19dThC1TC6ng6+JOiABqhi80hpBviAN2/xh23P5jL26S9x1E2FN9S5pmJYJATYOZ
2mLCSAC3RxFsvolSxarrc1DSO/Zr9EpgrN97ZqfJbIyXXGKeUakgTGmaJXtoaCTX9TxDqpIJa9xv
yk0cB9Y9P6O/AstZtkiM8r2v2RDkXZ61U0TOFIbQ/pSJR738LD7zik4KF1rtzJyqtwWzpaTgonnD
4KNYCsM1eV+lzgqpkYc/JVLTVmuyVtrY9PNE6SD1+qYRx5BIEpIduf5geDbQDCZhO1upZPtGvJe3
rwvFrGepztv1R3aAeNGiJQcGQgykajKbeu9CpHIWsPAMVjwHT2+7db++z6rUdmXUeYfwlxpXTSVO
Ttd2MBRSV/+Ld1FYNqyNRTMU+oLczJ6u9OoSBYLCgkBP0opCR8O2Hut7CNRXdvvsBB8xom/+G+wT
/GwjlRJSWHflY/5JWGN8qT+rCdBbcsVDWWjBtuXL1l1rVmd7+f57/ZEdE8tCAEwjRcO26kNsGKXS
XEmwZ/mUDHU5S/Yyd6JfYedGxJK4/m5IPmrQHbH6RrW472Sra7K7f2HloJYM+x2kXE1XkmUv/szD
vpLFXsgDJG5mS9ibgNj6Y6R2/7l3+BET1LStZ4l2rO70Lda4Xuof+SYAs3mc+8SKtVhEnArB5cRT
xB+iwp5apYoCdJYtR7rF75pl2HxE/VxHfK9zsMrzFnHRXHqjFAAvkAfmh5YS8/he4k7l0GNIVumV
0r0GFHGr10UsDNEUr3b7ODkyeS9E02/UnWRTFCLmqbgtjYewbV+3anx2LZoSPt5l3e3K2sffeSB/
3AodYA5sHmf/v6QOfSbBSQb9eF2sMnF3F472fDSiwCmzpYwILaqQDUY2niQN4ENWOZIckAtFeZNy
6YQj5NeO7AXCbIp6gNNxNT4rxvdY/xzmk8rfFHgFYQQW82kQcNn1otGm9SDTlKvGPRvO4RaiUMWi
HlhPvyplUYt+tRQtwGX+hUZWkcF8ND9pW1UcMxwdUaoVA76XIkIYuu2CvWr6sNUP3ISPxKqMJ2cH
xY4U5nH877Upsr4JvkBPMcx3T+MtVn+8vV5Z8pDGx6BiIEBE2+LRArUjW6b2B10MNHsuU1lcSnjB
rS2Gv9EtLdC2al32DFWb/zkqBHqgluT2RtCKmpZGZtrp6ojnGKJ7bOdgiIkbtrOunzwIgJGEbTnb
IN/AOhr5MQjIaCf0RFRQrBnZQqSzPDwsuEd2Y3TcaOcbMqUcg1//oGTILlxSqpy5fJdAX9XHuCg9
w1ua93yryui4agGnWjJPt5iIfqLqxpSA4OpeazrGfBZ5SCaK1RiljY1m7TrJmusw+njvpTsPcyDZ
EXqipKSbldQpY9MTXi8aAIhYqdL+IDe0lAGMHC4JNLz6ct6gbVHo1OCQkVq61OTRt73k2hruZlsd
oDz01Ngg3NWllnFJZU1NMFJiymKePbnucqWsU60UnEduPJE2J1XMdecgsyT91RoxvSEDgEojlrrs
ZNdoKq3yByNiTMBYkJrf+Wy1/Z5THOmlmBe3xv+96Nv9ZUXwqils9HSlMMxoiLmWWYtENKC//l/T
lv0T7Xt+G2bqDbTp6x4zgYhsaU5FniGWECkcLkc9ybkcmHNt+jjt9/90Xrv+sdzfQ9ISDQOWkvim
O3+si6bZo2kq/EdLQpdVzyI8POf65xvg8ZbGKERTl+KqlxJyl9KuXi6sna3ENxGuhdqLap2Bul2I
YtHyPy5U2MU6ek92gNcMgtzYAL1MskZHX+1Q30TvikrOBXCDsVjtcAUNaZnv5l9jWZPAwpTTFe0T
uNTqRHqw3r3lSbTPYoqq7EvtbKxEcLpoyT1yPUrwAP+L4kUszw5fQahR/TRrSPKoKeweqYW3AQx9
bnMMEjFVM3tKdcBJeh72IGqg/uSI4PpB4MK1MaHfVtfUJdNwffNSVw0iMMitpZRlid+cyKsBKX0b
fqsbrC4vHUd6XYDcAjZc0cZj0SzoDAECngMPS1JDKNr1WlLSvcPfq4SJ6OQxx+Ih8gCUak+0UZIU
6ywn8w+mnbiVgKDzUz5wuklYlfu0Yqd6LIqMCJKwUKHXomXjA8XYlVZ3/xkI5NUJetnRoUN9ERVH
r2wFTECQKFO8CSba+mRy76bd08kWt3Y7nkympQWFYmhyUJrHgka0I6T6OI7sr6fioqyvzFZPO6gK
IKRVg2zgnRq0CrOxYUGgFqAkSakBw3RxvN21Hu3o3UOyPGDxuWMkJDayAcYz/BMotVhlS8wG3TMy
sI+RnHwHipfSTQVmj3DHNdTvz0tlSkDNfjF7vlaNaD9GUrHvHtB/QHucwBszXsrVimHPPni0vQvv
9R3LKObH0IN6S7uSbbXTuRHsgjnrL8jLWwjzGSutqrrPxHt5OXed9oF1aDrkbMi8RNg/d/uDF/Zf
KMnAx6K0m2HtmW0bfq9L2jcnB8qirMetNHD+Zz52diTGfYtrv6l5lo/WfzWVC1OU5g0Gf7eCAAAj
V6/toJatFFCIzlUeFs0nhEpDiHXhN9M5oBnWbhl4gUNz0+GE278B3wNkdRMmUUkZDSTcr0N/7zL1
aHmWvwctXGUW7BUwGSzwM6QcGFlZIaY81wV+gF0/x93EXrENJyQfTIiI3x4eqp5K25qJTOv+13Nr
Q2/noicSRRWtuEa+X6S3qldRXLmAB0vxLHSQnwaYAnemc8REmNkj75TG08P9dZxoIDvj2Rr5euP3
kI6tU1e+zDlf8ewQoI9PpOB2UPhUjKy7hfBRLtBVYRQU9gsUGmnTPa3F3WXccCi2gaxJ48/IwCFu
CY4nykPK347lJ5TDuu8CMHPxA/qRlMfE7rvKjlsgnRhLVueEQ/2lNw36e9Fk2z3Gr+J4P75krefH
QkZLaVBnvxTRPGisQrN3vUjKBNNnbSBhlyNXkd/6W4TVebm5UOD78qKVw8o1XZGqT5yfoSP54F9I
ndW6r3LhgUBL/d+k6GwbEIcSXQmvoA1PjzTiAQm9WFm+CGn+oBbf4rJa5em/wS4x8GvRkuikqVaB
uYGpWFTfMjr9lbsdOwFv5eoKT80D2KlIiCVMK/xsqn3JLchFagN+ELJsJy/fc0XJqDJwuiLF8Uno
AnS3wzMFWACjEBVIHP2Bt07H2jX/fZkJ6mNjK9PjCBqhPwOawaeI5OYCVP+nbBvd48RDq7bzUpAW
3mbifPNa88A0EeNtug9ebMbD0txGBg/yWRiCaTmJSVm3XlzmCyG5TbeTak9XYybswUqHcfkfckKO
Cj8yWtgqjqMZFNf2YbenWRZo1RSsAd2kWSp4/JFYVdecw2ukXyuQOssS3qY/7gg1Uvd6xjpzULti
JpgeezhFTsOUTLstyL7q6JSfNhRyElHBEOUPdSasVObSnv7Yu6uIiTew3wVqkcInCkLuQxt2V2VL
rxnxoH7kPL0okmwb0hB/foCxKV9WLHPgTOrVf1oVKEelyTwBxUSRTc1SFF45xZ40wTR9BXYy46Lt
vYXsmu+vrJr+5B25KgaMcFanlLC/TMtUAbpGU4p8bwH2W4lYS7buyKIj2RKhYN1ot11eux3faMOr
q7d0vr9qDkJuYml2srx9d7DIYE/+x72xuwhfvQxSPICe2TUq1PFZVM56lGNjB+uZ18nqZTgveZeo
80pj3B6wR7btIsH50+CZUzWLGuP7dA6g2Ob1cYRPvw5EithvYc+/dSED/MQrPhBsk5Ac3xd8CjZN
bXVz9vmY8wFow4qE+8NJA6xUSu9HWaOo3aUq9E/H5/r4tfEjENfKoKcVc5iEcljSJzk/Tx1jIO2R
kWvYikAyJG9b8JlYbnWcq5lcOp27xGh6GjLO0goALEFuxVr43xotHs0N3OkWDXqTrztopzBQCblr
BP4SHDk2yrODdbjZznIh5CrGRdsRat2WsCgupuLbgcmO17vPymPWKt2jFcePStc+2Ji1OLLP04v3
ysIQF5L+9mCAkSkPXxh2KwOGpMPI5Bo5oSVBHi41F83/7Z3PBKtu+l7Sz4A89Ck8MgD6Q/WUyjun
aI5pxaZ9RW/gn5dFa0qm4T+e0GSP4XbCrYbhGwIwDiMwpkverDXi3lxTBAVshnKFvvtjqKvnghkr
4n/nQSXlHwgLHtpGXyvWbWO8yx/F8on3pZR1aySrcXtrOG/jZY+vAYKd+n68/hcEpA19Z9GrxFOe
DOI6bxsm5wkoC+niPAomPIY4SXYdGKPavpvYM+VpF1zbPCVIKpLddmAmwj9uQ0lu9S0CfT+azOnc
tGxk5644gsowtNpaY+qoKKzBjEXyBPfFfdUlM77/jWQYaZ7D3GkZsUowqnSRBnWW3a4V05BEapMZ
BoRAuADWuiPncWS8xUb1LK7n5gyuym8TLjTnAUPA21WF9bsZFAnjqakDJWxtdDfgL2LI9EINkV0G
Yhc3bQLGtBx2WBEZ9fDNqm1CPLpxAN/8XkwmPRlyjn8JjkFW+zk2tdEBNANKztnxSnFRHKqEX+P8
3Azlw4OA1Uc/TUCeAPteDWY1Ymgnnhcd+Z3LKuXo7+k88H1SFwZquOKiviuAwrJ+5EqziljQQIHp
49K39gAeHv2mcXtJjMOqwakmYzxjURNXLdcbmvr25RBQ9xhvCNl0IdsPeUYpMDlh8DY/s6WQuCxI
EDoKe4pfYTbKgaqbU2LlJJ0IMc+FUVyrYnQZz35AMtq6e3ZhrQzy049SmDTeeSvYjmx1HouItv5q
qlmHCqYCdtsDOy1bO/gcn0FhImhPyQigVkeXbzfkOy3cCziMeTT81in7wKQgilLXe2BSuV3rakmk
EUFr2AZFHejtwbnoS7+n++B8wkBB3urpCPb3woHUAVj/M0ap3yAETTgEmD+sTqjCqyxWKYYYDY1z
BMfBGIZQngy4jWpz+NYZ+KBOjVk0OUPhWGMm6zCqQrzdtITgBBsar+a6M7MeycgNF1e26Z3FJ7iq
PwKXFIj8uxHeOrnwchMhPDV3H30/17liOsmUArYHvdhC0k/bb9SdDaSuMJQLq/KT+Ezl65w5hRds
65o7GX6OUe294p5GVrPdm/IWuqHP1zLeUViEnbHr3stb72FoF3TArawOMIHERaDlduXxuAiww+ME
lYL7bu44VumGpJoL4hcXBgsnQpC3m90yUuSKpkm5BazV0srO2rhqTzSuK1K2hhGcmYsD6mMHeQA/
Ahh1keKtPhJsHco5Z8iIZ5NYgZUqLK+W53SKFMvYuoON8zuN94cGNuEn53n2rISXOLsRYrUBDDSw
QiCiyYC2Wyy4HulfLySR9F5FRGUPaBk8AXVaT0mkn3PyiD5NKM4trv6FtCQESujx6liMPPga5DDa
WMloXGJWPnyNqReAyDaaosv2aXDjYxTLsuZdAc7Qg+KXCa4RhE8oUKzExv17lADOJcJR/9HKf3c9
flo99LZMAlYD1rrdakD8Z+jlidVW6EFVKGskyyAu+wF54wRnnfQEEpZONIH5EFMR0PEs+fJrtqI7
KH58+wy4PKewJXQoyoLAPETAiiWnq+qiOldFQHIQ/n1pf22umtqb2E/kAV+7vCrNzOP9sLzLLEiC
JmPBxwjql1f1Fy8VO2KH+StZYBZcv8EqlOplt56uIhh7a3+BkNZVrVuIfto9fKIYz/fyQa5DuTFT
l2DpiwmS0bNkP5NMKVzXehgrdh/Nov1ivwbzOht8S3nTp+qN9zMfbEtVqHL36VdCwVaYvU1O2hmB
IOOh8AjMush9L5Wse9VnIldBu/SNFVFY+Z99n+DEo6v+7qyvB0NmjDe3Po9k0nwvrtXgEL2/ueCP
NFEQ9wjexFJTDoj00PplW/D9S6k2bOfGVtHPxXrFZMzgvssjWGs/BSK9UAeoRU+7bN1VtZelo36X
Kg89gyRekycRwcq69qKm9bHLv24ZUu5h4ZDifAiBwNIrVs8ZCJd/XOxxFf/FQf7IOeQJNYyx214i
oLFh92VwYmqbfU5fs4iDDbmeW4Z3jxfA+BZut81szxXOn9TX5sWT5Ci5rfI1WzVbnGSAKsCrhnwJ
/kk8ip1evya1yByyGLB4fhhBebai7CWLMK8biBPyAebKgP4I2ws0WOVh0PcEybTqS2TLdtpn1k3G
i76XOXr/4QI5Z75jzeLFneMN6FEbVKRWEyDMrVRXwMiYe9FMmeR99Q3W0iTZsp5NcVmOWAWeeppF
y8tEegQljWh0V511gCvu/REH5MF+E+j8OFRrmvthPJLPm61JUoAbsrgSSlUlkZOEEXfWFECgM5Hr
toh8mhymOhgOef6Oy+igrKZ/ztbmFoCV7VjcyoMdmDagL9sMLV/C+rPEAZdvf6cHsJffuDdEy+1j
ePjkmyKZ54OBeraefJG9GhZsPCRe6JOuqmXWquvDJMBlG/rgIQ6OSkVWV52gX/SW7hGXYCSASaXr
BtWo53H74TL9h5F0wF6z0oXRe1rCmruGOGtZFqLNlVA7Z+Q1peFR+TV0wSI6ifnJhDZ6+dyUswaH
jcOrEJvTKE4pftWt8zuttqCswI8+vIWoVo6KL1Giz/PP9dFBsmpZve+ya/YSYk7ATLP/CVfHScMs
0qxziVk45epg+n1PvB9TzDQ/n+XgvoUdlrerT76kwk8GIxdxkZ/6xRBMGAfvbSRZ16TTvQcJ5K1H
XtiLM7crPYFHorAMeLQiI0hNRYSN2O09KKgnE/XkQ3NLwMEaOvZ0YGHsR51ZXtYw9Yrhk4166k+G
pg1g4kAqtINnT0PM34cZhoKiYf6PkHCWd5C+9J4487QQs3ZbtseGNn1aKtGjuQVZtg7L4YfJqlGD
Xai5dOiG5AcX6ky+EQ3k+BNz7M2btRDungOr/pd/IsCX8EcCGhohBidgkW6mWxoJDlTwANBeCsyy
Hcn1qN9CoPH0hE3PoRTbyCS4PgSeeuR3zhzffcqIN0yoJH9akJLUaPAFgYiuCu9mDy8LsufmByhr
8VWPO3EbqKCiWalb5tbKgzJaazTomONqWnQGJDHUenIiXgV54S+cIR6u+I4j2WUdgXYKcmBx/6yl
V7zbNGzDTB83/m/OXoUGgodpP2buk6NMqbdfFLFPSmIaxAm/KqZTaCaiY6PEHB12qyZNM4uBZtOk
bvERd8K+LyQskGTKX1SWtXhGQvrCw8jh+tF0mOvkEgk2aDgama13bpujXMibMUUl70CKfwU2lMvM
/AeQjXDAZQr7BaMtuAt3n9OEG9auB+P9yAbaz/lE/dFU5r5Kiw06biOYhN2Zsvfjox4KD7Nm3gCc
P5ggdAY9rf3suSo3pM3hirYZrcb4fPBgnePLZ1i8lo8P9AwZ/X7zLyMoQZ4JvJ1sgTjbM+BijwlT
dmqo6Ff/PjFFozrPJXhMTW7J8B+dhFebpn3HuNaIlXz1u1nr+FlGcfe0IdeNcOSJRjkUm3yiYm1s
nWKxDIbynQuu9frkBXXevDLbhJzlzq8Sn/nnBZbKsGYxMR2jwgbn+3uBQAJooBTXaekWKESDC3tk
GUkzjbZ4PeodkwxyIkQdBdR2NGdjcxW1R7ayvi2Pg61Sm15HQqreIsbpnLmqLJhzPpG1yOWHG/rJ
baPvPsAQYwZ5WpQhSpt0CFUyOYU5ghPFLDJd+RZFnxltLb0mBKH1P+MThahlzHqTZrnNU2i3eP3b
yBOTdIL8WZdlqpgR0ZV/+B5JFPW/5/31g+Pz0ifWSA+erbi31vH4VIRQrPZbLTCPqS7FF3WJ/ok3
IT9d/rHYrdI5y/id4rLKWgQAYplEP/SItBa/8T+1NgRVAnaJjqhtAhE4npz0RSP68WuQ6XfaNnQr
LyGmPste2LfXacSU9GS8HYMyb33l7kTe09Z8GnMcEF7sk2Hg8rCTo6ZLpbN8xQ7spZDxsvbz3CYv
oGiV+IXZqF2/zo7IlnBG4Wrpoi6kN3g9A3MRO4EcI742Yi+0JaNPGvGniMnyuM6wtT+uYi60DT4G
NBECozqX34qNmskXulN413SnzoGoQgKobU9MSBTzNFxKHZ65Ha6MvP4yChb7YRwqTGOiPMkI8WA7
v+Z1cMb71PkU/yisLU1O/6rl76Bcga3WGCpAB59vUgQ3DWD5sg3Kpk6UVDoDQ2cuU84ORqduYCv5
Nj89+GezGlHQDgw/VzE7aDdcd2HNuyVuU/QWUBjYbKwUYxcZY/7iOw2jXZr3tFWCnDdLyddwh534
fnjmtkg3ekO/98DR5Ymsg4xqc/FcSnPU3XrZwdgLm1OiUZtmsnNvCmvYjFON4+vo6p4nq4KPtSiA
jaQYLRvZmhi4+uI4eP0vh4bvGW0FIQXEvUnJ1iEFedV1yTXsXfmfWxAOOiMhbdEy+uo39XCA++id
5hMbx4sBTaGfOxL/mo5Bbsr6hONKhSPUfvTnJ8zCFRfE5zz4hIRV+JeolU+X3QPumC+kNKOwA25h
rM5ESRgyGUUJOtwpAP7drG9Z9uueE5tGSamhVlnupC6RHue0StClPLcyOE/w8Psk1nv+52Ixw2xs
L8LzgxAGJsVjAx/EQhZd1qdZ4srRegniipxvMREY+OOdJD1fu4SN5spK/8P1Xn4HgWVxcAZ8Wq30
vMZwOEWEpRXTN7yq5r1QslRZKtc9bSm4KPZ3/+I0PzrOBpMmYRPVDgr4Y8bz0BUtY3WqYG1UNjpe
oCb6RBJ2M+jCgTfNe26rV7o4G83kdFOg8mfn1A0gL9d2zzMLOzPtZNlf23kJNMfDCxHtcWXfKETg
etHRQgx8nw98qz/wweirBNweopPHSfwb21XnaVzIXyMy4lMXGIM3DiVdl4LE8xUElF6QCFrQvvkj
STnZxjA/oS3BwOcKZD65ofYlIek+BU4lUYHjcybwYbESIK379NJkqYOO5w/mRt9Rczy22NXVjg5Y
uJ22ia9b+MqK0LNix/NBPxuKPzS1a10zP47H1M30FEUHuIWqor6ZUbn9DQkRz9no0G1XJ5i468Aw
XkxRxdKbJ1CNMDrGFNCz1fw9xwDzArhqfRmI38roVYHNJy5zyRfnj66hoWDt1oOGxCuQAMUjl0JH
KiCGlREzpyW7roxYMHtSpBY2F+Mv59aOnfvZz7P6cv7xzrB3fMTkixKlNS8xklyqeuUFLXJbVNnk
iMtzklnShepE9CsCnTYP6VKA9xa2xkKXsu+C2IaWm0GgtGuH58jlMlxNliI0lJZ8LSrQvrkXL24W
YKRJZujmXdSeU3Fjz5BTMwV8PiVhCYR8tWBZDEw/R8wpK6+DQu8mWNlbllVPAvonHw1/Qw+Gl2dk
Fkwt/Gb48meO6i78GryCggLJ9KbaPhnfEg1cD3n3X37Jewk+UFY4hVbZu+bJAJbaY+LFdyTjWN7H
/OMSg1ib/8fnfVuobDhUhrDF+loR4FJ529JQFoa6kIuo+FfgKbLnMZLfJnjL5c2yVGie8dAKr/Kc
piHeKK/QupY4WBWR8MBOws4Qd4lnISF5zKeuQSE9BvttOKL8cGkUO+ttkBRDYmJkBWTW6lzcZpoY
grZrH24YgGvZac472ayCskhEQXXz5epy8qiUWxjazdTs9o06RzsB4nvFsmCL8sc9dYAg3PvrTdNg
MxzMHw1LbkkFqqJTqmkR4cAd8If+pWD+QQMh7wPKf2Bh8/i1TLrlM2GSZ2fip1BiMFwLXAVbadFp
JEasDOkLmX2W6W2gnxQn8p2U1CcXy51nbpNzO3FRcvSgOdP6mR3W5YEiyVXUtiBuLrd+MKsDI0SQ
zX1oCV09OeY9v8GzwIIooGUIIN04JR0RgNmnm+79sD28TbvefPj/LeYtp+PpGrTSNUKEGy/aRSeW
mJdN+JfldZHQuLkJ83n9FBJCC9emmPnq8dxnbisBcdVSTRrHWeJ++80A3KUD1JV7SNYKhLmrN44x
ck4m6AUoKIPisHOnYbjMBHZCqT6PJoOedWYFsj+avuvZ/WqneUGP37LiesgUNfFS5erXxNfjdzKS
faVn9oL2MFyYQnyhLHcOT1tP2LCNlxlrLvH6EmLGR8sR0aF1J5WVf1/dHPylnO9PDNO5QO3mUeZ+
SDJ5Rqm0I3SkcV0uhQ32Hv+sNEHTSslUtGX1KiQAgEQr2gGmZR1fMly8ild/wikvhYclftKvYB2b
swS6Lgzpf1d9Rwfn9yamGUmzU0TZD3MCKqRRW0qGwO2rPxSrVHL5qU5Gzmrl3TsILZCsREEUI2Ln
Rd47ML/d+bNH20n+KhMipLva5tIjdfnudMIJMptLTYDhrhS5tdRb8vkytQLf7KSS/dmCofHCDA2+
wb7SFfqOTgegA+6ITbiUbjOntbzUM/8DGLwZlfS2ckmG7JKM0cJRjUjIui41qGaCnoCNXg4Wg/1n
htstvgqslyObP7woWUH/pWe03Mn16KEWULrjuQDWcUR2VW1mUosJ0IGVe2nn4NmhCzz31nDAK2ml
Tuvab4i1JSauT6KlX0U3EhDMcFWxbLcyxDp8lMvF6KyjskA0XDML++1gz0ACMSOFJVRVh7cBCLI4
PSPuPOASZCIzqdavS+j5nbapN+ix1VEMMPbP+9xhgIaBKPFD97HW9nKaE2y+yvlviMIIQUqSgTvp
+TAfezv6zTPQ09bNcLTzMv/K5We/jwYJcuSC6K1VTJynuP4fVi1J9gqduuR5VUv5teK7ExHnTVEF
ojkoBSpHqd/JD+XWq4jdKXghTriMlGM52lbx9MrrIcGGeEHPXpFKFKz4mwU7C7FTjB2Ch2V+26wM
QUlxoHNcEao1Tpi4YDa1CKAt3iMOB2/nKN5OmZdYAqIZT3OdL381JM5iIHrmGQJeVHDslT+aRofj
Pj09sOoKwCypDn/5QD8jK1AsSutcLulJZgvsWLKj+jbt/I+f1zmGmZK1FFTF5EezNesNgErY3kkf
j0NlkgZR8puZW1GjEgKEuwLyJ8w2RIvgrjLDplvRyb23HEzlGYzbflTbUCElDzkV/SgEMLuEjp43
DTcnWvBDzKb9a/H64ETDx3Ub7FEXO0t/3G+7JPeH1TJSR9+kVBW8qpNjVTI7z5B4ixfdrfmkwspP
ytK5Uuv7iHZin4hWXQVWixCZVAGguzdu24lRwBS0pe0oaPxPIYF47+PKIvZRSdmoEcZJE8x/6p14
fgnhYDv6AhE1isT7ethGCpA+Jf4xOODNxbjOSasxA1gIV2TwFowW4Y0EShkJ8h+GPMBrfjqOPCx/
x/WHraYKmIk0fcqRYWoATICydOll+qOaAjgLSJbmsJmyrLGEDW6WaVhxbboUrH4qmQtJyRZ2KibW
/Us9LQAdQoLFMp7GFSWX+EvngPf6j+/ZP96Yh0mk2cnMMBEzBy3Mi+YnxxuQI5yftUp2WhEH+2o0
LMJiHOiLes3BIFKQEy9oZqXEWIvtvtnuCs73qnQf53l0EDX4uQq2Or6u8HiIZ4UuKIaKakIgEwMD
xtr8x7gfQdPf01VL9jefnKr1k+1mSsb6EeuXkjWnrwqqEQklCCIOms4vnzMB2R7OCVJTjkuh4AQ5
JkrjOinkgDXa16LB+HKSTx1U1hZE2a64T35FckIe4fYaf7/XWDD6KrrmqXXtZ22lPIN5n6Xso3Ut
rwAaK2OMv4Q+amSxUyEQkZ/9VNqSpR4q5JYjunV7Af1JX5E8ENtAv9HhLXtofmjSWhuSIKsTKAAN
Ht+UzcbnBtcGT18IB+fLdPy73voXzSdAS165tG/zMlvK3UPxd7qfEReDwmDD9VMMCbdUV8vPXh12
elp2HXEZ6u9qajIsst7rPm6BiQIoSsLfzVEPjMtvzsfClMZkgu5o2TEH1FK3w8HRm0agzbEkECEm
iwcClimN1kR2oN+UDL7ez7KoqEv0FAQQDoOEVUpKyoNKvaF/GldNvAL87aLa0FLkITh1QJVbCkPH
hNRzrGIkHyG0wpW6dAblDRAw3P/a7rVsrtfuQ7PeSxqimR6oOq+WUuYpQKqyHZOthnplmJzSisar
WGg7FhxZrBY6bbwMRvZx1rY6Awmbto8Qbilb13vKrmrzoPKMWHQ3fqCtG4gTm9K8AWT4j0tJklU5
Rxh/OzXBwLptCmvbdXjv5GlrFzeQ9kylyJ1w7/7rIlZQs1RBoLeoOIJB6dm7R12EhV6mTszFnYks
8xeDpJhY+7Ne3ATj3HABLt7hPi/TaCpNxRBXseTegZ9P52WTCAm48ef4kxeP6SmHyaPMm6TX8TZT
ttcVHv5ybQd4T34TEyO09K8J2zcagNGndscbhqy2iCLMTf+o3JRlZ5dvgrfRxF3lrSWuw1D4EKHz
Aaw3uby5/60xutWICZvUnaxM7QWTNmeYpoJL/LziR3VaxRhiGXRpad/vVDRibDqarO4NGwou6UKF
rQtYj4NzO84UG/ajDJBP2qXpndoCvJW37FDPaH/+KlpMKimJnUR6y2+Fr0qvSSfpB/fyj8S1xMv/
d88utCJktWjT946nNi/5WSnifcZT4xn9PdrWvHOm3H7k6Gfz+YiPALmJAHEq2Jh8qWJoNY1lBj6t
OtecAZneva2/GoWW+BlplX73x6qwDXq25AD/UfB3i9DACWdyaBnnW708frLWQJxfbLV+WmCrLWl0
sdz/6dRohAylwESwwf7+zQVn25qeUgdspS791AdKhNe9siMO8bLnxnmkk5dQ3QCpkLMUAMdMfGU3
3B387OQPaD0Fba7va4ZxgSeD8wvVeVTRqof1iiWHAnNLwLCBClfhe+0xnmCpLjrkU/50CeqaUXeP
jAbVUkeoc8Uidlv31Cvk/1RfWuUZBTbjknBQmOAx27WiYS56AaCPEf1pAm/YWLC7Dw6uqqG5vAsM
Mw0po399Uj4Pki60vxAD7H+5hGmDI5dbSR0qR+i43N8L8RpenA/9g8kWXhugZs+o8NUc0xpaXSpk
ojN7uKAsNCOKTmSW3PE6jnvveK6laB4n2/YRusvLwFOFlvuYdlz/A9Ph+isFGBIQoJhz7oxIXQCN
YsTICqWDmqbjE3m/3M3fVfmjX3Q5RK/FIgAF7khnCeYHEo7oS1oNJzQ9CHSUKDpOs/aOA5qqZ205
VjXd6Ok5EmT3LeoRd8Xd76fIzuCULO6sa/S3pEX8U0g5W9vZmZ+PfOZBFDeXYbb7H2wOqG2B/H3u
ATuqz0hOfVUXm1iOmkB58S3gV8huoGYpcBbWyNojSXza8SZ5aSN9qJDbnANVGK7X0f1PL/zTNNnh
rvlWDcWMNFa2brOu/AIGpMOcPfPVR9zrzFS0I7/PGBBGgjntLNy7s1eVmMz9K1z19eVsvCmkcmS5
zEr2kSctX7NzC9rxtyM7qTUVDnx2VrEbyKv4s/7PNiIIBo6tfC6sW04NaROIgFI66x1UA0ioSrXD
CQ4sB/gyoDiSfDHS+DwAVoeYtNpJAnkDFiqdxsKHAPFt9GKHnJ7g9Vpag1iYazTt8Eu+qQm39qFj
CDz3eqHkJJwfZ3xv+KB3topUdznkh5ikzw15Oie8uxtLh8MnEbZRPf9cazuFfwZ/mwYcpUfHB9cR
6QxpnvH0DkBDz6gxlRwCBcbFmNoXXkbqi1c69JZrfPqsf6UPfIQgfkeztel+wQZ/6JS3j0QQvJvm
k5pw6x8jV1MI85ZC1SXAHstZumBMOBDOGtWwXpjOOSubYAqS1Ka1ybAVBhXzZhoLUVP9+Vhq4K/M
bSGxV43RbUoEs36WEDQqOlA8+S96Fxp6V4vYeD+n14EaEQXJAQ/NcIa2GKIqdVBmM/CUTNeCuvHc
IUKBHPjM++UIhH7jbiE9LYxM3z04hQCgtPdYYxITeF33zUAM+lZkjGCDx0nLLz+gJIPWRaI6rrWX
6QVBPByKqi+EnBZ+QXhTwLy05MG4wg7ZuLXzDYwEsvabjz5JMjO+hy0whq+CMuB86xhQhlyOtW4l
iMVYW7XGuoIBDcotly5mXVNlfw8A+jCX5q7Eyic0HYyyWmmTaLLkrREAwoa1ZYiofiWcHfkIORs+
eUkRfU5BD1jrXYsKRgwIgt6iK21IS0UMcGFafXJ3TocDVgJNdfEDpJ2+/+JNd7Bmcxm5ImMNDtfz
saLYH7P5YgpFGcUrSoKvx/ozQRT0vwwLmPZXCdXlPr9Ob9VLym0Un2iAP+BIGwmUDOLlCmD22Z4h
skfeMgDu8C2rfLjXHswaR1vAnjozDipRrH9l4JceEZRM4mwoNSOch8KQJ8085KNzdSkXfImPN7uo
ZU/xAnTMBj5iGJyi7NzcRoenGQtACZuCkmkvuLS/PcJfO0zLmKP95uYDQPDgiRf69LyQ2sIf7elW
IDig6c35MrzBAvpAoi7+p4+ZpU1AuyJt5kHoXcESAtk2i6pCD85n1BsXdFKs8Wc5PXKI2Ihnli8K
Pm8uOlWkeX4XdqHK2LG0g/QvX+wXW5Q2pEZsV3jKIMyRW25XQiHdqu0Xtj63lMJkadbq3dtF/HBY
o5cPQe1nPYXLuAgktwFsoJojO+ZsTqM/iB6S3kDTSE+fYWeJSKExz0nXtKYxFG2gia6MMuTIkuDE
JQvHuZa2+K/LgdRRWfXjOPMvw/pp6mOw/+/45cY9b0ZWvs+MtlG9aCvUiZtXwYF+3EXNd6TtMqln
5v6GNix6xNB7MKcGhNOcoqw5HoK5LCZOLJeNGb2yvrUEY4vwAN9gO5FQ75nNSfI1B0J96RDVfA2l
I+TOIa8WxtwB0FgbH0+RYnN6C/e569t07CKbE2MEbY7n3nw5O2CpMy0WEFAF/RrtDBaehUv5huQc
MCoxx1NnPcrO6FYbpS8hCo04IB/eKrTpsgu12iluNj0yicyU+vIHKsCxPsOo4TqA7/tX6uKGGsQA
DPO3w86SsicyT0ODSjuecoxaXPazoXRGnGr9j5faKot3J23LJESesAd8l5zlspMvh3jDjauDteXe
/mUHH8rOXB/Cm0JAmR9QitsDFgZQUdPOrL9jUckipLYoR6Up5gLtkY1Mfe1fb0TLd0l2moh/2yHn
TDF0Kl8Z1oy/BK2enAT9afH+F0Q5a0BEq5MimSvto0qh184kf0xbPtLm+W5WS95KxJlumSvXpbrG
nlM17uD8h0mgrBO9YQPIlrf3vzDHQNJzq7TARm3+BKwTmn1/QX/MeDhh2eXmZardQ069ARc23JVX
afvaaM3LPqVEYo9AI08CARvrStMYQb+NYpNnaHK8QuEmY21e0gREXSRdCpHrApmE1hvL3rQC2g8S
OsPJa7+P704delVBgi/cAUFRcwn3FLH+VQfflI5bKQ/pYuZHp90IbkunaJjdlEqxjTkhUDOjGZBI
VHz3MVmD9X2oAdxO4XdtsmnxL4+rwjaefTc8+yfiSEhlDM6XPUoGkJRlRoI6525yl9+zu1OdCQab
aX/nRUoSsvYYcGWMwegSthXDrhq40HXeLihRqjmEFAhMGyopL0hkhLTOE6YsIMMnFQv8KZ8bFqvI
BiUHzAwWWX3HlayClZq6OE0oMgAvLs5OlJRzuyllCHGKLCvkOtiO/3NgKRK5zcy5Tst0ZFWURGs1
Pp/2iAXqMhF9VWYlw3nzrEUEzLxMORxrnHLZaWeY6zH/zJhRRGlJT7yufPqa//iSiH+muW+Hs/Yp
7MecCDRwx3+xEyDySLifcT0KzmL1Z0z0ihgXOkwpKhNuWSi8c7jQHPHfH9Ue0vOcP38+amtBu5WS
0+cYVOEiugMNT7yin9etrwfIOXmIcNAZ1+LPSlM/n70DM7UwpiinvHKiah4Y5TUVDR2mteTBXFZQ
2QxDO4pVxSwWbRjFJOc7OK2//u0pbXUPbVdXt+0pS1CAzSRg/iMeAsVCO/05ULgsAuMxmlXgFrbg
Kr4ORr8lQ00dMLQ/Y9pI3KJlvT58vDsSMrvXkG+QWzLWNSzDFlvgNPT2HI/bKbVjj8I1mR/QJmJN
2VEXoanZWh8Yh8heogbbrABUYL4RlaypNvrpvudhUnKJlPl2xNTDV9waCE4xEX+nIFoohiFJqL+y
Dcxe4JgHlksa682u8ky4k28WsqnM3IUo5toTlvBo/QvnudevZCFEg9kuD5Z5uOIr4lC2YpU1zT+K
pSXTydW/N65tk9uORFGrZqiGstUcHITxn95+Zw/VRiSSAzcIZJhTEbMZAGMYlq/QsmFlkwiDy6P4
/Jz06Ian1ml3cEdwtYzjxmBWljrIrLFLugbXIbVTafkj2XnoXXHDwJYqQ/rYkr7WhssBzuO/uukE
h11qNUmPqGvQe4ErYxx6pf58Jb1a+T8AoB4uXl9sEbQGHvZumNbwYP9tuVnuzQ9p/oxUDLyqw9+V
3JGZVOLBwQtocbYqxSw8qXoiA9WonFGjyejpckxvxVxfwWqCH0iuS+iN41dsOiE/dQAIbt8jzbix
z+aHk70b57jTgJzhU6eArTOGH6DNn+3c+8ZjdzlmZ7lQ7gn7cRHJBPKR4Z1qf2hRKE6vzcZppasy
CvLr8aPUZUdvdorj4o1ZRzbRt87jKOVh4ap4GW3H1yYLAj8IYI1dPRo+kxWVMnP6So76jaAnjYkO
MiBDGi36xWdXS2KXN/v2wdk8CUxW20DJxEhgqIWFzY+cmmdOC1f3R7kEGS7DiSrXyTwjcmF1NoDk
729/YN4BlyWicUxmGtovh9m+6qCzWGK2bMg1JJ+OZzyT/bKLvpg5sLCqCt7pUkTj5asAsAVSKBzN
lmL9wn42+qE397YyedI/idia22RjZThQ1m8wuIdPthLpmTgyv6abMDd/MLqi3ZiucyErsHcfJYQT
AeenspOJGnd1u3HyslHUrgrD/B/k50kzFPm2SxyUBRaTsLIv9PV7RFUjb0bdpmsvPHXl2VzfT5Jx
43nSrdLVRlIyV5sN84GzuZ9vMu77EwkIKlttoM34CPXsRWRnakEF6kWlR8XGy0GqJt7reJeEqyr/
dkSzD1V1EGE33Y5WDfHaSu+oN0eCXbpSIU+IZemirtTMckh7/JoY8+X4jWeyVkLa80FOQaXqTtOK
A8S30Ll7iUktEQ6JyL52a5oFs2Lf/cJ29WmVKSe0WboewhRUDiCNBnoBl5PM3y98ooOaCNRc5Qtg
pJMb8IrwLXqJlzOTNoFHjS9pHlHXsWQ1ow5r1+8MD9UCvc4Pz6zTWBjhxiQuAji0kqTDQceBJaTP
h4uJfQt3nDUdLWRnIwFodp5EtKPI2cQPfUc3UKxvansFXvMDaLB8vy+9/CsO+VV7tA1Tg5KLx23i
ZV1E/OyQWlPPRM/Ta1Pmc7EVQdmAz1Q3+perQdsX8WJSahvQ1ymwVWSaU1x+JdBJhDQMXYCLpqgp
3hbrPGRMn1akm3/OAj5cgQB7+1y2NQ6rASwwgSTDKzmPawrkdS4EE42I7Y6u0j9vKcnl3jF3tw5O
gJdqd/cCjgoPRbUuogHf4lEZf92CRIRiQcNM1kFQDFRuK0rUPog47hPDwS0TqsPq6XG++PnI4/5l
YrxY++7/F5wbpWoYtQj4wAViTb3yDZjlLQzWTOGIga3RhV9Ke8HiFg193TJa+r7D/ST6V+1Uz9q0
PT5dacMIrSgtovQ/+0+wJZDRWBi3lh4XAfW5w88JD90Qb00sVoSslLwbe5vAMDFGgl6w0b9EF0zE
pW9csm/CGzgP0j+j/XWrlRxBG0sr4eKYQ60Tpu6HejJl/J8i1YElcRUVVsfuOJQpFiBEdSpc+JhC
TpVsWoUlZzZGwoRD+5NrGEwcCUNyAABdG1Zs2VlQQRXCt8CXeXolDBLaJqRWtnwheMvJOdL71tDk
5QrM77QdmD1HMiOUBAd7YtXT4dC5/0jnTgkHRIAdqhOhFGrd8S9f9MVfAgwpdHv2G2x00ZTc0ZRn
m+1Be5fFmkg6kxcXR6RkkPYiGjN8uaFDzh68hdQfltYvTIMAu68A89k+Q0kLA/Y3mN+crvuzp2W+
cXumJWU5BctnD5tJjX2OdlfC2J34rrSPRu4CyqAZGbGh32FnJ1idV2Sh3SUoaCi8PCeHCFC427qv
0BqMxEfSVcI/qFd4KmqGZ0HrMRk7jXhFPA4Mig/eGysSY/hDHIOAK9X/uy84Bvu/NzvYZPlrw5Y2
saqoxZy1rxrPmePjxFvRthekcgbPYEubjA8q/q0AHvt+144Kr96NmGuGx7qWTuhzRMdg/XExZQyU
3tXeKII0eiveO3lu2Vbxdi1YNdYJuC8AhTtiokXdyXspHRUt/xev4574YIDd3b4N+rlNM2ed/rEI
HS3n4BbYUwwIkdW+twdXGcJIw5hiZLUwPNMNtom/UICKxB//UbE+UjbPzQw5jdBtisGESiwUZ4Ov
sqDsS9is5mu+XwDIaRoRWEg/EndVUNqEHx+sF2mNmgThyugee05kZFk+skHj+eQMuD9Dp3jUC3Lz
1arikDBTGL1/4NzQu4b0klLLMDWhyrKUzS12h0gVDAbcN8XDUz9BJQpVJrbKpFjWn3/IeEuM20DC
OTyHSl1FbUkKdYJKj3uAETJ8nutCW1JRx3q8nx+b1p+6zt5a2rWhf5zOFaEgzqfCHGnz95b2Q1mr
pOKzlxx95Id631pfx+WjBNLmqO9XGUFsLfr8D4R3OzhQyCsEOAq5jVDHWu8myp8u+STfICuERUcd
EvX/GLbxzkHK//PLfxrIkHW5QBLySbDk+1QqvSIcw66BhRUVTnXiSK4phZntMETl5ZJM3j1szF6S
UTISYgXmEDXlmG0oqiDUUoMHXxR4Qn/ovzDCkZAMt40+6PuSTLeIWquhq1O4UNgue5Erh2qps1RC
NqU+oVD6Gm+c03gfw3J2NgRE7IB460SJujojPD7IWx2BFTtBOTGKOn8XFgRiSrrctKbuAQVxNyke
2bG3/TAJGHXi3HFlfFseHLcakOfcAKo31XWDfPM7s5OzYZsTFicDuDatgks3TdBuMSeOv4mYQJ/K
2mktMwEvWqT7On2iYPYX8MS1qFBgsihPbv1OvWik9ptpR2S42HOLRW33Ri1Zkf02Mn1id+QSE+so
zNZlGHEo+YI2Ke2xwmM1HXuLQYPJay+P3juzwOApkgFjecnob2dvKWFCSAVMSizPBXbqyK+nk86v
iiuDAwsbU2Hiyop5OfMxBHq8JTz7T5gKk7UM3osrl7yyglRCUBMSTMDQn/maOAn0SJ9b6v0+HU6R
leSKkUXHnXH9SguihxRo+p76PLqqAaUfUBrNBXE+FOFQB+cDVsm+tdnaWK9MdbP3ZEJntgkIh1kZ
pMAPIr/4wTmw/RareWAjLcgwLf+tapZNWElbS0uynUwotPQADOjdIYYs2S+0NkBXyjjlewdP0IlK
uoyUjnzM9SI/bRJWxpbKPHOJgNawJdhfoyZLapOk60GKn8XVSqEEq3+N70ncFG6PEQf/1rhi+bA7
3tSnMRIj3L3UZb5fgR1MbqUxIi+DLDnBQhO+Nhc5eN7s9P39b8sENTOmal5sTai+pyTbcyhCssZK
9aorsOybIykFcDrcH3jhRe81h6raHp3Ku0i1JPyOKAPHq2aaeCe6U5qYqJtIiKOtky78KeD6agft
BDRJ25QmCmt6MrLzTwYMSgBKd9O3SUSXRKx3AT4nlh7bji8p7gLe5wJWC90WB3IA6xU51JevPREH
E1V89wlavDqGlsv1jzifCPmRjmhawvkFJwC+5Y8xDYGWZrDZkiiYZzFVFoPIzRXotDoeLlGiEGXI
57UlFM2pNb+oKcbmAMU8+3/nPymc+44Gy035wUBgNzvMnZYKGX/n+O9JhclD1rfpGRhZ4yOCjMrk
W4Qhhi+ljSb2/bFzVWOyjgItzApSyKoLhA/8B3Wn2PP+qSpcpwZ9EcrOSl5seavCdwB7+RagDffP
9ljOQLawPMoMFHAa/KcRqlntSZYNKaEVqwripLXwZ41nZVf2b1gng28talPo3RK7+38bBdfVoyRa
H8DsF/6R1K48XCevWLhq86HT7bLUn4UHJioJsAPaSGbhz2/4I1t2AE8jukLld/Uh9bZmzGQvenu4
J+0lkwlmBcEwCXBnATQ+rL1ZY6e3XkamnpNqgniUwO3hkQOAYrYyLwdGbOz69wxMewwz5vuTooB1
FZQQfnUMlG3nTTY3vWfsnCCJJ6tJ7MycLSB1xmmYfW7nszxKwI0eZqmugfRmgGcPf09siPwnN/SP
KZxaua7Vitq1wPy7vLQBavtYwy+CvkMyP930JnQSSIFo2zbFrlGUHC6GmPekh33rp1cvcQGjY+7y
IAqQ3/UAeEaIX0LmMRLI3+3ofhttlbsBSoNUyZ2WSKLPP4K9UBVxl+paP7tZseZIK9gVHq51MXCN
CZFOQhNw8+rM8vIuYDJW0cXbmBdjm1dQTVmK3u+evl0kh0kPeUoAxLzNeWwuBk1SDUVPZGtKP2TL
VhxYBzK0wNSaSdyq6YkRt98Aejm7UkMVOTdg9OHi2sIczESLWk/oMnLmd048jAWmyI6c/hylAbCw
Lj2j7wCElzflUtHeHFtBn0i/XmDFzcGMoJeNBdx8QkT6dTmid0adFDxWhyxg5qmotUGI0oJ2792L
iBwLde20qpKz2RA87Coplkgu6zPf4V+fBa7kfZvlvhJvuSjuBmWmjH/O+fBRPornQoWniCT376do
kbeuW1aCgVARB18kWwIHx5IW3rbxLBfCX4nLJQW1iqTZJ1mlFskh5TO7oLPcH41l2GQV2msffQbu
LLLO2Zf1Eqkm1IJ3HVqkfzSUMIdWnpgBUYRnD2sGJ7AQnbutxFjVbk+2mMwvNyO4Hfra8hguUABS
Jgu59bdLgRrw0rtxFHlzY5UmUmGGTdm8iH+qurebKTZlBbzXwH0ReXZlm6+DAwQFg7Ss3TnjKxHd
K/8XeVDOUoU/YwMBXAeQQmiiJ/cIaB5yvwbqNhHN6i1YmjDcnsCeK8vgT+fT8GP9wVkx18OHNkgL
rBWZ/Ki78pwk6hiteRX37n7MiC0+7KEnIVWPsxefat6bcvhBK/cI4qcQ+rc9tjm+Jz1LcgwJSxW+
vviuVKTstPX0O4MhdxCOS3B9MudLJjMoew3MwjO1wpf4VpgGLO44ondJUNTf12zMEO0i8pDJ7o4A
TjOGt3BNNvmcfKfm83auCIpOxPtjJ+qRrFRnEpIGUcOJ6ul5Q5qks/2y1FDBDKi2nvINoLH67fhj
7cvxK9Q/6fzNNJ0AEOZ5XQELUr+ME9qqktionZxv4Rj9tdpRcEb5toiDWZliqKRs4kgi+BEocQI9
zrbr1tW+41cCQd4lmPz7DWj6yQ2Xw7coEz+eYCSaJxJBbzvODybtW4CWh+habPD095EzVHcvecNt
uwAC+U+2Vjo+6iq8BSujKET8zgXH7BSpkoZw/a7jJLJZ/DEqHhX7xDGZnG07xxlq0D4Qz3wiYCTz
+pG//2vILHS2jomGn/dubS+giT/EkkEM+54Cd6V9QLPZATGLcxlOaiuL29r3EIXYJqedXSrdTIqb
m75moBcEFTRt+QcE2oCaRRn2nGhfIVYye2uzOXZ31wvdO2A2mqFXJ9cyTVGGmAfXXces99sO5Bxr
EKEehGegUxxJQVFHA55Nso4e0zgRiDjSvt2GowaWKO2A1GnGu09dP8ovEePfT0yn5jAXYe3DtUxi
SUEyPVcLFlTS1uyWGMZHBol4AoNzf98RwzjsLSbiiHEZ9L6Js1t+R1NEYoLEvGL1y4H5A4NIWNMO
I3rxkyLOZTjlHUeCM9ltjqrsYlOOLUdbxek3zSMuWhKoZPREibPKYTBtLmi/hefW2Qi3KW07pnb2
Ecxw1cqGpPSbCZick0gsORm6FwiJHAY3qqX6AFQCiCbZSXcTAR/+kHdAVIhrR7/m0j/YfDTJyDf5
c5aVFO3Xy6m+4VPqrb2W8nk5bhaxME6GgECgEa4EWvuVoPAU6Ci/qYT4EmpHx6uwAeWVXI2e4T42
uDNJpC/m+naJuC+Zwym/+M5LK6GxiRX4yhDznrcv7AHOBYK0t1FUVPxL3yu+hM2SjfambqeSHFI7
aWND5c1qhOBbFaRYnhsKAmirnSZPwo7PGJWi3fiQpv7h9bfpkAkcv/UpUNEwtpBtj1jzh6dN7OPw
reBdXsT+fhWjuoeG022WoMIhEsmn00CPDYDzPJIoLc81Fc9+sFsX5yCe0EfY/OSBNQJUdkHeF4Jd
R52JLrvvkZhw+ru3h6WLbWeLWl3Pf1Ld7TjrshIs2H0jQJS4qikQ2sNE1Oz8DHY4ijMiSGLuUvgE
/Ve3cpQ20zuYvj9/QYTPD4y5rc/VojaBAuhKW0tXFfafH8o2QdlIO51FNWH9WNsUH18aUE/AEMf5
jW6mCwqAE4kRbBya6AUCH6c28n/EddhpF8GDaw/77lTDRbhB1alcLJfNDyu2tvHWFdGoJIZHH7cR
v7vGGFkFoy4NAEnIoEFYtqGRZ3rdn8xrlDR5/BWtOnCTT8do0S1DcM5y2DNINWrJKRZxq6mincxW
hhQFSJp0YTDuf9p0HoGkxGE/7WzUgnZrMFCEyI52sMHP8MxHVJtXSyiTTLyhOcOmn17T1yr6aKIC
8X6tvQGfdiPkLrLk9o1MpZ7o2mM6qWWHvHEG9BOs5G8xdk+lmw5NtaeAlyQ6JwQgU3b7oVd/DmQG
rK0HIsm6m/BnBsROsg6Cg90SFKWGsuPB9bkJxpKsUKvP4eh02hlG5XmykPzsQKcVheL906NlJp45
2A3jrzNbUItFnXdLJ04d1B/5jV6zcIHUFXK/8x1poqj/+pNiUS7Xu9OAVgIvvHrmd+94L66tKMGf
vCymw3XCD7nFIEvQmB4bknEE0EEC4PzGJmO0MUYrSofsXwXJ/qsHOCP/rfrPx+4X5FZ7yHnEutw1
PEjunW2P4+3lm2LAhWuupsV2xxoEonYTtKfGhcxDNLsAivPlf9WAtaPF+cay8w9gPQBcBa5XzAAi
xfQCbhvQ90Dk7oMXnBnya34Hj14fPpokuzg+raOHWK87pBDdJPC4iedi+9msEkpEt6lxsOENrDzM
fcjU+skpzTCxFUIF+be2Xh0YD+l6dTx6KQRurpcZ7Q/lK1OP0If0wHwXuGkb/D57J5LQNmNT7qKF
8/LVcwyv4mGaSAPpIyFK/lZ3TrpfgwDFsVJTUaFYsKpKGYlvBiLIG3mwGVyzzzCB9RYbT+sezOOM
nMcjlrpfzpXglx5M3Aq5hG7Ehnjm07Kiirb58Aj7P/5ZVU6agwk3uamlDTPJvCDBtT5TCy/1I6Nl
2Gugrv/QubK9gFbiTXkw2t5d+enhR6WlbSZbepgD6PbxD9gmzF1QWUBICg16zQgCv/EHNbAHpeZd
G2r9P1Z/+Myp78VrDdxSge7+jefGFurAvNGGtt5frvxR/V7pfkp/jnYE1Igh7Y5G+PeB2bAt9/fM
HB58Io5MuGI8Lf8qOyUBBLBKE5rCX7SI3rGmwW+MOXpDFZzpTWt7vkAmlFOQI0VkaVv9BnCLN/Kz
QaQBIsgXePhqJbfZM4iLO3ATcDp88UEKWfqXtflS+Hy53Kj5yhNkm7HkDSMB/SmbXVc0pnWM4tEb
+xaeYssKQpxowtnsQXrR8v+r9PoLIiZ1/LPR1vOR130XaCriQCJy0ojIlGLN3mGysuiCiHOJAy9I
zFv3pmzcEU5Kka+K07TU6w9yo8+NuytbjCf+J9SorQaROBsVojXlZP8IvD0h+a3pPgZLKomTKSz6
QRvvNAxqJLLqThAY42hxJt3+duzcxuNKLMOZ5pjEoUOe5gGZ9FbYuvXgVIdDnW5Y/OlGA75W7EWU
41Kl/aifuCID3oebHgIG66Nye/qv3pKH2/UvDqsetcwP3VVZ3STxdaZ12WudRlg2BuCzT9B16G83
XeMRrBTVKSTUttJ6tEP1UeiNfNAjoiORZygJ1RhDNvcZav7vf+d/vJgXb1tErWIWPr1ng6gkYgfj
nOFNeei3qctJ57CJaBlfbj8VdJibujXgG4shscqpXDnFphFKoyOh8wdTbJ3rdngN3CWChidMZGjO
NDLMKMd2BxQnP5MB1ZY9ST6ho6Igv+d0USGb/hSrKolwbKwwqnpgZWIXy+bQzl5Ra8L96oEcoPed
iJHY2fP5uWDFndjWS5Ncy62tPTUA176Q1xdGJitTc7B5STN55lSZv76vBnwnvuXL63j/2RnTjaQd
jevOf9sgQv+z/4ChP4StaPMAfcYBV4oRTO0B8ffTO11PMh5u6YQs8GwYvu0q6WmP0GrvgucrJdM9
svdWfuDpoQjetczX/eDPei3G9y3rTuog+bobTS5rVCkPif8LWoH09O0XFuO43/uK9kcyaN15q84c
vFp3c3y/YRjfHq0TTgarlYN5ZJWhspZS8eYGIZC1V3xSz747T2xgY2YlCmiDtTzzTgMQQqxnMdi9
FqDVKh480i66wOmhPlEMEfOpRxwssNOcRmYHCMy3Ejvq5lZdMVRN8y1dxSzpMUyF049BY7lyM7Tq
0nld+TJozppVHbKsBOhStfEzBli7zrA7SaTtEV5//f04vpkFqJvegyYI2eh/4sNI7IcPsu8rBEMZ
Kog9EvwOvzAofNGuB9uJIGTGplxU9L05kVg6BX8HPxFnB/TKuA2/JdG8C71Z3/apwNxIcuzD/EwX
nVOzKCt7ya1IuaJ2u1ZWD7S3Es+6VhYNQFxnb4572dbFfjBy4ippIWqFvCbouOR1Bt3IcyimNOLQ
4jgEncjtLQYtNQ4KseACRs4FvVmRqBgLnGCAraCF+PzwggUMrcvpxzv1ezcImQCPbP1HKQxC+0wj
+QbRu8cXxaXeFpulcXvszWLtAt+O//uylrL+Sf5sofFUdO2A7h0byZzEjaC4GP/Up0VI6nn949fA
y3I1/tcxib8fxP9+xELV2idyDfGYSkLLK16eOEv7LozenCf9H89RmPN0KiwH7guxESY6iOLhGcfT
K9SFRUYIpq2bO54iXKxaCoP4W2Gw8Mj/9gu/yYJoS1Bt9AKvM5W1OJFD9jK7Rw9nv3AgNRoBH8O9
r4xbdlCZY7YdGJqDnfpkSWtvjWc8cSudi2BsWpaRVOdP2cjfS1+MybnVe0B0Yv3HuApi5C/fOcUS
gqXCzYFU+8VvIgZYiY7UUPZxUoJ1+SGUzl9MDZIWrMCFGId3oLsSai/ozCLTawPuqsuHbe8oBdvy
WrVawA+dg7VDqjdl6SggDUOaPbHLIIuwDluYClUV5oNnRL7A5sMQRxkCynknXa3vpQWE208bJ96b
Qf9Pq4+IBAWkCjZsXV7NiWdQ+/Ca3Dxpq95CpJ6TlJ/WHKy32BoOdI+51sZee6MjQUEGK7oPmzN3
BTHCqnjDO8TSp6ZbT6o60HRT0dZexfqsROPIJiht1p6rX+zqPKOpN1lgHHrQZSGUUig4CZA0qpnH
5/wV19Po8a2ymTFniVvqEniksEXoWOVdOFWqySsHXsCOaEDEPmsT0fyXzmRBpPEW7hB5t96MSkMU
juO7zDjXyyGz4LYgRdcv50sjcIVsPYgYtLrBBlVeJcMlZHUSO7cm7V35vflqaF1A8tK36cVfnrHj
/EHTQSmgfeunOU9es+Lysz9WY+4cJoQcOhDjYkCDLM67+AI42N1J5d0Eto12jkzwmRMXX1SY8ir7
ncr04IQ0DcxJ0CyMZrtRvtyghsAtsdALxvcI5ooKh5DoHfg0Qb9XXGj2iTxIGp7STSCe+GLbtbSY
ijqLYhjTduQci6MqQJKlODxUwH6Du8raJwyZaaVAir0vlUFz9YnfbQf48+O1XMFsjAFZryKwfB0L
tdfjImY95LmZTefFhxbQ18rymJpca55Z6BpyGMPoDXdG7nhVT3r3k/QTPzeiuybV+G4qE+9kHUX3
CKES1x7TKpjJ8Wewyi+eb1uSnviUp/Pydd/bFOh+4foKCAt8kZbRWwROkMo5RnccJNygipwpXXjy
6Ua4l8eaJ7By3/Ij9TX8ikau8/Db39Q3mu3GV9jDsdajSCF9Hk2px8dt9p7tMnjgsubdann8zBtC
qe+mV+ayDfbUcPZMWJxHKHlOuFVMGmBaxibNhuKOOZXjMhZSQPl2t2t7VoXnXUhF0H6YDI9Vbbgu
gXuOQ4i/o/LhYE0LU5PGyhUoP2E16BT41U8vJGMnbIfi8ckeZHTXKjQ8IKP0HxEnsJ+S3WFj0Iom
MqK2sOdokdWhRwNaZrmA8BQ1BWa8dsuJ55JSDw3XCkkxe+1HafHxiq0e6CksBByjHaLo0WdbAAlK
iA4olQSv3NSEyX3Kt2ViqogV0Q+poCs0oC/hzvjxaIDU4yRXkCzVggvzo+sQUxt3Q7nUm8Lclq9M
k/NrO7IXLey5A4dxth+DyaFyWS67/9z6rxuHJGNebQUQ27ySGkXl/01jJjYilIIxFMjaYq0Shx5s
pt8ycRER182i3inovSrdaxIBNeeYwEgtxMf8t7hEuDINY3smqXJqzYCyda0enKFE1kRFh+HQY3E2
hMwSXbj2ZRdCTKcPJA+3PbiObCTEbJmiulMhPBuCKWp/4uAxCn4UYh6JOQbtMsJGTOzp1OJSA/mA
VTVSP5NuyX0ilM/TYy8tl+jvjAT2EJs2OJqmSS90Z1d6K9j91IsNPeq5rtEKxBMZX957wOARaCxe
loitw8LOU+qUYsnOhVbLuf3imL5fIqD8Ek72/mmQAOPnNuoPSbgzo6+USDOsqf03Yyw2wfLwIAIf
4TjQA3LU9XbbIcetgVCaAhcOvKNQK9mvlQczPs73USbVb/I3GT4rty1sJCRnmRv0A1tsV4Ec3iKJ
VJ7S1kRxL1f16U8JVZu1y8r+wEQJVx5GLVjBXg0UYq63LyxVLjRvcCS8DAEx7Otr5Nznuw/UER8w
vxVtGWT/zJyGpPxFkGLGj1xOtAFwi3TjUJvB0jSHgu4f6Mr07a/Shxf5700v6Kxcgb9Zq/MScuDM
9K75GhvHyfHqxcjJH+pr4dgyJqy0CDSbr0bZuqfGE6EkEUkEHeEddJ3AhrKDz0fdee4elis7CVE0
B/3qLkb8DOnrnTM8GWNBdH6cqm76/3ZA6izA3fAfWJfCYA2UJir6InznwOde1L1viGxxGgKCOsik
/AYGrdV1kf054qwjdXbIdgmlGxBwS1yse9hqYVoiQ75ahEkjdY+pgQrBc5zoLn4B4obAL4gHVj3K
2B68ktqbfM5hjGAiW2iQVOUbhRv+F0KErhptBA2qcKsEbALBwUPEs6K+e73KpPy9b9JGAK25Y35W
HbqwJnLeXJwfEbRyOVWkWX9CKUjbVTGj3EmcBSZXsjDNbEw25ZlFDBaH+x+Z+vb+gyVvGcmutOcV
xn53qKxnhpY6Vr5YDfueoB4W8/seHv/rig1knQhWdY2MRYptdVBwBhacussAO+Kp8Evgeh3tP2Qf
L3ZqbtWeqtnvJkWZEswfEjsqFIwJkvDeI78n1pInKtbKwKp5z7SGL4RVKw6bpfBveno8cvNzeHlE
nVglo9IO/IvdOBD5PSAlsPcH6KD/sKwFdU+Yy+LZe2JKuiYXLjq0nUgA0JDiKhlQy1j6EZSsRHKW
v/mNyFwQ0RDrzi6pNhKEYI4IhbsUADUGwIdEsDdHZHbKF52l/hmsjiQT0Eh7B+zQVb9Yjew+3dWs
vMGlp9r9RjpBCQYqCTS93pp69JFVUixAYgwbDD2x80ZTkvT8F5Zv98uIEpaK8oF2xaG1I2At1rEZ
WSE4kF+o24j+XCdhmQS9T5M9XssJJcmMjsQo+1UA6UYcDVYaY5akA8xs6Mk99k5DzUz81qLH44vV
W+v5CUrdFFoW5SCm6EEw/FZ0nsJJhgZ4jQynHSbRFgN67oTO++oWC2N0bZKKn5k3cmrCOQ0woNhd
pGZrTv5Obmw1cfLv2gbBn/+wwP5WtdrAeBoPjic/U1JgouLObNt3vR7SuwpuV6KL5CJ5173Z7Pua
c5RkirJb4lgAed7qeavLYiQPQiL4SJkNY9Cde1VRg6aFxy+3ZQQbVIhB1A31YFXOg5FIMSazb2CH
H6iNtpaTK0b5xnDd5MN9RhCznpYRqpiUSRLL4ZXjq6V6+m15YatqifyJ0Dio43s/n1L6h2Z00JGC
K/sxt624+QLkvDiF4XOHlY3pUZlj+IyK0M2MrjJsoF5o/nVT4CksR8HqExYKUYg6KmqhSrR30HtV
XYdGdMP3U7IK9roW61fcPhiX69jSRrlSxEFPNiElerZ27xQL9HPdJ0k7bSN+3QjAT5Z40OkSe1Na
vIrQRwnEcD2aC/FDgvTOWnb2U1u661Sv9GwFvQMmEYGZrXrINlr2T2r1EnxTFValCoE6caTh3Cp6
ISPcJpZYacZo73Aph1RQz/e3X8q3/aLuoM7uAxiwf4GINCrLftxZTKIfeCrEU8kMkEzJmc7Ya+Ar
KUnMaUYN1ZkJ8pAgipMPvuIpnoKHPkNuvBuXtJFgvnRgOPHL1rtrlcS+PRb91KAGIMFXfk0ghYF2
LLXO8Exrn7UwUEmHgUrsV71KzzAipIhodQCKAET1gRILQMG2d3/98DoyELcld/Fcm7FuN6jbirMc
K/RkxuX9ePrRvu31E/9EDSuG9hFn2XElnUNEm8UmuLT0ZQavsNgqpWO6rjzZD8yrP4TJpfzJ90he
YwvUYNMYcp2kJ4Zd6n5uSS3JdUzixxIpQdHCi5rikpKIpYNIztI2NuviHykbx9G7micmzQOUoLGq
tDPBRGr0N+3DrY1aY2Ld4wZO+Hz0e6VEe2B0A1qJWoRkFJn+K2hqV/dxSooth48sAOoangMnGslI
58oONxzgFflwHKDFgIIcevn9NO3/eZ57U4dxMMfSqGTp4BIlNjGQZNZqSHOEZqaXExKQmaV7/3lx
vZeyXgGXAIPFwgS/nksAKhdSIrJM0Gt1AtzcqwVfCSvgk0NjsMI+//uDtInBvJJS0hNeQglhkr8O
pDjHGbDwyKXHrUsTZEuXT14RzwJrWNdBTAFLH3OWirM3znbAUdDhGpN4vzNruALi4CG4q/jzsqzR
xUrHD3d8y1Kx8V3mL5hGqxaKsinLbi48b2AVwC4rLwssmp+BveKmSnl1CftFUYO3UZLnABdS1xCo
eAW0FohA9ll2tkZ/Dc7c5LTmdIW6Qm7XMSg1O+GkpgK6pEYaw0D2/FK8F+t3/TcU65bTGotPDmb3
wQQQ6Wpw6hBd3/UmCU28lKp+OFygZZFYfCn2nU4e5q3MqGfEya6dknb0pa2JV7DCMOPPa8XcLfwj
/j4JFwknoZEgrPQOzTDnPo8JMd4rvzSnxP7D1KdqVK2uMabk7wA3vcxwevlVFLH0RTpkVvrnbcyi
1CiboOXBMAScRys5aqwt44yvkH+qSmLYaOmu/6eV5s1ov7Of6VPNBJz6KHFjB5KTexVZQICaVtqa
QpPQNxa+GH4UZP9i7xBspEvYfjtNGeircaG6dfSNi8Jjwf/zlZGv1yPxF9M5l44F63nsvh3w1+1H
48EYk13FLsnsbTGPee8F1zARw2TBf4AkkNcTFXMICaXF/a8nAU8UOIhP8TYSXZ1VHiPCNVVKi3LG
kaA1bLdXfwvcw6Io8LED6RruRSWeEzRUW9oOdLh8mMeVCF+Tr1WYXf+IpHHLVV+F/+19wDjfWgF8
ufejXGris+U1lonyWLHqMK3oOB/xg3BmpBzcof4JBo89kPSmrPSfuF+sDfvu2AEYh4SH0fX0w0ar
LZtYZza7pSzys4HC8dxBMDWsntxWVgeVCgt75XNqRPFOl9EV/kfeZa3M/ZHowiaw4T9gxMn2X/E0
28m4fkNSNAi6TDiMaT381ev9/4nxEj2eklo+d8qWSUHEBkA1GT77o6jcGk5p0Xw2Z5xR994o7QqJ
SsIjlmOD3vpoDdD+fMCJH0UtK+qPfOcjeFPOxWz0Ry51fnaxiijpsuzwRisBllOdexVOLxxdQ0+a
E7uP3l80VA37l108I6jjfd6xZUw0FCVDcYwPwcIsf/DyqgA3XywD5m8XvMPguQDoIl5UI0seOXYs
gUQNQmwvRoN8/vW7mVg3fGBkrmD4FLp/h3amyS+Qm+qrlnc1ExXIg9yFYtcrIG1vbrNOQsOF4xTO
sb99eDiWX/OPC5CtgAPbXZWpd4WeNi9LcfN0TSEJZRBhpYaWSkvSSWRGEo4ZBqG2iuybCzCueXp6
0ZpChlMmRoYpxxwJ0Ign3wQPRjj72bV72jIgvxac0L30/6y9PwhHOpfvK2tYv9GM/tiVcZKR9ygJ
Yp+drjG9QSMViyek4om1KZMMCEe984HdyhV3tdEFy/CN9AHPROx1hM3riDskNopCbQUGrBDJXqmP
hCwgo880lnNz5vubBSEt1eascaS2FRz+9VQMyUE4z77eq417G8eGnWMfZabOkA2D41XcRJDscZn/
0Z+0XzK8FWcxFIvyhf+QlIqlO/c4pZsknEfuqXtvXO+76djhbL10qMbVYEFpd4WjRxD2ryITawg7
8bmoSZpCq3+hzkYI01euwWsYbvDZHg1FuPSPwMWYfdkn0M+2JlEcWz3j6uzBjagFSfYInv83Wq/m
LzcL+YiSGBo6CRfTvWmXonSZ9D7axxprxoUPzkysWgl0/vtGy1MYfnPacVxnrCSor6IyiNm/J7a6
+tKJ9yKLSbjLECGeapX8oWWMk8m59UTk+3oYJMHPPFPWqd2MNY/Ko9UZZcJqnluLmqMqZuvT0f2w
jRUdrErZd/0/2qHLqeq99KuBh6rZ2qf4sekwe4awSvixB4rNiW5FBQvZPAN+oHC0DvqIKjGVeV5+
+sG/noNUNNhbckQjQ6ckVY0SojbxkMaGVVCxRaJ+wssRz1SjH3BnGXH+5dAYskjFjhQjOrbbFrA4
HGTF4ugz12D2Wc5GBFv5yvNQ6DBxAJojzczaUlfT3DbOIRIEyWoPb/JzQgJ3g5MU+H5wN6rgdPPN
JXG6Zaa0NkGkm51YsQW0q130yjkbxI5HGewVju3B77uoUAVRquOe7rjdZuAOSF4CqJ9Isa6s7CvB
XNrJFVyHCG9NgJzu0ap6N6IrMV3J88IkYgYCyaX7Xkm+UNqOqpV8HTAATv+sbOtAc8Kj8KPGCNRE
v3IMh2Gn6bae2Zirab9EbJu9vkP5IhrzFEMQH4EjkiJ0vBVUyUsIZGd/2nr9yI1nyfb/8lBcZLCR
IHGVQZhuqEQ2jsbAY/dkVqktyqna6hAaIxNSePHAEI2YGI9u+k1n0DZ8xsfU2K8DfhN59rz6nmYG
O0iHJCSD0Lp+NukBrZ8zxDtjJGWBk2OL46h31XjJsr1MPweCA/lPCMVSAs47bp2abuzdOvZ69syX
7Nhoxo46Fqf/kO0C/9MITlJCCzHr04C+srZgV8NQGuhWPsinQ/Nfv/EQG8OKGGCmQ2cQAR7Z35eJ
u863VdKh9dV55PYDSGNpAq5XpddbfgzjlC9PrkdNvRZB+DjNpchQH+BUEmDIJqI6nCb+3Ndt4cUS
xXyoPgmPc7oAoDSm6BtXn6WcBUNuk7RUNTgFqJnNJY6Fe0N0cTw5EqmK+VBKpXCbaoV+fPoe+Pg2
7noNEKidsmLj4hPH2lHN2nxb9Qfm4BAN55xVmkSXvJpL8APrMvVu+H1+OMKczPg/uMaX+GcKKTeI
jHXA9IifmwErniZz3ovVLe4TwVJZr+A+sm7MfO8Zn+YK4X+5aVhrGzO3bj9E5ks4/VYVpvGW4YOL
KGAitYiLuKtEwF1fsGLG8L86bQCCe7zUAylQzoPAZRDmqT0ly7CEUfSMN4yybgPzWdamkuMlhFdr
UZPMQGja1OE8zG+s58YFiZ6iJgePj+u+LoBNx1gt966ELk2dgci06Z3u94xMDVHTLMe0dTp1uVgi
wBjZHKqK0adU0TKWMP7IJccNrHiaROifjjLi3ZBNcxK8BlAxOQNVakQIsKOS/n4PB4NAfbw8D8F5
e1UuHIeZVpA25o0jYv64bfq5pGaQhNjKYViURaFBNDxSaMV4ctr4ZYCgACT8I6rei+Ya6GPLTAqQ
ZWTD1J8mrjQDD7J5aDs66V1r34q6S3tCp9Pk38x7HEP/ex9ZcftOzCrCHZJUWUf6W+jskMCMn04s
TwDPNsKMyobF8kaO1UYSxFnUIBEFMFNgEFpebv0oEevLHSteyhdBRIBMhIjO1stbCv8dmogb0n8j
V38Qt9UsquQL1PoJJynq0/1/6f1L/vvP7cNGj23LMc9Ny97Xrdmz9Qn9Ld/vB+lTIc0UiWDNSapH
BWV/BoqV6EC64ce4aVJjfB9fOIMcFYaONNlSSeEps2nP3uu/7HEiKZe58R1d/zGqoEAYM7yIagSu
1eD/a6h+EPiegreHKv4p0YWlR3R63tP4XgHn/Jof7AvIqJ+qQiVBm/oejZsKVVBdCzpZwUZGoisZ
3NAaPSK2VKEdTHDqaeZ0a2VUesOR1Vn7CaTTGjWO4FnpDh/qUcWKAl2ui+U+zdO+zBCjFkvhIWSI
AOtxtUsNIIiUPeEcKLL9kC09Brev3wasLtzdrbhGPOWK+70JgDvCyjAtSXQ3+Qzqwp9/GmvLESog
v2FZKZwy/ZcruLwWpXKS3xfak0ixMtocN1TgCFB6W9llEyLRuvJnXCLUgskdFtvtFmimGAyWtvo6
gGuGxEQ4dFYUDC8t66LJLSy/UOPEujlddTCIr+DmQoDUDkAgwpeELvzxca34y09Qz37fzmoBwDqG
mUmL+5/4fRY0EG9Ekm2ZEDGTowqjJ9d/qGkWsooQKLjAXgckS7ufEDMc8LQ+hLXgMx6mh2Lqo21j
vO6wq/Y0OA5anoUnzNl2zKAbEZrckDF08sBEOacRDbbCzX6mwSwfOJ2jF6QE+9Rxqnxhnl+OLC6X
uvTUvILB7XS1nv0adwEX0hNOuyMv/y5JKPKTCpvJVMmfGTOvuc3ShkrpcRextJMBOE1oV3aFG6aG
HEra0cKbUHEXH2MaaJUlGDZWlmMlXn7+I8m4XJCmgG4rkc6vRWWNOvKxstNb0qiwLOYTqy38XpCp
lAiIKxdZMvfkkLwynuLg4PQC++dBqDaAHk8Q6JmhC1FfgVOCqx0klDO/u0T+g8rgI/E87kpv94KU
oH/eJVUho7isD/iNFYD/vwQ5KMgn140Pz1iV2NGqPtlaiFS5gy1KoWOFkppqUm//RVXihi3mCdMd
KKllrBnz7+JhrMde4+ywL2rEC54srAOfTMf3wfu7nVJmJhRmNPiY4o2QSuQpmhBI+rVbZ6SUYYrz
wEaAhhltt07q//dMG4X3yjZUP71IBTyT9YlySWxXWM5YNZJhuz7UWy6SxDC1j57zCYlYoNH4D03G
vhf+mOJhgtgqgi6vXB+B3eruD9/zg5kaojcetkD59wtewLCpm3ah6Z4qFQieKe/4yQXbPtSHB32B
JAERaYVJA5A2YFwsTn1UASR1rcZs5TMIBzLKDbmE+7BzVo59CWNf27wZXunHGEQNHme5/f2sMbsh
x6C5YAnFCVkmKeQQW1S99ozWtU8OClAAwTGIZqmAXL4f51Tsap++WaiIYnL8Aj+00MbfsZRT+Ilc
SVYIL7b71YOJTovA4Yx9/5LlXhiDkaIt31qcKXeBxZUCP5xW8pjGDrbU9tGaRLlocbf/d7/CmAoY
9GsVlHLCDgmVKhChJi+8065HiiRvQzPR7sHIieXnaOtya8jNQNzDefQNf328mYfjphIcQfGwQZKV
jI7pMIDjzU/lZ9cLKOlAi9U9A/eXggGDaDLUMNS43sMbHsefVCJcMC2gV6X4x4U2C+G+KJsUOtGX
92bL8Rfqv3AhH9aB3cdRWXY/IG46NxiGHiH5ir5J1/EJBb0xHm5DTZWyS95/m/92GI6eq7P2eBwK
N05IalwmjNd1moscCuospg2roHjiqlLL2Jj7NqwgeR90XI2I2NCOLyB2CYG4/RTBxlTyT8jENqKd
bzx8oMBkbmgeXWEA6YsOR5+pjE2fCxjj4fsBQ4ot1eItwrRWsEXVHr2pf4t8tK1Mz3owwa4zDelP
rlCpeXa6jQW4mXBaPig0D8rlIbdxZUFLxVlbM47zQShel5f7XkWGAH6urKQYALW+9CxxkGfZT6s1
Mb6YFLQcpM80DWvOon3a7CAY/WY3osprKkHqHs+itCaQZ773W7cqlw99QdmHupwQ0CwbKdp6YVY1
6iwGUt53sUnVNPeRQpqS5CD6KDuuXPZ8J9+hBC+xA5cQpgJ2PC+yl/POylv9wxd42ub6lESRfPpQ
uGEAovN/ijBCWDrX4Z5W6zv6Ub2dsh5TeQT/SyZsDs/CzjVVEyv1fvvgY6iUv199/hwSPpbIZ6G8
CXDXUIGVONtJpt+dYY85jIS4h8nOQ7cmRdQ/AuD1Aju2F9Z3O/pKq7RzcMJm9dI1KSkIIW+5773g
vp/jZLFbOF06cDhMrEMJd0dgTPyN6/wc25U2j0Nj8m1q13bqgr8AvBHfOmw6Yti4JQI/ZPLONX1w
ewEQu4UY3ccCIHdh0+KxQRoAP+01pe2MWfDytXfspaYvctG6cAYHihz22ijH+xKHKqcwtPixste/
Wt/elfN59OLWRZ4+vJxWyw8GGYiB6irlW38L6zxcXXg/Hzlf94jASNuxvZv1sOc5zk1FLsGnxCFR
qriiWjc7bD9zB9vcbT9f4N2U6EVuCKKBet1V/i1MF60o+CngiMOPZEwboewt1LERHY1tvsmJM1WH
Pntk0Sh/+eP8zFM7SkfLhZpv8joe6lAf2G0HgrLb/35Sl8JOlifzdJvbH87dmjEZyHX/dz97QZJa
vhgK632qI6aQ2I7ftFi6Nm+AWX4X7wyrEubN2FV8+KNdg3oRShjH3zvCl4x6HkYFGmZ0OIzS8GjC
vTiZerdUcXB5npXZUTnWxh29JwsbS1l3wleepxYMHXTxgcgTePYjvm5w+eUWgQJHpZvMWXGZoe82
gib7+VxCMG2lStUf8n78p6q39LERibtYAyeo/BNnWsuRr+4uxf7ixQCZBBsWtE8D7YJwjP/IamhE
l7XFSHx20wcYGfgJFk32iteQE9it48LgyNgSu7saMW5Gl39aZJiAdQ9xXb01bwUaNueqUVPHsfk+
/mWbW4EL7cXig+vDRps7K7racNEV78jTn6Ab3qWEH9kBK1KtHSIF1ShdxKVl4IbXET5gHMHjpx7R
BZdMNlzgNJpJf49ET2Ay9ScIzJE9KLwU/HYKH0nqznaoNmjgdb8ZCDGctsiIS698Dy6/CdfnxhTh
S71LmzjE2R7bbn6AcbWuARNYEpqnU81p09S+tkmzV8zVF7F1jC/f224qG+1gElGHurpIoOy7HwGR
f8oZhEW7z1Jw2wU0MMN8/dyyqkd3Vfqth2Rp9+EasQJRnbF5gS7F2Mi1j/p7l2brHcDJcqhtHeTf
dh0AdnVqCnviTKnw1dHuzhKXOfF5SxV4hdp5E/HJg85JhSFcEQYIB+3pU9oCeIPFKexXGBI1vlti
TetqYTCLkntTgTA8rzGHE8fwkhYTwjruz4FYfx/Q6NsTYJJb8sd8u0YCwTyn0p1CKQmMQuTdL8hK
zD1qhkeiylIxGWMRrIyEhF/AN1V7vozKt7bjKjn49AmLSgYKEsC33MNQ8fELXp/e0VkGc9qjXMa+
0TrPYoGqXSroxDuiREy22ZI44Hy2OVwuzLgNSn9HpzdLOm4X/QW9QwwXVmX2npWtq+ZXveL2PFT7
xTgavNqlE8cQ/2gaimz7GL2yhLkibIooMV7YrSIwdDLaXZOs/+JmPEwabg1AqERv/uGOa6fgvVMu
sBqg/QEoMDqCl8pUrYQ7luLqldK0/85MPTPNSdVI1R6lt4H8PsquKq6eXVFvWFiL3fQNyH124VHn
JLRPdJWtwlsQzGMi/up074xAiUYExSPoA/W80oh39XQ6JF1up4C3IU7odjCNE7n9Y6MsdT17GGbC
Dl4QYAKEjXyab9HMhyeTNipi40jpPzn910INDEiwA7+jbV4WdfAcKBJsArTHFNLCM1lXfWZ0/oJS
a6LP6pRDH+yqW8tZYkPBzwwb18Urdv1qZols8YHrANeTz4mgUbCODSL54Or02AnehjVZazaktXTq
Bz70lY6siULh+rst/gRHTEVxthKymF5o87LvV+XPKcR7XFHkf7FaIF26RceewkfwG47MH8KUyCzO
NIGZ6kh2ZZlrEHyuV8XlrJpUoRd3KAxMbHtJBh+iBYFmEbenWkk0wbvCIjtkgL1rX9Ce5akvVLzg
ofMxmL/RiXFhZC6A+C76IkUDlcu6ZtLFCfnDpX3ndGDnxXFxVsT2n/pBajzNUjTQecJq06rE/Icc
wCOC25xzSVflz1xpa6xe5/NqWjxhM/fxewdC84/T5kfzoX/HmuIDIi2T/KYUGo+nZT46szxveqYF
RR/o0RkvXdF+kRXIuJq/0iaLMsQOpcZ5//E3PWZAFAIsMjR6GnuJ2rhf22WN/W7t23ROLsE3bJ1N
YOPs//k32AxSIiixwPSdPzFy3F1qjqRaAS1EufItRNF2LZQuIJnIfKcVwFhsGikYd0jgd+FLPkOb
kfLfjXy5FLBo57j16b8hlkP6Wpq+mmCp+yEFKkrt/l8i6pig/id5FSGhiEWpRx9+ApqlFWTavDQC
SA2FiJbSJfBMRHQw92uu/lHV3/8XjtWsjRzFhBLaKLkHZ+HqtUGyZTE6Api80672Q1cjSM8nh7m9
rOL4T2mDXj1UkiCREYsRlXpmwk+tcwFIyn6DAHGAc3thTmCixTQdDR0JhHkIYBfdqdHhg5g0HkLt
ZpX0ny0oZOI7P/AqqkXSKZtLRirSAh23Lihu1dMGbBVueDd5XTX2zTYKDns6vV76DLFT12S721re
aUcN/u1lPNQZWR2KCabI97wLO/uX7aOFV5B238wxSEW6z7DXb1W1MED17HPSbZoeCAtWuwziRKnl
/7waUHYXLXzZG23At0d+fLZbfTv27xm6/3VG93hxNvq3XE6CZ/bDSvwbK30jIAYnFPkTmBLk3/dB
jKQvxpqRdoui/JM5VPviHhcR9hUf1Hp62KQGY6hGl4uOYOqdA2EmUVKl8zff95ep0OTm6luqplW+
O4sGkfeUmI9Qt4EJSgBQSZa2jPnyqyonIIqRhUAQh3WbtYfCeOtTNmXt3nXZLpJSXUtA50LBzPXo
TtUEzJe+RGcKB6eq/u6jnWS4K9soy1t7lEHvA0XXcBZv6rb+gS6SSj0InixgpSRLIZDWtBInF4Ah
wGQeuiQsuvi5uWbCrZC3lsFbhINLJaIIFgtnegE1iPnMp5xfbHINpvdu+T/SzTKSkYIdz95IwYDu
0X7dDlppYq0RZ+FOnxTGiRlzyVxSqAxEdJyyZaUMTEK8vhgOzcD/ppqZLEuJXAPNXHG7/aoeTPYP
0r/WJ7Fr5YWni04fErWZFNoAiOe8dXjzdMkvNJpCdSX68Wu8oUv6JJRRQdEHimGI8H8z4aa1VWyF
YRcDvLQrYUzcZmOfZgPGP14YHyM1TdXTXpXEKcz5Fqm7odEdLUhd8x7aFlFdWRNdYKKHcwmDPovg
rbOiWwUZ77A5N+/ikWYvwmT7tc5i9mhkhygMlwQ6VbhvtKJJwSuNZjDtleXFC1hVFrg/tKRSP+yZ
xhqBqJm0tA3kHKym9SsMIXTnbqR6ExAqvWHfARzmhaspv2ZhDqcklZsNKnL5XI/uQH5Ks1gSSMbe
Jm5heLigfNFDguTskli+6wcekzcqHpltVSFr7Hu0nagRlfkTbXomSwKJGRUh+EtbQyHT1LxQ3O14
Czn7qRqaihrNr9STo85o22Zlt502k3C0TIWWpLgZAFg3iQ97LwyDcJE/vTq76AIVKkpSqwYERHk3
210MziselbnLS2LtX9koY1TEa3yY2BpI6JRxMniW96mMtqwX/anlP78vllOmaD+6RzBVyEDTsr2b
4eLKzXuS6znl5AVkXZqnUivMpXHW0Z9rm0g6M9zW1V5bAajvXbEorpzJNZD4kfSl26ypItQqCTu1
oUa0XBWFHt6FGUJuOc60Wcwu5Ca2a+v/x5oLmf9Xm7WwHziUXqVspeY8NOD2QNsbXqcnzNpa9MNL
N0A6DoYCDifRfo4jmBmAtacZw/gGmk3g/x3zeIJ+xe6pJtz1zsfmqkzyStgtTrbHhARxlJoEKTjl
Y6dU33IyojG34OJn4BmZVGz18Akl8Xedgbhp0Xu3AvS6wS1EOkG1z9WiMdXFi6xpen7t7cMGjpgf
sVnQMVAzllKtbk27JOGWayV0jy2vZhVktl+qppRPzj/FtAGmuru9ZYx28hJLC2x9q+wOIRBpQrat
RiXYnbdv2UFR5ikEAy7R1SUxQl5Bjn+qfbPduYATPjNVHpjsjBfMW/0ESpKuQByTsYGWpELYHQDx
wAYpPX2ph/VBc+km3dMuvN40/W1BkYaN/rilZUxL7WC7dNbHxOxlNj1WdQl0PhYf8yYpgLdo9RiJ
niyugigfey0h3yDRSF8IGLvKJH3wuolYxZW4bNBrwtmDX2yYCyaS+hvcAd5vtwI6OjeyVs21hQ3I
/GB4PJ6SR5OhNpAZTO844o9iGEYxldgRAKChgkU9FW6s0D2vxpeNgQ1rcK6PBIQh2ox/MfnzA47W
wAz8id1zhX8JxPUiy/yU+sU5Jisl5+r/W8qTtTXIWvEB2PtCtBxLhtPAzND0rSFE+vsCb6v88rsB
hch/H08diKvbuAd6MDMzmwrT1tDw5Ck0Pe/SYfxvnIZNqcNM/aFm9PbVf1FZE+7sf+gQQw51XRh4
M8iNyz+9hPDZtQHNh6M5IwmhZSmZSsxyrKTmg5iVgMsuAIN/ZZ52xctCVu3UWJrpfVIhFalx+SAB
clM6m1KSuZJhOiwph0ljHfeqKauRbPk/ZT5+X0L9GnNyYvF3DPkpnnRe58ywLogk33i8Jl6zB246
LRdi7heBm/K55VGd0aU6YuYjxo+vDqVqerzTAyTa74P7FO4fSbLgKwTnrwMz0krtVssdu6LN7IR1
SzMMA+7m7/XIpjqQ3aaUSzZeFYb37oG8r1yKce+RjPzwGH+y4rS0t0L+fuRVW6DJBIo9WcQ9NE8G
8vUxSjFDroSJxvis6xY25SR5dFm9EjtBeHVQD2JBWtGwr/WgYlcRcqKAJ+4kATJzgqqA3mpLEkLr
SLc9DdyQ9PthwBMIysy0h5djYTRfofKL0D8abbzUHting6SpcgFIx55ILiFftMXqVdSM+ze02VWj
QeeSHtdMoNayiy7yK++dFwHL/pswlJ6uFwXJ4VvhMEYXkAtfT/oyhaS6Ce9/rfKvmH9T+iVeP+xs
jtEcQp3tCVBzF79OIcWoQL6UWp0cV1RfDJlghfLeyWLx90x7Y9CbWPbUJQOyv/kvY3NdpoPQOZfo
xtnceV1aBSyW+YFDrBfS2Fx3dmiPKmQFOO/l6reptgXaMB26FnpulCc7UdHhcab5KVeI7QuPQfDB
TTVOu7926gkYlPNNOw9xux118FQEPgSdK+L/iHVSxVGKcgj1kctK+Wilfuei2KtYP5ELdXQSQ0WS
l4HyV9d/D3aWdG1iZWSNP17uOXyJAc5Pq4RYDvpwpGrs1+k750upGwqGuz0LJ7M1wAqNIF+XsumM
aDO31cHjAQILEPrydrC2UHnebxRZpnYyZvAcvAJDo20AjUim0aBDSx1bvvViOLMOKNY3Qll/V44k
peRWnDvdgznUQyYrVughJJoYg5bXVYhNaPDbqWdpsvz56h7BVTuzF8qSIuvtngpT01QoxhkAsvyf
CNpPsD3fSWbhFWthCQKzfAgfwv3hGunK2WoSngM4c9wkOWivCtYhF2IlfoEyvKO88n88VmDjgES4
2JcHM242dNu2J+ldm+CYO3rbrRKaXU50h6wkJ5qH91li+aWBYFgjkiQuae6kaF/NoJJ4hTzlVd+c
GP5J6JAbSyK7mrZN5QUTH1HR+GN3Us1aVAW4QBohsTuxR9qILAqYB7vlz5RYT/297IVMYitodLAM
QRS10nPje49NhxLHfDLDghr0ltN+4QiidMwYNdezOZmyUftG92ytqsQIfrA21KqOGfw2wbFw9EWU
BRGSWLGVWwth7giEoPi4+/oRmkgwdKwgos3bMaD4WccmYixcTUrI6+ks0j5zv0eNi8edwYhkGK6S
LIDxvgHEnaNGhXfsYg2i+DwGIyrBK4jyst5L4Y+y8GYw4aElFcZQ4uNtVN5r71YIgpVlzbdUdk2x
XidBi0xsZCFnNIA4/+l/63OnUmKlU5f4lBngZUXg0JcQ6YOXL19G7QOKoVylYY+c8tjFauFBWHq4
j+JWOPW2vGff6/Qa6dZuzzKXIyhlE8zZNFd3hLLRMn//D+hrP+CScndeVW81Wxr4099RaOIXvfcz
PNRiBchS0ZxFO4SUJhigq8nzEyOF7Zksp7XUjThVO5MEMG7QxDotduj8pDAgfIibjiueyX9GNsaY
PwSXzHo7co8dCQNqlFDaQH76G2YFmcM/1t66ATt7oTUbDLMyNV657ySW9c6NEjYBrhFyhFxN2Pud
qICz5olAZGYrSsaYs2M6IQp32nRBqsCR6L2pwhK6OEltinUw8BshBic70SkOrAa4aNG3xmK0l7Hr
cYtagGxE+FrXIrmvth2O/nZxK/kDJry3VUtGQ/UsdYE/15OZHmx1DwD7EXgV35bpC6R6w0kKeh1N
Sbh8SlNBl5TlnjOs8rAVdH3KzkfPmaoMOhbvwACshx2+MItjxFuUt3Of0TNg+znEhfqWNF2VALR/
2UU8d4MMAQ0RKNRS9TyIQAJRilbI9RbQO/mrWgMe5Tjq+Z4YY/1WB6+puWSioDuIk2S8vTKX4UaL
0YRfDrR1XLDZbX36KxUn0rZ+SzlHv2P2337Sx6fnfOb2PIix7yi2vEkBSWlHfUVxiua4D/QbWfqL
1zL7QcPkckYoW4C8/GoOg2SL50sjcBvN6tC1arD4Nm1BdB58w4Y9+J2bU1WYE0MOU4BP6uD3W37O
kLvIREYsRQNanuVIa35ZjdnG3j8Ou+chWKvAO4i/p1wwNILx0YAYPNoETjiwJ53vecHj8VmbTfXm
zagYXboW1vD51PT9RULhIL16syqXk94HuTFzrnUv3K8CyDO7BxeJwq+N7qhDyWd837x9uquEAATj
QOJlc0k3QTGTE9uN5DMP31zMcMIEtqav2IZQShASw2y94ZhNAa0wnLTAZf1kcVeFJ0KNGVOUrroA
SEKJ9dRwf0sKe7JE7pAd3RPGOoswAcl5oYldXN/5zvTaYQzwaeq4UtpTgaiL9leli7yuXTzgwvfn
t80JxRrzqKC8kML4xLn6S3s3CR7nRzfMVmmxStThp9pcXnqfX56dzq6K/T02Lw/eL325od/mhAKj
fSCGDbBplyoTa9lhCggdNYiG28HN7zgWg/0j5eNXTNanifElWwYjNP0CcJcpGZnZ1V2OTvs1RrhP
xQ/2FJPqvhwJs9TF1cMenE8UscF6NM83SwHXS5NQKkmcDc+tw7azlFqaT0Y8AWhUdpQvbZ0mqU8R
XYxG3A2IOTl5CskzAN9f4QhGOgHbl2LhxmKg/HP9eCeRJe/+ysHYFpxjpYUUMxg0W2CyUgCS3J7Z
2QWTwZMuNHlVjzsf7SWKwuVCQ9FNSqkK1Bb4i2NOLO7Cae7w0+Ccp3lp8AoXNjOSMRbm7/jeWCpu
kQX58HgtY3Rb8mpv13Zi1dwKEG9O6iBzIwJ6Klf6VBNU+1AnXNDieQuXwuTRLYij4EhZk643nXvp
NsVLHJmnetzof1HDRvnkqMt26bZtkVjFumr9ED6qCIqFbPC0wtOVKWVHX00s7OtXYp7QXvzv5CuO
aqmpw5Dft3obXlzz0tMpAhrVAUO9jtAEB5Kdv6juwGmXMWtiQwW8gzEGPo6XZxbTp1Ck8z2MMNMn
4IscCXxfCJB1ZMIoowuvSrK67ONecrf6FR138lNPg7iIFfiqnYe10dkDgoJZJmBa+3Moga6VGYpV
6zxYfd5GHr4LOc2Bn/shyKEWRm+HBghLO0Eujah+gUEG5Pg+ks9hhz3S3YMV0mbuVGogd1Ys4Yzu
Z4D2T4KCWEf9v9DaAl5Hp6WSYIPWBaW5YCidSr+UywOxxakqgIMCMdKHCHlXS3OmpZ1FoDvK5tEr
b2D8inMzMUkZTUEJuTkCHChLuDDB5wC2OZk2tKwwavxdiv/6o83d/QZqg2Z44YnX0EJNvxvvfTgs
aJqWINu9kBl3bCZH7+YthckMJW9gwtmdzLaZ4BSk7gzwGXG1FM4rucqKaYplFI/QKsiDOk+25kJn
fjXnHEzHc1IlgbrktfeggqFjL8bqJrgi1MVSCNHpw94HEJmY1FSYZBULnke3qEvsqQ6bSI6XoCmy
9fQPrdhXCe+nUtL66Tu5ZSWLd8f7WsXNY6G3xiktDufwg3Cf6RBiD40Bq6oo9MspAWPv5AbZanPq
snoWS8uWUX3fPbfOFwSd/8XF/K7jhQsCvPOF8EDF6Ld0QELS1/TddhHzFGh1/Z0LoKt4xXoBtk41
tABHtzbbElQVn0a7NvV6X7B9BRE3O94hOGXWLevOeP46YUupO0hQBAuoibcHIQz/iuPhJRgNLD6d
1IDhOGKlemxqRcvatt1FXmcAm0gNXn2yb7odhqQs0t5jPoKbJRtVoND7U5Kd0nzUs+knQGOD7/iS
2jAvDRN/VUMq4UI0buOXxCu4OdesKJqqTCoc7WQXyXgrik831oe7IE33TVwt7pL1ZpWvxbwYFXlY
kXftSAnUcWZ3yfVff7BkG+0yzdQ2gMiMSC1OTCV0XHh4ZopOrNr7Z4s7MLKXz7YvfXAme2NjoL1a
NDbXbjR6LVVERtTw4hNxx+jgOKoxEYbh4RYaflFRV8iQ/sjD6ZMBoadsIXMOly2ctC7oViJ4IqZ+
NdcKjdrtMgidhkbVwUxXXC3yWvYRfeOlLfA3btn6kK4SK/lFnoImm9j2KTbuJXnCmRf3UtkXHR3p
TJzQhg1bTVoi3tbQzOPXubL/4s3jEe4n1WJ1pgxgv0BKlRKRNo+2oUKtnzSf4HFJK++gfhKO0B6P
r6IH1lf7VXcabWzhBCsH3+bB31KOsPcj1b2YO5cB74yUV8NoHTYtwBlwwJPP/VfCbL6X1Jq/xRK+
VJCI8TDBPHpEfoO4Y2xEtDtKzqOj5tYURFzXQJirEqxaz/xR6CHp0HAUsObzkj3GkuKZ+O1XLXU/
Q2Oe5rHONjRw49nGWyR2DvItPW2FDb3FpIvj/ZYEFe2/M2NA1qnelXxiePnPlx6uZH3z2gqn1H/1
SRl757kkKuUATuh3jkD1suKAYg4vrbregEahchFqUmAfi9pelin07EHQ8+7rnPQ4oQdt16P3kJjV
Q20b2XHeM+vXRIwaXZz400XcsfmyqfJtFtVh/K26545LlIs2c3OxEfW9wHkA63fj9P7jms+SGZ0v
fR8U6YTUsb7/Qtzs3v/IO/yavf4qau7qsGGAB2osg6KRsjZbYZ7cE2KrAoZujGbhDSXCZfW4Sebs
8zN4k/XZkNFO9e4Qy8nCdmLEzNe7ZxdECsn2q2dDp/wY+yqElrMwi3v83b5XtYRZIrwRlBQO0rT+
r30nrP66DLuuF6n2m/vJmIjd/06YLEK+Iio8/QnBEXWxayuctovjPBlEhc5K7Sk2FqpRHCXZ9X/A
uY/+44SQr+8q5SGkt3mc89fUSqGsSZ11LPLc7CLCmPARYhUzcYddxpwkaHHRClZrs3gQZZkfrmsb
nDl2xw1MB8CIisJRyGxXFdLe+ohMV5/A2YwhteQACFZemwT+32lhPgsDZ5xzPBT2is8xq3STaIc3
NbcC8x42CwVZyKlsPuGeAzK14VjyevAPBVHo0TYCmHutmaKVNpKV+Oj+pKqEcWNmwn7Erp+hmBWA
2G3puldFEARJwnarh+QtOTufqLIOKfbWmZS9EeDUMLuKeiTHAwCHLY4JYMGMNUqKFMvI10fGT9nw
EdnKaSRSxRaftG08ECeRLzPuTL497ObNku70nhhSlNZ3PtalUqqBxYp3yr29kd55tFQ3kF7iO1Xe
0yAtPyljhA/tLQsp6JLqKCdZSOvU30D3FkD3pGYhXPhQNcYg3ysrtu0b/cFm92y23U5Loddf3r9D
Zl7Hn7Bk4rtUuk5kPWfej9asNUf+Vltia5gadG8tkPaJV9RbFE0zT+vhlelNMmEzy+UoEWMSI01a
VffOd5v7lhz6sShzPFEpOjBrcGZpdoVTxxR0D0Rd5AONhgjWb+7PUQZFsJz4j3TZBRIprr/RBbon
I9Vx/m5BlRzPMpWpL3D+EbxYT9lL22Ze0NrOX+IjGTRXYPAnZfFmLGewZPC6awEFwm1xQaDXL2yu
iTGEhZzXxErB5yuyGyHAV/HtGcGf/f3FP1gYYhGxozhLsDIkSQWIBOBqWXEj2eogrylvfAB00gXU
UKuJCVWjS5pFBNASC4F0cUcemtBzP4KBkJP3SIuJv2X+mrr1f5mvw3QsKq7t4xE2wxTW1+4mdKB+
Iqf5Um9kLjtDGKDbJLtl5xYM6L2tW+MjWC0Iqnn9djSbac2L0QcuS/8WLm9GbOXufB2hfPjs/QM6
i8NDnAQxgRrf089k/8EWqKH+snpDGquUre2neXVsM7Koq+mgvnfsPqG/hhGUQoVVWfQHa4I2ulus
SbRDFFFgHssX1ZFd+rM+Zv7ggwftSkfmXVFnVGDPn5gNUWcbAcLhGLiw7ZUtRGLtw65kxGL6Pf1S
Mj+sM4qZnfH7hXClbo08hqRWjvskTkI9AhKql7IQDT/JDdEl9HjFYTsFBi+VNYJUZqyzwzBg3odh
1X5GVm+b5PW+MW0GBo51MmUnt2iNDVtca0MLhYuEABxuBdsQcoBdNG10K091umdHN9QME49zIbAt
Nf8ZqTWR4dzK4+pDWTX0kMh428kwGnKLIS9/6YOR12qURiE065acA0zJRo9OqiaYUYdrhMWDWm1h
M2YYDZUHx/GMSBn6O5SljwNE/sCn/jcCWvAnVtkZz/abrmzJx2kSUzDikAHVvkGPW3cDemYt5pES
YB/3V4splymnWGL3T3VuBsIpTI/jksFbggoJ/0Ctz1uqAgAq8H5WDqC3C/vf/it/yGPTbdTMpb4V
lX3n/Bn6MkhnCS6e8YCb+YXkf5cFKdeOWH6E/wMPgV6NBcqS34El+0ctV72UcCDNBhzXPKAz12TW
Q9MgOyeDnHhDNDOOXzPzP3t1YZANu2rg/aoA9MvWO3apEVQiqjCKbmmPU/UkKFfBFOIbZRUClDFG
x+XL6P6kk9VgYfmwDAuijTmbXHIkWSHF0hxKxKjs+KgK3TVoFOV1flQvtjU0GA/j9pmeuvHBDWy3
O83YAscZ0DUb3oiVaUZqxeoYuho2yAA/v/CQagan4xcCq0e7ncrfPBd9O5Afdkc5ff4XcQOYaCwo
iP6FXhrfW7eF8Q+9JumWvhrLnUQtEo4PWNJITs+pgx5ic7AkgiWIgWhEz1i82tYAvzYuQfKNtpRF
HK99jrIrth9dTB6Kq5bDtfj9MB5pqgtd594Lg4pfZxPrSH9dzTPNHurfvG4JUsy2hvMZgAB/EhLm
7zAEAie+u7VSU8cQFPhPSZQ9kFShFeufBAvUsMsSXJqmoYcsSCIzuqeexb7i4WQf66a+viVdfC1V
34ef6qhSj7A5R2A1XjvrDj40F/iMPc4vok7O3mMf+EP8MuWRCGaBKCdKFg0kWLwWx8WW2fmrdXh4
n5vgvaIDKy5JcVtriCf4J2nG9SDQ3kjOFWz1HEYhBhsfVHopCSmsL2fRQV4PNJQROS9vyRVCChtu
hpDBfV8m6yuFjUbxIHX4JSiiUCtC4c2QnccrdFg8OGTh9L8rDjcSDucwuI/2gnXfa2RenTKHG1C8
K1jMAqXEtTSrbDUeyjxi1ZITgcebN0VQK3akeHvJ2rtBkq3/OaflN3krP9BuIBinhPkai1K6nU9O
RlJ0tuYd29CNX5EAKHoSiRM10BDhU/FQXPLZZh4UAZ/bPmxU8CntwVhVSb4f25BKySnSuI3MaFiG
/FQ5vH2mFkJV3i1eFAJiBsEj6JeuWGiGlJt+p4YIYtj6CTzwWl1bbXPLeKnfXVPxlhKmSzlJfUDz
7BBjkpG+vf93QkCGL2PbIRbHCn/Ywt6UiTa6f0Hhza35nA5KI65g6fh8Owcj+7Bu7CzUCHthA6gg
IgVLPzLIWWbLKvn+MN3qovadwfUxeU6FCPL+MdpvojGVo96L/EUAdwnWmSTTJjOhaSFzV/FF64at
TM/guceynbxXEQo3p1piO3cLeTbBxxxErEC1Zdc1yIBzN7Q6iUu9B0NsqX6lhK0QR9k3XYUvivb1
0zgBs+7kq56e+Ac31wbeIfEnnTIvKrpoEZaokHl1TTjFhlJhPKpF9LR4BWZzbZpgudJKs9J9FYDv
FhWfqtDU6Fz9OvCQSsU9FuwWCnmJC52dvJKlt6/SBcUYhw+J6oRVASu7U01Zyu0S9+MGY8P8rzeo
asObJd4Cp0FP2ZOxter3Dd6ADnSbBh7UOIKe4lld7nj4qNLJYqlFhUT3GjaSZAhjbr6l6GYzEHlF
mmSk2Fg8LqHinT6YxdG9kV8NKlroEdDp4MG4yyAtuUSdKkyLn9sKKlLL1N/RiHSQjH4e9il+pbSD
RPWMEBX8tD4tVIsmUMGiLnDqAyYWqF7zlpAcl1lQHiQiv4b/9d87aUjBuX1IRv/HHkvlMrZvEUJE
7CzUHJN+cKuuZYqvygRLcaYJH18xvdVAFitZBCrffVk2zeO2MhyjHSp08bOQ0cJJnqi7BZvR7yce
9NfQXnNPR1weIZH1sZIedxUHQKNBtH+Sv6fkjxe2RCSFluG5Vbx9QiqPGDV8SyrXQS1WGtYHMRo9
6TmBFD/MK5cr7v7ELkUwB0V7xz/qcm83iW67e4bKqYg7ACPWSaIMoFFdgQzq9nn+LZINrjNLGgkK
KchyCOWqbYyqAOs7nKNAhYiqcLWtW+LA7fxuEltH6Fx3XpwrvOITVXubNfn1sn5K5ztjTIEVeO0u
568GYxRR/C7OURLfvxsiWg7eKccu3MccQCksxFU8EYMyLHHNDfzqRO+s7pZPXDEhTyPMlcXZov9v
Onk3n4oV8yslftbfZph5wlhxmhe3U4FlOFB3HZNsOyugnozhwycQrixiZMi1dUQneoKlLsllevW0
qOZF4lqf4c7LLImYnK9ek/Jij+lNDdJ7non2adOXNCOzP7iu7MrgBgh58UwzMoFkFVNg//jOF1//
KA2mzO85UHPBzSQ4pBj4QjUUYYGaVzlJdjboByfVQm/Xe0H3KbyAL50hALj/itNS7caqlO7wDF7n
/5z2GKjSg0EKFmTSUkxPJm//hb0oUhVU+uYMrYwtdndDe10Z6mse3d66v69hsND92vuz9Iwz4Kp/
ae0c/zvTS8+L57ZygzNEAK899CLRbPy2YZZy5nNB8l9Px5ZqW081UlBT+aOnVu4oyG3I6rBMZ5k1
MjvG8ZemMgP3tFoHa4u88ug2xlAKvOgWCfdT4CL1jMn4sEzPZJTMXgtvCU/wmx6Vis/qidzlqBb6
zH1jpjjLqbkNAn5eroZgYHON5+2sHZC0UyyT0utvLiJZveD/NEKGHilrZ89qxZ9wljNHalQ0jvV0
pTWNNA6tdp0vzmcMBKD924I+JnMf2ULK6DYOcizWr0ekg3rQistOZK1Yoe0bE/Lybkqb+nmxFydG
yDaY8ZU5m1gdQUdqyambKCakvq7wPLMUpB2a9RUKwjPWkjLnYj12DC2tGs+J8zVYDp7MEJOdLKbk
ZyvBYuSUBavjTJGF5Y+Vrir8Pwv7CSOqh9woqJohiIMIuzBhuNncn/P7gWVNSeKJYc47n0a4A4QG
yDQhzdGWZrziyHY9itQHmgV/KTIcKUqTJ3PeawZctHmPV5AE67KMLJxRjF5hrk3E6ILdaVMs9GD8
TaPJnejvLHeP4UgsTNGsw/wFbX/RM6NcZFU/2VrrF8Z/NhEaeJgiZSb5m4lqsqanS2igPHSU58uP
cbdaZh1DP7AvTHrY36+OzM5CIHJqiszBpgslTU03E5rWA5chn/FJPq9YjOSL8W3mBs/cYXzkBI/9
QlRVXqX+ysBFulUivsX/GMvbwglt4dgQu+YtgjbYy8q+vghCelSHEnA+45aWEXEfT27DMegHfyT/
7+Uc1x4lMj0NF/wsq5kW966qeMlBv+W7ycOJ/5Rsk/myuSJra9UpkFjeU0ClQbFi3NMRNNThXS2p
q+fwhMI4m3oi0iouAearBphSj9tnXQN+lgZEOBIb9Wf9MwITkjjiGt8s5gDE5mD+jINL5fVie406
VXXwW4QICdigb3c8LQz822YoIkgDfTDd4cqRtYZT3OmLGX3F7joDyfnyseAiFhrN8iQ3o1nw26q4
Lu6p4vNeAFJTNBBYMNcVBfnKtenRxWmEiOMk9ldOpAfFRJXpzqBt/JLNuTyip5XunPOyOyqVwCTl
s9WHtbXH0EvaOrLGcTtSL6/vhU6QBt1A39BE/CTFoNccZuh031wJSzejecYD5hDv8/3N5hrtg30t
kY33ck1npREiJfTV/8c10tNjBVXXW22W9LudBrP385rjkSvtHF0ViJXvE0tmAVEFIj/NLTdmqDoX
1HH/D/VKuKRksdeNUjRvVrmGAlhodi4uKLaPUVy0+rpT17Ak9HQzcg9uSUWXHERC+tGG7bP/tI0k
C+pqkAu/7Jm7oyRlf7LjmsV9Gp0P7KuK9QrFA952KlEaS5wMU9/gkk9d/XhM0kVjiuy8T2helk2B
J8HMA/Kk5P5pns5YnBrY+vYAX3wa3dtQYAAXJPKgO0RdfBqXcU/MaKmTDqJ0CRz9eY5EfzEtT95p
UYcyy2ClnNhTQ66twAIaY4c4hC2crrz9LCNxsOZKB1ntqrhOVtJk25YNumouxqrSbRLR6dPs6DhJ
8MRpMzHv2eST3a/nTZIbzR0Pb2S3tCdZB8pTVebJGO2iZbBh4UVbvomdoGhQAza13ffa2SEFR8sP
rWzatOojO6H134Oy0FuJTUOKV+QEQidK0qLE2aBJ/hQZj6wtadkYEMwgd7TWVGSHdNUjdExCMn2l
wHBUPLC6dGVdIp4Di2Go/rQXCvV3G8ThDaiyBWyPQ+dDq2M0JoweGRO+wwH6uhDm2UB+2NsU/H+E
SWzCKg1i8whbLNhCirvMYKUTVjSF4cM/O7JbHTQ5h9RtpT8GEAIOoAiTS3eLW8shIS6EJmwL0kUF
3+oY3FL8lVTnjlrW/MSB2KvmVqRCZOAqtugPUVN60SPVZ5T7eeSjKJCKSJYnHdcgPF2OMy8mgV1h
9WINpscict3WtzFu87+S2Qp8P85EsIwm5Cwm0s3DnKLxnXcLhRecToxE5bFDcKSvYi0zbC8XAkSY
B/qHZjSKp0dF/f/oe6LXZphdwnzeBP6sh4H0fnbj66nJ4i0yAEX6Hhvi0gME3Q75mN1bqffbJY8s
W4JymKBLJlvi33+w4+Xkn+7Y6wcOL5RXkIAmKs3FNcUsh7KI4QkOsda9zkjqED/j4FQ3Cdujj2Mb
jAM/d2jW0900xfYBHq4/L+jWqHpMOe2l7dJphkuAmGUaU88MyME8ZMlupIjR2UfnCf6XjIlG3wQU
EYZbuJ1UZVOKm6baMyBa0YkKF0AUymr4mreo/4qNrMj5eKC/kGpYPtYK35L4bW0VoT4AodUSn8iS
YdxQu39sb3ATVvLAbdQjuPg7NClCpWw98JDvTKYhur784I/yRtB0y2T+QgDBEgPVO+HFY3F4z/vx
ZJTAi5t9S8vwlOVsOVExvaALiDwaRbDC9FZWh+FYY2TBAR2kilG50doaFpyNXlkTpP0/T6YyGCxP
p2Aj55m9nMY1L5LsWAeQx1KM8ImtKie3g8ZEBIVmuz6in83HRohz3mT4tf7maa/Pxsxk0nEdNzSY
CAGWoEwJErqpDqAs6UhI7hTny5iJI5avlOpZZJQsI4HC+JvwaWlfpGNTRHSb0ScGrOgxTNaqxHd0
nrFhJYl4fU925UeO7Fx/SjREdVy2KVtDM0JALb8rFR+ZC5HmS+pPsqmRai1Ce95Xa0zmaOvz0Hxt
zBfkd2fO0MV63HqQ+foEPJiPsXCT6qAv+Idm7vX1Xd+mtVJ/qGHkFdFfaTkKVpOv6+ECQpva+ba8
K3opPlUxppe/vZOXzBEZtSyWphJc1e2VtG6BjrN415VCtT7dfeVlEDamAZz6+KFbjonfyo3wW9q3
JBGLt5+Src81qDyqL+XBqA744gNhaaqxh3A4kBa6c0c0F6d4IeorIDzZM7r/xT6Hd0qop7w0dAjF
2u4p7ZIdSZtO8EdepoqprcnDeBKAYxktSBTCbK+yCemgj4ttRw/5v4+kfUEpZqhyxKJekhapSqBf
ljpT1Md6l7A9FQYskOoJMhz5SDHsqQt0N13/q4uVa4Q6GJzG+NKL0CUeCXVaU4udpfd4/J9OZ6At
vMx5LK63q5Iekp79KxsTlQm8JyVZHaYjwU8SSvd48Su8nU0bmAfHNV+d9fnevmzIUBSjnFzgsB48
8tGg7tEf3Ogd7mSrXvlyG30fgOAfAQecZy+wRtukzaOr0O9X2cjgysyrYpEiRRv4tSOQj/IgXp3P
3iB7PlMp85I7aTu9RfMgSrCccWBHaOZoCo4NnR1ufmAyaMrwg5oDRxu76Kq+F3XD04WBnHwtjXam
FiWvZe3i5drvSAdMNOAJFXXaGeGCJUZ801NEPb5alM4ejZ0s99P5T6aPjmOzUdr1MZs6prqkI4D4
uaJ1Wu3zNQeHMIXZ+n4o2kEf6JNv0LurSWlKajiC4NLHvj6pYuw/1fN4EY46RrHbLd+ZLmZ+5uhU
uAXc8MGpkhi0kpmzrNqQ4Z0qkWRUj0rDVBG+rSTpXn6uJYWL6GtFm+KoracpMKVjXQfrLRoOOk4b
xbHsLPpwCmHEXwR8D7GEfrivHR31F9aVqpXvG4t2J+SmwTLi/zvRiO+paGWVxVxdgAbsLNIPDqIY
b1p3Blof6jmkkMqq6bardoiTbhuxA3zJxPI73cez/P0aoZzZpIptcmQ5f7W8tIwtPCY1rSzKiMDA
9aV4AouzDmyraxCAGtMm9QEVzlBIrfn3Lm5U9wqqkXUDcNfhk+hBmy+5SzFCOS8o6MZBu9dLCJOS
NNUeU6J8RP1j6ZDBLkHPYN2cwaejttovyIGhbx4YaWPlDWP72KIc+62GnpcQTaF0jMHm2OyJHmT4
VrUv+yKe/AFzq2FDcPmnzyMiX68P+Fp9mw92jnMkZxMYMu+lzdICXVvwhosbe88Y4f96pKwI6iLY
omaiQTXe5TwPM+kpnjK14phUjVSarBr/7sRxKUAcSDBgEvJerTlOFY/WXy3MrY/zOADs0DzDT1bb
haJNCGU+OAd2gKE9dXqALpys7Q8WkdFhsmPDOCCZNYs8tmIJ891PeXuRV+whI/Ky6Io8Z2H/q3tt
0+LPfcA5OF25DQGWT8g6vqjRZffvgfyIrShUJ3SQs1u0WEQc8v7CMOBk2NyYcL1UHaBhXoFOkt5H
n450Yo3xG8nAlM9v39XnP9YOVmciAYvoC8YIE+ypgMuEq738jxSkpRld/7as2bOGGQcoqa0nN7jB
UwCxTufuo1WBb2+WYXthq/1GGPmi0SocOlBlBJdAGikHCZ2GRSFyhPwjsCafr4tpCjgxS2DqR9yZ
cbcBa1TjV9poeh3/k2gNLQ55LzsmE0856ln1E19KDllvcwU+a8L0nNEYDitzH8fvmRMIiSZrjp46
t9o39S18FWyYylFf8MXnDGto3nHpJg6pc7R/AnjJOSkQEoomgahEKaK2N4+mpecGk8IiYWz2bFQN
y0kVcYV3cSKMsrxKC3kGL1TVdd2cQPt6btOUdCBI5CQ1DTey0x3maE1bWol6/YqbKG1UxQiVnJEY
PlUsMp17/Ytu8jYKYcAhRUW+LYUzLbefBbRiCXW5gs/2V+aniKxM3VIbLX850iOy4kwhnZaTUGb3
cZTBoV4jfEtwGsUXdiKeTgeei+LazbMhlStKVlh5qZwYW8FHXmqSkUncQTKzcK8oRps7oEkd3Zob
IAa+5/wqVbg2metxzc/HQRlo74JNSKYiviQ4R7phlqtIZXHdFMnHa+dddre6mnBaDuzr5CoQNezr
v2PY2m3xrmTqB1fOOAwRcP7MWSAPy8Nt1PJ3KMUpc3hEvTlirhuGFqyuhcIu7gwnIUGl8Sh6Ce31
Ptz36mikuGIJW4yczv4xTWAGMKUJsIM6GylNL7H5nStp9iozxkYdacnOnStBK0s8V0a25XpX3hU5
Lva0cBNpy7zThyvTq72/22afV/CQS+7FeY5tcOAh012Raa4cm55/nCmGD75Fi0siGliC1m1uATzH
IHZAxvbGoJjpXsavSM2leE+l4H/1bXVlD9CbbLturtwUrUWIvP6RWIJn8qBFkP3pfzjIb59Q6Skf
FyqHS+wiRGqNZOuHliZFlkjnCN3IcANsYoaIGJP5cDo/T93q5o+cjGNnt50gnHupqh7gcPAEORyb
8kz1AFRf+rRM+fju3Rg0sImrxGwbsbt+cG/gcgpyEjixS7CrukidKNZbRsUd0TT9weth8QISvCvM
qJaBk7RYTYlrn/Na/1Mq9Q+2Nx+TqmoO2BOZsFjLbikE5HguSr9juGVyfWvE4tHytnm7YgavFYwi
eqL6jT6FfTcuHlf4zQC4uOheuAEF2A0KpbDOqAk1q16AQqQ9br19n+83NKBEXEvWS1IacknYc0r7
0p6xykx7AWdTfHTsNzGHtzRrRjyJY79ni26tqK2HuCz/pQi2XuqPOvwwBB75Smfoj4KnumVyngXD
MLHxIRCH6xFgOeVgarBhvxOFVMNX0dwmgYihCSJlCo0xqXmHhxwcKGq92gPied9CKYAFA90zulSf
gFwyk3JK6uWY4Hs3ppdJwi5UlsJeOAVkfDZnAKSyRRNkZGr2jjWWBk5WwS/URwezZzC2MjfWY++X
uMRCxXqWPHB5hO+fchBUgkgOeO51T1ZrLr8FtcRjOrbrMWqo5fnY+MFz0N1sNTmtPLjzWoQgyGb8
JsZ4WFv+JhO9W3x3KjcC8Tp6PJ90c5yRp4NAP9BJ4MDi5+kNDmGx3gGy7b+LmjHcITHsNCPPrNHI
5z+zk34WcJ1gbW7JzGOuYuzK6TBIz8lbc8J0J/39GbspdLdxFUkenxo5hSqHYhwuvWrHbKN0H6PK
FaUQIH7I7ERojLKBrEiYySkkFCVXzRiW4TqgkAF+GAAaeQxyIPsddXmK3NgPjvXq9zY0apqbGFgE
TlhMOzbbEhv4AZEatu+/FDxstjrBdxG+Cm5fbRnDBDzlcO1pA5Wee2l8f8ln1Hy5mZTAErUgR5mh
oxtOOxeYBL54KVPSIofUYY2hK8WamPAaS4ot6ElfcfAccksX1sAEmtFBA6mQJT78GkrNqidOfzQY
GgJuK9yPUGV7fyQ0yGHcw2SN8a5hxS1YAyxokqcZgcfdWHm2W5SedxjTYgQBabL7Nig1Zl3WkTEv
H9qE6cb+5n6651ffDaK+LgnlPLzGOygDYgPAgkMw2BQ3/+KZ7njDndBPD7QyZaIfSSMUdcvonCv+
xyHzq6QtKTKRZ6pqOeUskWO9saQfg5YBnVrVk/Q+2Z7X/USXTe2zttFC75SpDgfwFU1TtD/9YNNt
Ldpj8IvX8NRNqq1BQ1DSYKCQWTPQimwo8vLuaSv5G+rnPPlVY1sIYvzd5GvFx+bOg9lABalcKMGC
O/RCn9oiD+CnQNzArp29amfhnxDYjuk3h4n5ol0bapNdU0jWYosQchjZgBx0GJCP8+v7kKDMWxOA
0x9E593l8UhUdEjyb+3NXwnttKlrjBSFvPVbKqnrIyvh7fSBEwJB5q1U/p9QxjmWxZTadi/7Ymau
vfMG3SYmGhBjDO6g7meEXNa2lrurCf/JRTqNbjbhmspmR4VxNLCLjUY0E4PsYoF9EiyN1hUeXMTr
YeOVfipzEpSvJ6dFcJ0wrTp2Zf5BJPJum3Y0w0Q/mU8xqYbT7w5kMkriDq6WT3OhXGk92prUIjwq
950lXVRl+V9/5cTFl64dUSBbpMszQGVn+2npPhwXX5JXDacyxO7hSmslsk5Gf1Kilk+U7NVd/W9z
GB48qLy6Pp556ZnoOkYeIxBRTvCNQctvAk4/vpTg7+bD6XwViRC9IOcAJScGyU53zu+nHSH7KFkr
sdw6MDesHhgTIjPV6JAEej7EXr3+Nm3AF6bQg+ZBG7+cjmXscXvgkV+VulmXSflASJl3rGI1LfPs
A3Kapldthu1zTNjZGjMGGVR3S362Xn/WKCHS3Zslt+NtyIxzmW6m2wyQK467dd1QSpLUkl/V9uWW
DZ9S21QQLnhn8ABVNbu1lR2Ytu1/zzxJGFngA5f1NrQ6cNnhNAaZht16XyQVqtESYpseMyIlSjil
WQFQMECFahvFu7JCu92hpcpJSaTCLwubrwf+Svuqf71kvZlveiKE3vSJM2MOzs/NGVc8xGFJ3tZB
bxLCkYcfyblUjc3XcKRJuFYQR4Sazdt/kCk+UMmq9kDHnTL7yBMCzxbKrjg0UXfGqBPR3lnrTQ34
Ut1j9SVomWaTnm8qnknvOkJR8J4TpzHfxTiqz57d61IRxCHaxvPYkjse5M5Ddc21uO6crEh3J3sM
t5o88PegEEcmpe/aK1L5TDN8qI0a4OJFJewAwloAtcuB8hMDCriAjZ4/ZQ6e94GYy7mA6lkeXDmt
i+alHU9T9HcEnwhvz5DZ9865fa7/hslk86HZKS5I47V1Botzf/Vv1qTnZwIdrw+oIRlePMY7pSFD
+uFhWrfGW12gVzqBXLhcxBkPrxuUtUDZySjAWO6MTZv6U27OE09lwKKstmr5A9C+KThemZ3C0hwF
YTQqZwaUZhg5ebObeYDe3LmZNWv3w/1ujdrvg+qRrAtA43tUMhEyKiXaHGn70oLMD8rH8a84Mw36
uwIS/HhbIgLojtgYNYcd7xf/4/9wogIBlU+nzrf2qEKS8/v2kPiOm25x6e7eQuK26Rky7sJW8Z3J
ZBaaUnLktcOnFAPK3tEnXSaa+TJnkT78ztZ1cC5vvPf7NZRDKYTT6YT8vAteNKSH5TlbIbUoGyZs
1hv5Y7vZLTShYz+vCKaxQV0swE+Uk9qS68shGdI1IWWCUejfCrCzqK15n14HgWnhHcQV4zyboTtT
bhKKqSEeeAyPZ9r9udNhFXaQLANZ1C8QACcEO2FJiFmv2Hn0irBcH+cXDgpFQzfBejWLMEMTpjZX
ro5ctOQHY528MFTY9+YXBQLuI9ykoMxBaFf4aHwz7Xm+GyEAwv5iDsBjq56O3yDhkUNdaeVS18Y4
mq24iif9JsCZcfAflWfoqVx6h5ynCA9xzABVGrUiLpfebS/e+qt4hEXcAp3N01n9EGDOsNsV7u+H
LaoO16ECMhmFjk2RM+8NHXOqNb1x+Z+TSVmYRSBX5XrXL+ghAvA9t3o5YJakKJhceKPov0CtMXmJ
J7kJKvnjUlNii8VADGY09SrsSIPKJmcAy/b5Wwn1VxeZlBelvMg11kFmiUHHYfgd8U7idHIgv476
afErsUSDy8/tzuxs/76HvJeMB33+Wp9kH4J7SI9w0W9TsxZyZjxWloZn25TYilLliMKmXsUPBInn
6rlXgioBhbyd5gFBYGWzDCVfRirauuE8Lxxhv11z0aRO18bljRSPzM3I62+6WIXzcDXi/gAmkY4q
Cr8UfQrJf/IVZ5jdtgyQbRjmJQQTwypoRAyirpIhOk9oHSxM23p3U3xSGK6xbFP66o684mExbogA
LvLHhtPsbr1tDRQeM1CE/mIEoZm7V1ZDm8QRrLYc+a5b5E+t3MfiFZKIM4nra2bHiHTGi/VTOUdL
+6nkU5iCphRhY+LtxIIYTHX/bgxpEga1FNFgS3Ulc8JFR3Mgx5D3rwNyOmxUdY9Gpn50NclqiPGP
XMGqZfmUddU0p7jRwUmxwE0F1gLZzGwQTVJs7vCwLinmIyasIWQXHaH2NVVWnEIW4fQ2Nyvw/hVZ
D1Id5l4X7PqwiDdzb+Bzj/EgKDWi2cxdSogmwXBNFjc/pWFizPlkWowzzr3sDlocvibL1xMMXlAf
7BIUoEh6Qze4Huf1wN1aGIxyJMA4b2E0DClNBP2WgwH8is1DH1wZUdBraM9Ag9McGJXWB8O0jS/X
ym/gBCTw9QE3T8exiWI1ZoVg9nvouGtcSI3Hdc6xXH8A81Gi2V8VL/gOZcuRg/yLwsR6oMiXd8xM
DfHx+Ss4BjVmE8IL9aKJfBAUaANdNa691SqD1DS2jNOlrd1d/MjfNEd9LahA16ZmLMaVUKD8UDef
zuB34C2Q05MidVTjicu4QBq3oCl3VYmm39B+1QJgpLYTu4CFUCWyTXg4BQ9JdI4a6sx5YF0mnEYD
jMMNIHurlWYiJx/W80PZeWV0j63MxJJw50aX4xvYqfJaQOG3YVVpvmPLYnY+XJ4XK2EAVwUcAKA9
2YQ3F65ynIkXvnoo3ppKA341fm4nfY1fXUl6rsX9Izam5DfDHhrS1mFQLsG5Er8tF3Vhcm2C4aLs
efsaQxWf0Utc0O87miJrTiDBMCYrNqGra7aYPfsRZpkx39gb9usFXdH54h4WkaOUOhfjGP6AlWaC
FEHmVKCIqzbMvsIjgTlFlWzWKaPpH6MwhHySUbCDJosxltXzb//FN9IeXwLG3mSvIK/3BYKfZvWj
aNWn9ZBirG5u4NKfQQLVeFoIkoAEd1nN74w0LUivQis7KFosYSyjz5nYNJEbEIUQ45srWVbd6KjS
Fcq/xNfYPdlSL6OJyrYFU8zmS9O3liJZPVQqvw3m+DafsI4ox+ACqLy/kVRkZ1Pdds5g/9QBAzcM
AUgCtc9mV1atS1PbQEH+k64h+ImMJWFUzaLr6S2PK8bbUTNiSxQksVM6L+A+buAopEZ/JRMyjjlt
fwAYXdb/vSb4/CbM4ujIwnGqKrq+emH22FboV7MX+92FoT+CM9Jr4QyYpru0tiuFh2QGixCXaQ/V
PmrndxcONzgUtnnIeFqytRZ8LqxlyBuXC9Nr/75GRqfStyH60Il7RXzeao986g8pXwyA0kalxfKG
AVQ5slZZuAwhCeJwblfOpxJ7vUMVJb639g2gUR9t47tmDfn2g0MqGwF6/tD59zdm8ghRFj/2Aa3C
Ie4gBPZmZIUjD/k/1w4rAgaVDMVLhbuuaGcD8Be/mPzQY+wVZclzDIbHNqKMwbatDFBIEoP45+YU
5uhji0elAFsEqksrkoUr+1hQIlosG5QEovBnW1UqCbXVQLG+ESFUsEgJf76rVpEIgDN5NhagqgPf
QVD1S2Zz3Xm3EofGHFnCOF6zQ+TIdsRw0VgLR0mv5iZdRxNNPxMWq29pcJuwc2vwrGO05limpb8O
TvaI20hK0Ml6h1i6eCsAfbnQ4U5LnIoMb4wKW1Brn6ng1Xsz+KMGDdNwBqVffiqO8KAvGBwM3V2U
DHKyutgiYvpxQ97oxdHMdRo2jifF/JpnUqVq3KZl/HNe+kFkNRg+odLL38WsltL0WTa3fNME0pf/
e30li9MKA0TEh+SPo5NrtCu1WdqR56pGn3OqVLPPg5RoUoC95chT80tlnqMAxs2U9oYTw2AttfYj
UKJCAG60MzllMaevPvPkNOPcMdV9+T2R/GNtFLL22kyMRviReRh4hFDVyTV6N3Z8wTnPNYHs8E1W
G1owONyWeLeLrdCaVnbVZwT7dqKZVk7zsgVFK3sLm+ZiS0zGm9Nqcn6V2f3nDGimb1v2otMW1qNv
nbJzKtCLsex5XDHgstitOOviXwewwctagZk+9cRbO6wAzoervxjosmf4R5784b8reICCRIBFxrQW
QvZATBjxEVg5eskfZLIETz/Rlic/Xrq0RWXWUlmqJkQi+C7JyEH28Unfd7t30tzc2Me3gAzAg5mf
Kk4TiMVbsaZM2zl1B74q53z6kC5TBV/gVTkixfPHDkECCDq7b0oQBkjs2BfnESH8CytMjU97o6id
sItvz3Dnla/D3ROg2fltR4WMhtsw7+Q8n1OzmZl7GrEDKO2BohvqLSGJh0stn9myFfDkoxY3+Zwr
FEY6UnKpjzMpZ/9ZoEJd9XDhdH8J6rshLio6Q/XT3+4JXY1hjTGxq5ovOmBBlNyJhSVKEZ8XI7O3
86DaUB+UhEDVjIMIyOslYd5CGNxtbdA8YnJ7XISyZrb0XIxFdQ68ZwocyCDx/LG9QvtUbobVTxoD
RcHfqPSOnUdZzDDXEQuQjXHeNgiRhT6fcK6wecpfDTznxw418lL1+fcDU1JM87SetVTrKGZKZ+TR
FUPQOGas7KcADCiH3Ua3bhs163X9kTZNXc46cIW2/liEcGcSg/mlwEm6nzMLvHDNFIqswRou7DuW
Kj4LZTzFNQOq9XBoxcHFK7I6WvcbmymLGUhpUy4RnKr8OdFFSiTb0ONgsZFH3ifpEKvimBqTYkp6
7ddfKycG2pHDjecsOuCgUiM4hdT7tyO1IP0u+BKvF2ar4YarcaOEKgbO0ZZkcoChOHCNXpHXXAep
jUaJTuoPMjw88PVsOXMyVz/LZV/TqAEN/9YzQNbhHLqogWxD69wQPfBAFQA/ktuDZFmuguDUtRUs
WJLmqj/t3UJjPtkXgkC4+yIxM+rgn+LqK2Ci9q3eYWkXwxTCR3Hvij8fYWUl1tjUOVxIIDU/tkA7
pjhkPRB2ihFsYjrGlEghcyV24UH/KOuP21Nhl051VPfjH77ysY8mjBpUrDdAJrrzWRVBIdeFoas1
zoDyq9zMUiCFj4NVSlMxUUcSYymnENSpTXn8bqHpCJii+9lI5NvZFNkSamvPFbDd/A0z38Kf5Qv0
uX23xqK7X8ngkXV4HGcCsqlyuBdnZARmZVZXLlT6XMcHWScqgIeTY8Dcp+jD7fg/iSZ5x/m9WsWd
/2LNIfva5zmsdxmpw9ZQDcUNMnc9GN9qZuxPm/X0c4vvEendOYH/jYhNp7ca2svW03odmnsxTlGT
Kk04vWUMDt1rpuv1ytBOuP2dnTOcHz6/7pPm7+Td/j3FJNrcf5IscxcAuUNFjKXJJnssQcfNU+KS
YCrtfl6nSYhhv1quKPSIpwGk03fqP/WNUpUD2lUa1D0Eb7wFvRmsFPLJAXdk0Uf8Sv4LbSCU0Lqn
BW6B8hx5HWZWxHABWCU3cJcrMa4TrpoEKbIEjJai9O17MXlK+0Q787kLcdPGLVs+Zj9+Vwrefirj
1VnNcPADKxkZ2KPuP+bSfYbmqFY8RxTgpAf4J7qxGGF5/V4lOvIOjXmL/1QBgTmV+DGT2pj3BtPR
vHGplWP1E5taUVCLotSNQkeTLF9zrBybqVDUE64MX1+YFUhqoYvH01Lr8F2r8Tj7J1ZoXbDdTBv7
wD+FluiRZDgfNtvobNzLtlOdztghYiuIjgXeoj4vaHar7XnmO6xcgyQtYaASb6Hj3xFlfPPt69YU
XbJA+dsB2QGzOwq11gWMKH3sgYgLLai1zUty1Ae/EqEUtBBdIt2oShhKIOElXUETUEh1LPvE95Mb
7m584euKSScKMD7poDX8OkKIjfRMModppUNHhHc0+K1EII4Bx80CUaybvnFvAULfeMBkiSFKSF0/
fYgH7PRv4E7iNa+mARFqW3N9yYX2+ayCnmkuZ0nYkPNm+r6Y/v2YVQZOZTO108AIC5IHjPOqmWN/
/S1T8zXRbrpP0U/8iIfivv4TTp+eTd9A8cfgMb4HY7rXn8MJlcBKmlQRdwtqswIaEeCi7AHU166+
53ORDF+Y6QZBwleqD9J/LoRzRgF9rTOYcuECWuWXkIU0y5bzuUc11t6uK4aw+jgrm7b+WVFtjmfT
OeZ5a7q/O1Ywax2iLXxNtnpIMnDreS28bgE/ISYOrJTd2uu3Oz0jS/4U3dNzcpOx8sHJXiFaRwVE
mi6W2XwJJRPQMUdGOtIMnCAm0W9KYJRZyGhx0qUI9CoX1QE2FkmmvW3uIbPI1QjLVDzDdZwAODa4
Uav7eX7/+DsBUNJ9sYqAhKEtDDofQnHx+jm2EaL8iOIZVeT1KJSHTKRJPPp33edCP/gJs/5IzDFg
c3/DvZ1lXulY7pgej/L+TlFNhPIqe1mTPxGxu26KmA7mCEId2RzB3x8PbyDNLz9BJ3fY0ZdpuPWM
wQpG9UeRcnF+iAoM5ipC8VXEZ+9gUjzGCuLbRUS/O7gtP1fA6cR1uKSFblXoA89kRO3jwVfXzU7i
AW9712sX218cgOXsoCBoO6EUIEayFd85FTSBFGJ2TRQITQeAnMyV6aEIBaPVYaFAeVOfZaWZ+5xM
yYfhGbi1Yj8/gUVR8ud25mNetWPZd1frFUKoUSxgYlIN5tw0bAPrdReTHuUXaivld6V1GHvS2rVv
Tm6JH3+g2bbZZ8Ilg8ettRgSxPvsBZv+yh2Rk9Ytg+v4bknbgQriqq+cgfqKhRS9VVrPrp0spUpk
Sk49LghyQMMuxX++y0enWVJ8PwyWMEq5/b3b11G1Zm0cXQ5UseMCRKdMn0PJCUdgqeR4HcVWCdbi
NNCeokQ+pp4M417lYGWm8n4zAAjRrH3HnhbMkVYMa3FKJb1naTcTzfbIITvGPPsrs68beNPYRsz+
DP4Uto0jaDPHSTPAlnFoVOOPlylMG5d7YW2DucpsrRoBKUF4/ANznIifXo1B5yNDd89+12lXkpr6
uvlEVYmwNLzLLc1yQpA5unyJqGyPqnAMlvIkEt1B6aTcvlTE1knwtUOSF2Fju5c3N8xKXZXEqzj7
xfAIGKH+paEC1kGh2XCeej3cskq0jsrEji7PlHh4PCudjQc8D3N4hnnhP+bFA4PIPABlRjLGxdao
+4N3LyErq4bnYQ9qj/601v3MN7XGZ9iQxP1glMKrB7vwrNN/fUFPIaJm7FbyqoHiNhQsvDxZUMYm
pmRGqSFjdBtj9XoDpPB3FdMpr47R3aICfsjF/cZ8hLLMI9Sgnmvh/kxKrbcNWco+B4PydJCP8oqy
dWTQQIKDvRDPwITGrdrQF+z4vfVpFIrOtxpm1H91TaD5I8QQM2se4qPgLG5I1Bniz1Q/qehRjkNI
SSetVGiWfrBgSAHGaNzMopfmswVTztojAFf1aemcYoZoZQe/x+E7s7CqZCcogqv/Fy5l3fd/9dM5
uyILu/txJEMb9EvXKrfLZDyTucvA7tTXZ5A1MOPYPNQsbep7XcblKkxL8gsnvLBvyU3oQtb+Fu/X
6tIvw//ocR2imriboTIWPiwoacbeYg7gDTraXZX12VGm01EU4iblibXhe0Coe0yg7QIxuR3gE+qu
iWppAfIT9qdJk/YvluCcbX3qTnzyWAVKLQUewbIbCs8IeizTaUgWYYV648K/wGTiqZNcELk4J4NO
d4wWIxB6jUBEdK6ZSGmAcMFg03LQIKSGu9P4mzLWpVSlzLkDL10x9eQXClAoq2CKcX/bjZGoYrpq
DrlZo0cKOW1vCEDFUuyBABarugxNCeEwkXSj5J0iSgvM8QvLGiAj0sEsN3F0woFt0k/UQ123G/tE
hmW8FLfN7jEzKaks2FHVKnJ3XXEqOfomL8QfFQKDrOHBlHEUfQEd4kYvr9un2rnVQN/LNlJv9InB
hzxWXY0MklhtfETW2azsPQltxBiDsPYYJ8za4brTBJ5ZHq6Zx33dweAOBHXoAhOe7r5wP4Z03m4D
ZkTB1oDPbJq7CHWs9NvtYi04EKRf49x0QF8H4yQJa0Gu6zA8cMyOOvorTJexQfXvHEOgZizeBf6a
lEd2eB0kWP4nYCV4hIqmGWkV6/5GSc38rVvtYnHMWLP4MD+euxM52KwEIUIq6Vykw15YpvkzbkOy
vvSoFXtr+/fuyQW0BP+3yAhm/nbVK4wyKlgilHlPb6lWGXdUpqKsGf+RCduaq6oHJDAf4N3p2MkJ
v39uZ2etINTRXI0KvXkhAq+bd1y7Sgwqk7LgLkix/pGADYIa3yKNDMTmkfPOhuOpCWOubOSlD9oq
jEqf4+Zbgoh58hlacFRhgyiA3fdOxDBmUgzOjR3uDU9nokpF2e6j6nt06CLRHQJ6p/6IxdZxl1Ye
BnhHJIaiT37Z41S7AjZWrdaCfsuRD9sh5IupDlY6N+9Ee2LD8geEhHt1fLxWWSkeqYzpQ/o5xy5d
4LUUnxskRA07CLs4xU5gerUHAk/8bBlu8Q3iKFpD7hTjpnnrw6IG5ZCe7YgcacYjvEmX5Ect9WW1
WX24ci5gVSWiR4ttc51fmL4mPpWUStYoVXZxk8F+1ZoT3ZZbbzefYbDbt6vjnUWNA6068Gxywr2c
pv8dhftXXlcW//FM5UMgCSDfKlrFOasmqocH9opsi4B0sgyblID1/T7oTj0KXYr82EtXf0W5dVTB
BaiYYf6jmyrcKubuKt9dJIm7H0qBmZEtT5vE+RY5axh7RAI2P6mNryQ7BhIk1JccOyMdwgJOsx4g
X0imd5jygcjbTLxy93xh9k0pHp+u5DkL5xYckh6K5KCVqGdKup9IGvpkZy8GTTIOLxZC6nM/bV9Y
4wgOtmP+rJLRCHravHv1GBuha1Yd2JgbI7vJP2S6wM1r+X/8r/d2NKgXuXArjWoJeA3oCP3EoQZC
TtEe8bKCLUHarMcgO4LGjz4fLr0roceROl086zm8909maQ1dl82XE6GfgBif4j7b2D1zt7pdmECx
xJWB6VERanvbvtjV/nRuVUQpUrg2/L4zGPv63Z08LHHd4twVnm9gqmQQCU7LDzsJA32srxnsut9X
qwUXDdyeNCrPDfu+2ZHE/+y/VKX3s+gWz6Tu1xBhESSFHQdvajSc0PbgP9dgPXzQ9IQ1On+kg1F5
KdONexMC1xPwn6x41NWbVtjdSR78ZZnnEtRiAoEWYEsNSJODsdyL9mOYsFLgDd5YvAqK/BhDWBDA
pwHAmp98jjhLTyuNMj8k8wYgVQts2n8HavD4Shb5qB+oErUPQa0dOGkyYQsX0eEqavD1862gAD4i
tqbB8n5Q9gQ0qAHsRgKO11NgxDuSQRmwQkQbXYR/XnOL48fbIq552FlRrGtJBlXPs0i1SbC3cUkN
EpujlNUiHlMeNIvSV1YkW/F4SJCuoDYptUlEnEp1H0M9G9sOlj6YO1pgEY6lAhQA5CqUHk8oP4YE
+6jflR+q14MXKqDfMSFyjvMoOcKhD/AqlcNCLlIiSDmSeQprulNRzSNoX4Ceggsae2nmMalE8sKf
2XPt0Tugcs52yLVwHSmyVMSZzyvonb0iVhiEBzFC+XATww4tlZyxoiPpkw8YO8TeRhZdUhKjVgmm
bHZ4Ef9bRU17V/xUrJKsQj8OAQQEG9EE/M8ocLCU7YqmBQao2HMAjMw2Lw/Amb2eqSjm5u0VBFVt
W5P1zPkuhSnNrlTeudjeEdD4ssovKSbPwgAhr1XW17eNLoodxcjV5sKdU8Yd33sQBFKMNA+swY+n
Mfet8K976cXH7fjdci2CfhyuyrZhHun5fCEvaetWXCZQ/feBjYTJRVZwFgzayeicSiBIOp0Tl66e
kxgo6wQPzwQb38qMvWJo7i3vKroVi4t5I/78Jv3X52q9ljRBP56hwZIYGFjrkzgacC0kt+H+7Cz5
yBQhsIbdzQfy1mPFZrYkpIEWkb3sQnepDiOrlOQ0GsWK/nV0Y77ztHpbLANbO1B2W6LfmLYwZBO8
7hb3nCtZY8R+eIz1H1RbI3BJ3Drg5qp7kQA5cWD8aMQeNNERJCtz+tsCjXPLdFvmpgBncH6E6H9P
+7ZpobxyZURx+W5yPjk7doc/Mt0GSqdX/WVtdSueHTOoYJUtK9gEaK1XvCnUmIk+4Yc4mbjUFv9M
X31S5s3wJG0fLYdeZfW9z9qWE6r/2xp1sdyn5t69tu18cyaNa3DAMrGaVacYGyIj5JTKnIxRWLhX
F9HP47Cl6sqm/olKEYHEEI+v6UD90IZ7ihefSfzRhNerabJjf/yoN8omTPLCNrDxj+SfIwupLuyk
p8oMSKoKlkIcIn62wDzQkaYwDZ8cQuQflKkL02FRSD4DwgAnjX1gtbgSbU4ENl9HSBeqlGblWY+u
b8K/vVo/m83YN+JtA1tn5llSQvKQQIC+tvJx/zTj5cGp57W3KF9N53gkB+NGPWMv4KY4D+LzEAv/
gpX9xRQnDKasONqYiJ2GBlTviir0qcXSZmvJaNh+QR+ZOsD6F+dWzCYuVb+JtS5d0lL7BIamRtOI
8ogkq3g4ngbzDwgieQZRobDiB15tPpXnFu4zT9AJexrEnHvTroBp7Ef22oNCNeROsj+jhpzdpO9P
Z41xd2n/v7NwRZ3NtBhvTxEIclrD0cfjvVj6cfHJzoB2Z5fjXggEQ2RgwFxDD9N4tIr4f7Goi1wS
2tFqRvao+D6lAeakINkSiqq+yHMfWRn/qpaiTpwpbUYvgZ12iBBnm4Hl2POvrCS4rH0QbrdJlrq1
gNIm2I07T6b4eFklR3wwMCFvyp/NiIFbMnJoA4SQKAljnRHV399Avfof/F2W9pe+TXYyMqxJcMyx
9KYY1MAc3xQEFw/yF9KBNMCxm9Vvy6G4ak1SR6ePSUFOzd0cfCOY1D/aLdbxUD59Q+Y/vfx50hwv
mG2+WKRXk4Mmh/i8vHKSyzYsSx3yUyEtM7ugGwxJrNbR5AtFAVJ19tuqo3N3QENUZM7V50b88Cfj
7nCjigydnDk6FyaS3uG/+pmv2YgB+gQVFzwFJDjX/FMcHNnMVbb26orBlLHBiShWb6ZZ4uMV4iv5
xu+AD4Fsx4GTboSSTFKreWFPERT11V1i6va3UTlAwJpwSslLlQTuGfcz0VwlGkK1QoKM46McNzk0
xa04Q5JwHqpp31MUt6hcQtxgTktj0mbcCPd+DUqbHHV6NXv1B8KFXHreJ79hIJiiDSvnv+/fd9H7
ov0myy5qywTl7O63GGVkjRiH8gmPQc60uxq9Lw+9ulpp/Ed76FJtVlgX748B84S6CLFT1obfvjMc
49QQI1ftyGwezQA2EmCvY9NDe24g5GN2GG3PVxs/sxjjZSEitI1+TyvoUUMHZkfvk+9NCdViHLjP
PUqKui/UbtjTm4CzWH3iv8ALI5zJYX4tB6fVJ6X57ajppNngsriBc8Cds6CxWvXzBWSLvHdsseHn
Mik2QM7rF0uum23HUjeVBsjzGXAvp4XE+Oudqva/8g51HpqdaCqbSjmy+ztA1mU5qUuE/zrH1VKx
q6ZHalsV4xCX1DIMyL76UkS7GTG+w2Z1v1g+8Tp28trEgzdjJzZ/6/AAjUbABhVUa4Okw4fknfuP
uTprgG3Wjw3Lncc6kTF8Z5QksM+qE6uooFfwx+tjVO4rjhMpp0ocXSkkfnPgVUcHPbf60UlA6bFZ
kbzZ1UC9fYyEguFjg+nmvjrzcrvlUFXUrbnhQSiV4eLUdrrdPKA4E8936MAQhp5yWpcj8dK5eFLD
jfuQHnNwYHOUE8Wsli1TR7h9f42BMJVSSlSwXZyMgCxC8lP2LiTazq0HTlji9C7h0telk3qMQjeR
i99awjAG1mGsLfgElczW4Kx+B7n4YOxid/g2SVxIHUSMSWjDyXxrfo2kLLQL/MKUdVx/Mnmi0ynU
Lr4heRfkbaairfkanb5LLolD4lK1ROHN1n+MAUL5XXXadsm7ElgUMWJiXsa+ME/XdUqiLVB7pT+M
jPGa6hiBgwjAtG0Is74inEssENT6wqLGRtXE/ooZR20XXe4LAWUgvXV1t+UxAAVbvUCKvQyQYvmM
7u8oKPAtetEu38yYgNS+VXfWXDStb3EcKn2qcXzozeDVFXqQRE5/mCJw4VKxtHFscjswXYzxAbGO
4f1bydlDxEKsRnYoI/37ZoNlkh5IG9Plcbk2wr+/0+j1BuAMlW9gYGbSCyb0OI6/h35wA3Fpupol
BiYCEx+8V73HfgGGnOxoSCKw2U7yzWJ/plscInpnZpaY8ineIW6k2UFhuqurdBLrBvZUFjD4hqr1
GmE8F5PGDoTUKflhA8rPUmEf7MmFQ6WRfEANqx7RyGsiBMNexf54Al3gjvNuzFNru2vZGOlVtaIN
LG2sW7NjJG4IPz8tTU32iAbJSl3OFy19IBNzv1V8modFuBnnxZG98yWGEk9LU182cjJ1ZD7rjj4S
JIBi9ou0gKw4Rteqx8lQRGfzLL29BFMo2X1ImhlVvsoMrwB1E5hTfcNt+Qt/6GrbPDtEPxRaoFeW
tjjfUyZhjjd9HdqsWBt+T0X8pgnVqBVELJNxvOKTk4YnJvkouaZXLUE3gr0J1evtaLTpjDS1Bfj4
qfTGzXZ03OYMBEGGemU4El/0tgMpX/ahpphwgAynU+3AAmHb1mAS9bGAXNiPeZjS8KLvFzUk//RS
nOPwLrpkZHPOuRO+QdnY/TIGgTx02ybS0AfkVtfuA5OYp03jru3F7LOmd7Obd3+Ejp4ZNLZ1QgzB
/mRIXfUUlqNEffLupEpJ3Rwi8JlharLxlfmzZPyP+sQMHpxpjR3U9meKcRXXi5+Nmt3vluq60LMS
m2D4NL/vnYIvZ+GUUTHuv0ItkV3q6JE/Pbil16Rq2BOjF4FXYuiNwfvwO+u8G1YBTQTkNTZ8/i6r
Nf4GhBCbPIoLw290q6+/vmpKUEcnncLddZqkhWg3WYQiGE+RzQ+g8fVvQCWuxZ8nEF7GM10ZwRtp
mSt+HZja3pcKJ/KnpIuSLzry83JeSx8RH1CREKiee2KZW7COxLNN5aq6khxMrMA5WtkQHl4/cMY4
wAgH1HhxBUd6OvGTL0dUFUeXT9qsXpPHEoeyMbeCyFMwJR/ykofgTiBYYTBPh23j8Z7sN2KprCyf
6wwCOqhXXFwad1ZbQdAVQe+Hjwf07f7TLtClfQT+EIgmlY9ByaXvbH9kdUfHDUPlKq7K/6+/ryEJ
c812BixCzsMF+2q0NSFhD+uukGqgtDlFMiBUTvN+W2ARheFarT4rdC4Z+4ogms21ogfpoao0J4B/
0W69ui0AtZSu5LGQky/8mJlrI4IDbtnCOmHE0kft8Vq7tSNCb+GOuxMvWB2+meW6sodspzWfa8kS
urEyG2P5c2mfADYeYb4VPjaTqJ8iDxgi7mEYpXVmhI1ZoLc/LdpmjATnhgVKRZ7ZDOyaBsrxxX7U
2YVkaM7HD+kc9HQGw30MGLULGHxCzi74RrjJfdRMKymKW/zwEOkRZQwJ4IclycGfCElO0TfTJE9/
/07a5ujj6cV2ot8kN4wN03WECB5HeFinhEyeI9zz9+/wakQwR8VNnEdYzI7Z3yomJBRMDPlS6OYV
OXedoFfHaCMGFk6jAH7Ztbd/mIgVLIXUCiEaNoGlWr5Vwug2B2Uu+qYb2NRx6T6/6VdG/DH3bkmE
Z1Pkg5bsnkG7XQLDC8XTg/+uePuIPEdrNoHGREofTjQInxOkH3OF0Jk9MHuX8DQ+fxD7cUR21fKN
aEUaK+T56l0xfkHfDXIoFstGi6CG/J/v2AxZoM2t0iEVZdtMW8Oz57mr99GBERqT+FPKtkzX6Yi9
H+TFgXKT4Cr1AcNITT6HdCRon5yx2C0I6vErawhY86BvXFBgLMyO1cc8+llj19RH/35s9G0dgPxh
PcnK4PKP3KxYkfNPL4JX5UDXtVWae4SCOeq+B5O2Md5uFkkLcby/YdMhNoBZFDShnqvcd4vgUN9z
JYDMjrq92SmvLMlNWX/12l5CsRkd4G+7KD5z1+QIbGUsQ5MxJE/TdatRs1on0RUhG6uOlDoKP2rq
dV2Dy6omk/5B603I0GlYdXcmdsinmdyscyq+mzIOzJrjDuxrnr2ZWaLOKC5Ue/Sux/qVrL4c4EK4
wVdhElmEGzE6ujDw5nn1FqO6lPIRAsRvlA4nmlZf8B4cwOxnqEBxCV3fBKmhOR2DSFZ1LdZoXA0E
qnwBMDdFFyBUbdSxFo91QgDrhb8EkN7AYUavlDtQ+op3047sQb1ZGk40nazW2q8RChcBkO3Dtwyz
EJL9NaMevr47lr/MXdoFZtLDwjslZIPOIHnAQolYy5A5CwIoGQRJ6+6SfgTNaltvmUcacMduazDS
GZ5B/6nrMaiCs1Ltn7ifhRl9mWCuOruk5AMPZKH/Z/4TPxN/x2qSSu4mMeCNHjVDwCelRUFl3cyp
1Mypf3sVJ60Q8pPijLtWKlpBYin3r3om5JRGqkJi33JQK7iHVZCxxTepD6H7LeQHRJovM7tg+ec0
WDVu1O6Zoagb9hRRvvDFpAE05DStCeAiHJSlS26vJ9XYd4XbqGfgqmtdQ587yWfBkRDnDnTavHwt
Jb5nMQDkq4d37KqxX7KXWwHpsPR/dVov6p88NO9UcrXcIaRMCgNhPgRmSh1wvvsLNMsMIQbNaSTH
CQ95Tz3szowiB2n3gGgWHqU/bl7tCwDxhmsDUgmXFFnD08yyu0AmSrgWsTiBKYxKC4FTXtQbWOn8
M0MUdOjelh2LaqDIYO0A7UlZTtSMjRsqm+YJxzZ7W4GUANRdB27zyA9jBiPJFhywuVdcCvSvJ/VU
v/eU1bry2MjGrXzd2cqiLiJ5d5LNJqxcDw6w7cFGGjwajNuWb7tsp9omzg4u4wvD3D6SmoYqt4n2
wB4Ndx5oo20r7ky3MwkHe76jJCV5iDDkPXq8JQ9RH1AO8PLOkcaJ5G2nuGUXF7Y3FovJaWorboPz
JSdZpMnucmFDiUmh9IGiAtc8CwXrk1mKHPGKHbOluhbgG0j6yVQujJ6ZOQLAa3VfF3uHgQuO7S/+
EBcNvXxUDJc3lspvANkht0+d5tQ7qiB83MWDDexC84RD6hOQ5FA2Z9scDdJzoOa+bnL68pMok26r
IMStz5dfi9nkSUa5Sb9Laj+wDPqvWe3ypQ5NFbDQ50j42Hrvvh01IjgdAiQGWFUIAFoxuPNaXRm9
/OhMPMk2vUhEpTH1FeWwCQ0TRc6Z0ucIGpVN0woMZkikLEopm5xcu7fw6AJgnO3yVdYdPSBuKMd/
TshAxDc51OU72fs9OaqYgz2OsPQHvOVShsmGD0u/hmvCJuekRL7Kf2Mmb6iQXa9ITzg+2j4nrNnw
vggs3SRY2RbhZIHocvGyK7fIHzl1GdZ8nuKunIOhy2tR+byVNCG5318KB32merMVuwQFn9EKTr+h
3RL8gb3w0l+F9mMe98h/V/Q8V+X1gbePPCd+fF9arWFLS2qhFJhHf+UgVGZAOdZVhInP5uZjiyW6
gMVvOkpZ7eL+sbWYJFDF/EjOpdqRlaF8fTh7+kURCLhxpzdz6pJNcVCwY50l62awn/66qbgyZzRO
Wps9Zd2fwNaPyXbjGBrrS39vpoufAzqIITeeJAtgWrHPNo8p2cTAY5KRLBjjKg3WXzgMTd2so7Ow
gycUzucM7BHKkOMLanj12Dq2UDki3ym0IUBsotJ2tbg7juf6g/vnw4nf0g/UVxtQyB4OELJ4Ge1k
l0Q1YLSZ01V2uVnMF0StKOTuF98lKaeQXbH84EoV0/ayLuobx33qR06oo9IlCej93IEjFfcw/DQH
fy+5sSE3H9TT9L2ghg6EZeAmo/pvwGzs+oCoc3U6itykOLH/R3mcMX51iamFh/2OKQaJqMgbT+Cp
QhjrWB8cV2j7B4xW9h3fZs2sPsatEU3RNnfKC6e3qW7MapUDBMWVU99cZN97r7CoHGReraGokOX7
OT6H7SZPpqiGxNwEJwzQZVokBm7hV1DsX7oPA5OPw8YP2KJG5lxR4WfmvIEZTd+eWI9faViO0IFu
QHqZ7JAL2aUJAEAztPVL1QDzqn2qRxO0UlQ45tMavqC6WuX4/is+hNK+NNFMWL0yHREUzexXQiEU
M0MUcQX9HnBKKxGF92OT3aOQ8KEW1i9zrccThjGTBGcxNJF+208UXDrggCbVdv4u3j/ydAJI7Yl0
bL5IO9xd3RyVd0mPBYktq+euFHbJsbZQxSF+BwAJgtaAnansNoIqMhX2fpQtIK64pMoToEEr0q5h
PH8qLMEUcNlVV29TNS0qjVrrtnSYHrxnXgXGc8JwHgquiYxXkfc/WvcDF7uxE+Bc3u7skkGKzy9M
zByQB992USswxhSypA2yjfKjm+QbSMFfJXpwv7Xr8OjXJrjO3kzjKT/8I5z1uxgODbnieyDS+QB6
mspPw7MuuvRGJhGdEhqJZ3mnR/uX1cBTgC0u+s5FqImkkqSEzzIBtw8Er1pfkBH7ghuUKr7JVL35
YYtgiCRjtAglwfUtRY8R/7u9r0E3BffeStZcdvB87LrSlll/iLjbZEmWr1pvLfmFWnY1ZurATNOO
B91nVdiQVIeUY35w/7sRc/itflpG0104G7zHzCbR/FT+iZ+65xxS1q6zK7zPry2JOkxxqAP0i/az
N4MoTlQt0WUZJtlQ3jccRF2/i18fr2egKv9vJZM4FKZ2Y5n1IckF4OmuqqmDSZrh60+hpSK9uzR+
YYTISw6WuzKBiKmzt+ij7Z1Tzci5YXwFICK/iHs8r/RwNidC8/Gru+hw/4bZshu0kO2RHRthiTsq
0isyphS0ODC3jjssH/FP25Tss2JgxzfbsITxVOhtBKLaYWolR6QR+y/ljGd2PuOgR7NkzsQg72A3
E6ulTXAHCmbmXil0l35koqFV3QcJzeYsvnoTK7rkDHzuhhSGeCy+kDtgT/3Te9VZjdBFDKAKAOD/
Ti3Fi/qucy/HJg8tGDkc81lP/cfO2Zsz6SiicNs/jwVGix+V4wUbzwrIOLylKqbFMSlW0C6UOtnz
1Kynd/ak7Nc0dTtLF1jVHa4whv/bEtRJaOKDEU6EQswN9Rh4/IX6sHU26Wb/1bZyJ7nyMp6s0QOl
nXD0q8fH2bXVEI9LhGsqdy8zaJGtiBL9lmw7KboBLJXnx5nnGNAKY5Kj0+r86o1wayfa5JnXADC3
KafMfRKzKBCV8YerJkiUyhyNO+784Azo3+p9iKB+WVysQMjrAUuKuOV4EZgS1skBBQzt+y3rNR1Y
LU2r4ZOoaCUqdnvur+NL/ALrPp/HA1DnxL/Ya0OzHlDnA8oDRXfUQ0xvMQ/yiyyi25uTxJPSsjoY
G6s4+eopnD8+Ju/mcLlkoN5lbWectvd5L68fOf6RiUJU8SjtyYJ2+dkFDNNqWtFfqhrtZ6pwb7EA
jFlZAOcQ+g5RQTg4QYs2mLLoBLUOw/hQ6IOe1D5teq4BmefZmDUOh/672N1Rp/oXvI/wkaXnSnzd
vVC5/3hyZ/T2SzjYOA0XAHVakg8+VwiOlQjpq5vRZ3p7hAlbIbm3kJSQh92emegHtNJ9ifCLs+rn
ywPkrc4AJxR1CuTHgLTjRAQQLq0kWQ2mRLBcPDBmliSE9WBhtswkC8JRB1a5wQjQ9PI/oRRlEa5E
+dCpJPLn5/bwBS9wT4R2NBCWi9zRGYF16BN55gjZIIO0onxx+wRRLas6kQWq0ZkJ0TB69UMqblWR
f0MQjckByjx3vbSE9OtM2b7sLZiWYXM28MxzRkbkv6wkL0cDuCGwK54NJH8E6p/6I1awLCzveo+a
aI0xA06awBxV3qqTBIzEh1vrmh9QatPcojUUASV2fXPvljeCbMwK7utL4zG4O1BID+oWJfGHwgjt
KtE+OMhWl9H/mlsXRUYSWuHhqKmD+7QaKaVfFQcxLH2+HgYA/SDyz6KozCqOQ+ybDJKArwyjbJV3
geSUb/5yIC8MUOTbTBO/cEehNQmB7jKm12HElybmWRtIzNMHoSS0t8L0PonV5Dh1m0fm8yDZq1HP
UQKBzdf43lpG1WaY+d8G4hF43BaJC6Q1hsMgNDrRHPCyIJm2jV3CBHVPoLNfryrk3u0nFC53YrOc
1KaIUu07Hg4zHu75PuXVzmHKFc2VEuPgEGew9TLH97rVokJA4K1z4oMBC7Ymyq8GY5MZ6/btF7Mb
lCIubuYFgBe4wdulZ+Tjkni/XE+Z9/6xsWlyLyho70MQbWyuvhogjzWIJLuOHqH2DowYGGiyur2S
EUG8VXL2jqGS/WCL96McYIi0z/0bqG3l7sWkEMDdUQNgHVg9plHDD1g6Gp01gaBMydhga3ej3ehZ
mw+e5diYIlOHcl7mTgWPt4d24UBPaKSxzMz3mDzWF4iJwNr/MFNfwt+5cXS+zIjuXkfRCUDU/xAu
gmR3gSLVvC0gE7Kp0ZQmQtZQAqY+ZbX3Xy8Od8gqLP1kvMIqWB42Yl+vBzCVOo25ub+AWIAv5DTP
YShDMdz+CD7+RrMYyxPD249987lFOa0TlygmJbRctl7Gj0/bXxtiirmRlL6z/laXls3OgMPmU1ey
9oADOJZlCO61OOhsWyI0yhGr8HpTBjcsBKu8bSxrF/KCYnY6VFK9NuDrjoakVtqqDa5eR6qjGO2M
oZ4DOB4Yg9UyFPZ3Grf7U0ogT6ceffXi6zDtumA0bQIpHUQQhiJEaoEWFbRJ/Gmb16FM0c58AY8W
+VRtywHjAc4zDLokDxJH7hUKrea0OhVziC9DGtyNkpcEOJ+HmQ3sQLkz6v5Ph0fHi2Nuvd6fhp+B
KpIdyooU1POAUmx6O9Xcc3TzPFwHo210uweFqHw/Jo2K77wMQpw+bxsGBRLah5lP59q0yylSZY3n
FG8CSjBALEdo4oTCKycV/orWUdwK7SCIdnU4tYrjLDVMLLtzWJFy6qRTk/OdYDLtm/CAVwVBXoDJ
PXs2aAuw9qZVymR2JAsjot2lhM+VgZ+/5d+DU3SjrsEYTOBayuKLJfZ1mkd2HH+6GaV8g5sDIiad
HX0YfKn9m/7Zzmxizr4wdxoXmqVA594KvGYLRmejK2RonFIxE3Ig6H9J1q+h+A/OjzJeIELNKF8b
2JaYNHv2EP8agtMrGumRtKAfjvS5CgGwEEVLEsQuUscAjRYjpaox5t7rQ9VzNR5rLBJhTuKgCw6V
W5QdSLUK4SvlyqcHCa0Qo3ID+QYg7IkBkiNS1bkbALYAoKV6zjI+mfnKLMExGAgrmF2gxM+ngRRH
p5nhKrSWu1ES+Ue/gpbJOvIPl79Crv/PqhOcUI9NCyHiynz1lS4wJAied7b2hGgsDU+GT2cEgWAv
dtuptWz6JhxQ8K8RWeKGeMqhzhiFGa8wssLreHAT7lBgiXWCFPPQlPnl9UXHe32V2T1DfBsO6gNa
MnFNEJBvQ+7hSeMXNIN6XhvWq/FT6bQihzPvfq3PAa8jk+ugF3CUBdVXojq1TIlwsxSInmCYu5hC
iE5CJWju1xuAFpFMQI71eCbDX+y3lIzioH7rsoMCCu9z8Ep4xrw183ku15jpX6UxnESULFTWCzEt
CBB6Ja9usTlyNw3Um6acynkNUXyU+J81c/Gho+AsSRzgJHDVKqnFaWpWXduf0l4p82/dbOtvJA2a
vbQtLyElDvraZ8AernQuBCD7MUnqwMlZ5XvVZUzYvFRmnVDv+bFpKTpJC0lwj9cgUAHz1hmdueFp
dcO6gBYn2+7LDB5TJAfl9ESrbUZwTW04GfIUdIF5FTIyoh7D0LlouDRDuu1unMc3D2yzQYCwYI7b
uMjqfFFUMk5hVA2LdAW67oNwljGvNHpsRX3FvTgDyEd3HIGRvyGeNHgOYGiEdjRGc+DeFA+DbxtM
GVDTQ/uNPVTm2ka2fRKcANzhTw1e9qOtCNQ0T7vm/hekfeqUSCltrycVyy1+iu60HlgnOMoXlRb5
lfABok2qn0OB2bL3t+typCWTHqEQEAPF3YFmd+rWfUIeU9hZrderKeW2NEgcYPmn8p3Fwilwyprg
K8nNyzCUQsH+3A6QDImGlhTpGGUNrSqeTSBaW7jhNSHXHdhVLazDiEJLGXToal09myEIk9MllCzh
eR+gIWBuAjLRTnzfE1D3gYed7OxhBPqC9pEi06WXS099L2VSwBGNf/0zsk0SWJp37VkZMIqBZMZv
FEs8FepeuTcINdG7OEqmY9XKeKP9xHYwFzQhqrjrQltZUzIJ99RIj8ysYDlltECegl+58xCAUs5D
3soweOoTcg0JnBvTGH2a5vwvvg0OjTPFo6F51eg4znMTdNv2dYG8SU7/6/Ja2PtnQtp8ZoKXZlOE
QCqjeqexmowz9k4uHqQkiNqK55Mf8/TIOmsWps3qfE1BgeOfmB6Ua8Kr/HotE3QjhXeEOGOGV6wW
4gbsMAi69NLXbYHui+VXiPYHjwCrd+gXsr4S+mLCKJSNNKiHC/DR3qdK6pFws5/MRmijNwNQkEuk
6tVdtUAUkSL+nEcmXePl0h9oHl/n7XK2aGtpH5emxD6PdlbrGl0zTD3aZOLKFbFK+D+nhUmyeNDP
Jlj5qeS1GMiX2f4ohRB2kHLbToDnL1ionvx8/F24qK8IJBzzqiExoJYiD0lZ/G65bvNgll93ZIjn
Ktr4U9wMtCmCK8287m5FY8qQAMXPKCRHBo4ly50Shv0eyiiROJgucqxQQYvInumeQ5YJRsbWwI8j
NSq49QpKAFU0G478kvb4XcTbCT/CkwwDPWvor+6AH+ueGtzyGcpOvb58M/JLEUNem2LK0eP5ZtVX
rWIB/qv9HNXyITQq9bZLU2vaeaSuvLNkC5FlSYbfcRrTqyMeyAQWN8IOcRakMuBLwPewKxtvhdLj
t4O0HHnrKBzVFAYyCVmRcv1r0u9SdMsemgOpZ7SBxtCuiS88Uk+0y515bF77aDa1LN5HBCd0rd19
Im0H1hZpCOyZo81ewKQ7vpEPlRjd6rsiuAUWwKz/EhdMn803kDrA23u+oaWP8J/wZphjD2V/yKO+
p2kiLSfYSG9lOl13CZLJfJFcU07qsrwDpMwX41sjc6O8uoUJdia3+8+SxO3muJLJ3ZQLVtfy90Td
VyFZYfP2aTKHl++fZYfvzoH1Zys5YgJyvXyyYUswczNoC3Tp14XDvzhrw5eHHxxdQR1xLTugQ+Fk
8h4jsm43AD6rM0jFTQM3ugMPIeMSa1zsq1zng24SD9LyHrXfdm/Ml6w08q32cppAMMpd7Eb+Y0iu
Disme6r+Ffo5yHFtFLv40QbXHzSqg3Ie5H2qAGU6JlYbVkNyEW1KSnnndoyP7Rty1RlvXf+cFIZW
UDfm2fsgSkY3YL7kgc+aEOhYLYIn2SlIzt01DAweUs8WQxEFyUHFeOygQ0nbJ0YxpDDCbqST0MW7
7VOs4H+QeRd6qBiTB/6hNE4ov2K7sxb+JRea1vggpQPb87Y/mM+3e4ZfqPVLhu51PEnLPyL6+etg
Y1LNg4dT+yco7XnnzNSVhvPhy2s/3VYhkYg+y4o7WLrRgYOOvEuc5YKib1wypAAlxJAbFmBj2bqc
bbPQ4aolAPdQr+Pm1PFtPkkmysWo94xXtwDsHDcKk0GVJEfTt2XklbJaHl50WuXxnSD6QL0fbZAg
W85fNy+rn/RoFd1Qq9p9uiOXvogG5zR9GghzJEs3q/B9AAa81Hgv+xtcoE+KyZdU2f1WHyu0FYxz
Jguy9lWh4geEnevJoqmEdHuMHDu5MQHmtMW5dg6qouEUfGQ2RWx6eMV3PSQf/5hlV1pio3VB98O0
cmg+9WOlSGcnChuVqkfs5LeO1gV4U/y1AOwz60z0z8g3Uerjvb4CGWTlPVouZz02Cq86Q0MSfeic
MYgTjhqRAtApecgRlbimb8KbaOo737PGOWracZWc+UEWhGcQZlL5BWlqLQmp1H4yNAWqSFmVOyNd
TLo+4yqLlURoSaUvp11J8xffM7yNzzkehwK8S8RCr/ZzvGXExiX1R/0e8XBwByxHU8+ffucSYfJe
ywdu4pOLrJz2YryHLg1U7TF9Al0R1Oefw69xndA5fRVdyV4u6x6flHrndQqVmFKL6g5GOXAqFMpL
P5J3XFlyc0dwERCQpVY97les0BIPYgh723cxOTk5rI6wcIOC/R4+U2JLTpff2kNWsRuPbU4KGizl
kocqzorwPlwdex+zOGOK7Fa5npXFuzG6YJ4JSCVy/KxNZFJSOeisP0JFXNU/u45nbWgAwG2P1GGG
vstc+FKpC8fLA8tkLBbbVSwMJi3H2lHWLOgwqUyWAp6vCCE04o4KuvpU+4WMKqWPEOUDu1MDLbNq
48TRP+vmcvy9eZJruvL03nH8Oeosi8LtlGqSV5wuqo6+3RQkRt3WItAvVQ4qTFvyWAq9RM/G0cxV
HvTESIBptFPBFG4igZF1Q3PnkwsrQ3ekzVqu2X6EMuShPRCWKf1eFXb8Pb3/wHbNhS2153hBBJJ0
xoDCbKkz8u5vyTS3ULVSTZZYOSNVP0wqfbVeQ0NVh4lJrLlZ8DYkskz5RKyBlnesWtEs/glusxnY
/YZZn/EuxKQJFdYHfaOBc6umW3YjzbxdnocZSdqyRFJcn+v+iEZTsIg4k9pZZXQujzyfKXGeu7+o
eEl5LTtExyqqjNkoOpthA+7DpSVYh9iR7I18R1K4HDCE9KEtq6SnWuQjRkqRX8YyUHsgNzV8q3Oz
5BhNL6bZrOGrtAq+AA6MTRyMBIYvU485A3H3SPMmQY79ljoZEX63FJOOMszkujP+gtYjZ4uqqUvM
oYuTi80MBO1WoqzxgX1qYerOtvB/OOHuiHvMVWdy0VEVNTd+3z8qRtPQcYsPWAtqj/UXOYrlCUzV
QOJLM8xo7S6S79J/yeYY7ccfvg3Mph/1eiRXLXeTHkHE5kGTWH60j/dcNjpYh20es6FU8ktEfzaG
4c+EKHXJ0Tvkz4+bsU4DtsRHnkRUTADFsxaSBeBHgGLPkXp892nGaylgtzXI+6+MBfrWUoKZ8HRh
TuGuSRURCGGJYEgz9MTCLpAbl5Gaj+hmpNWzGObtGJR1cpd1jqw91vkl2CwIDbNMk7U3szSeidHK
wJFVKJdFamDUxvfiA87vkbmNx9x6TCM5bHJ7xoUeAV57Tbe8hIlmU2BAJs/1hvUrl4B1PuSILwNJ
yPA5eTImDvTQmNTdFxoy5pueiYjJU7GVdwEIgUL4aT8eHKQEKYOUAmuorXVtFtxJY3PWI8b9r/zv
SZvqL49mxs+6wG2Xx+TCW4i4wIYxaRgvhaZcPhI1xfL8v08svvmnH+qGg31HpCCCMQB9x6ioxg7n
PXO5r0TflkdavvrqPYJVLvlJzp3LVwp/v2Yaexf3MuIYcsPIWAEuviE/K0t+diO8ohz271QZhv8o
X5RY6KoBXgFovQU0qTIHchRZk51QAf/a927wlPoMbTYxsMhAt5YsAGvFsc/WzUEBfJiDYMpQqnYI
0540VWSZmCHnak8bjwWH48XGX7sXTIpVu+QZrp/TYuS02OVdES2lC08076CcMxi9lhIcZqPE2vTY
zefAsoxWirrvUXHc2bBodYtVw85enE/OFB9vEq/BNnM/oatfybSeunSe3gzTstff9b5Ix0QZJ3vg
7idqMsld/YHPdBzkFqHL3WGSACyhaXzNfcepMIgcyU4BHv25pI4Gd6Ckq7ZtxKWWB8qcz6+lhHcC
1Kb3h9X9BC/LFDci/ahqHNL0zqyzeDEm7CLw9TVwA0THDo/JA9Y/O+OsGu2oeOTW5XDui5z76j/K
0pVnRMQs1ezNuxbTgepyD4Pq3RmmUNf6nTJ4mr/2RxMUXJrEMFNkeN9jQdI8nBP6e3zAk3k6/Wwg
f62c1NOx1mpCF5Ew3j2AkTXvkNjHrVfp/sJ77pH4ow7k7rxogtfnHzL/xgpayXQ54TRVtoP+Yqfo
ldkRIPacenkKIiCGiXgAiyFRqilFDgIRxhAG0q73UtEdJg6J16gUzVX0dQ60QIb/W7YsDgZNJV7h
vVeIRnK0Tma0M711gld4whwBZQmuHUELlwYjgX9EZiH/OhoxjbV+fonng2gm1auJzzgTBjTg98m4
gla82CWwgSJYhUS3UzZfU3Ff12+hvWT3eM061z0wxSioJAEo2XsnI3oK3xQAwqQfic6NjMmIKBWZ
zeil3QkTcRwc3ANoXmf69mxFDSVQPCPOrVhNFdN7oCgb5dQs/b3yS1DanmQtOzKX6X70mX5Q6i9g
y0m1qVYy+u7WYbgCvwNPfcl3ER0bKjX8QPFPbIK/zqY32bNK3QmOrLzG6PfLD5mHfPFPgBOXXO8x
BiG3PZ6pnjBJ6IGZWAm3Qp4mcJ8H2GjTua7I4xQt7G8kVETcwKdGWSWZdYghZWU4C0T8g3u1hw53
QCE03nhVeJoAt+ICGGV9NPYV/6fl5dFtktHw3A6seM8SkANTAVEYV+95KNjfnXZtcfltxEh8bDIg
0pvxNpsDrfBzMGuIRxTsHSxYmfGcHYG3S4umyq6WilGZALytHdXfw4XO8pG02/vv0DgGZk4TjOX4
LDiYORf07o/Y4N79yZGbYVLxaEli8ov+9oF8BibzQ1Zz5LNpRds7OR9ypXRTGxfGxLKNlo/c1kc0
vzSVtpxgjZf6OFGFlP3pLgUF5nnfzLGgjBfE4VPjcBZQPdEBdkhUniETS3rr3G31AZr9jk9Pirn3
VmacGLHVVdDL0LzuD/ohcO32fOZHYZXYHOjEdHCunFeqQKr4UNubrTTnt+DP+LNFjGSZvEFjNSbH
sAxgiz3gxDu9eI0oLfwRMlvu2FaJoFXxjMmAKI9qxp7S+NdyiDlPjTgX/0heKeWSPwLMts+d3Sxg
IhBZKb8jBf8oP22D69YQ+1H0IFedEdSp1JBwpzHx8SQ0WfF4sRocqAVAf9FETx+5LcNm6YNe9N3b
nmsfTtbhFUdJ2Ncq7xDayhfsIaI+g8TlKXOoujnpePMjkWo1SCxaFVmw2zgciO/n2MiLFUjJq7J8
ksc5H9p4zXSTBz9ZJZdUz/LzN4q4n9oJ4OD5dVX/z2r45b/LtI+Jxaf2b7WgNP2zTa6hIsOd2Bah
Z5zgzbrKy6u6bCsvf3W6pNVOc5xXL1DkxYiKa6OXUv/Z0Zmm9CTMEdawfagLyzU/FmPe8IvBigNY
X+2alyFkPoAuEETOXqCQe06X8F+uV4tyu+yqHtZl9qMdMYG2CTQwnseG92u5qYTwhk8n5qOCgT13
JjdVStBiJego/IpyOifF2Eo/xCS7bDb6UPTbbvOKnuKO8SXSV1mZZex6bSfIbLnwSTzcq+cH73zy
T5QtIhjtBF61UslngB//Cmg4K0dvfutZETbaxmCxwoEGb56VosSYRcBZcwrVJSWdQKDTW0OMaOIU
xjTRzCYC0g3bSAAzUfMx6k0SOrS+Fl1h7i9yzitxahAUsWBtpGPK28qdVhHHo3fJUvRnKn/W04ZR
FYXD7bx4HKAoz8DsK++8dW+seM0R6Cl5SPqgmC1jij4i71J7pBR/OAxXX/KCAFEBY+GstJ6UXPBc
dPtzw38rSDCEP0TDr3qDj7ZLPhaN4BTe4MnjBmmaxNd3Ys59wf4+3EOJfRrAGX0xbQzccerVTX6m
++FgkBjrktq84mw+SXOLQplK2pavLA4HjIIfI+ux4dFxo76GokGIlB1JOymiCKU8W15ukVIEFp51
0liZEjQScjQs5Lfk4SoenJwCO0PlL7/+00Ui1HyyhRY4CzkKNUqfIwFv/IqQgFLGCKdrrx/E3/fw
RSdkBNZYpGK0ZyyhtUt+qe1CbQvX9uCkfKcztepBwTUrjZ1sH1fiiyMmdvEL3NIf6C8XQP9GahCn
/dRkqr6VZ+AMSLpSKMgBVk7G7MLTl8BQERL+I3k0XiZfrA7eI8KCLyoQsfTVQUTIGqfz/FLMh5nG
sijKnjdxN6W7SYN6SP9vJw5n1e+me12qEuSgn/I7loY1JPKtOkYM7tg+GV02nrsUQ/UIRTo1DBNn
EP1+sHUr1wbYFMxesElugUHOyiAXheP2fBakCgmW/+cUIAe1RqzFoyeUBuM34P4xe9T1wn4yz54W
k07m9V8uugyZwZEP2vJUSpRb7RO4XE8QNuph9Z2YS/sCjKcY5B5SvTFYrlW5JVPhbng4VxBxNDaO
/6Mv4HM77tyUu+lWbf4BEFJ9URpe/nwvAWxSRUqy0iPVfjLI/SDGTfoUrm1Ec/Q8QX95MYirzUWw
VbGlrh5jQNhxzgvk5DPmDDMFNgYjIf+nK4ITp5SU2k0zsLoSkauHsVHuXVcuYTpjL5RSXeiXma1g
0eECVKPzreGqjPc/A5kKVNxZpXczM+4wthHxN4QFA5i7nVN+1USwnJvMZoFBSvtywajpYqGeBNWq
/Pn9CF8phXyxjvzXH9Zkkh0X7xhP/kQToDUv2RZ2YFpDu8PmC1mLvMmc8GXTOJHQ37Qh6WAkr4ik
zIbSKtTJt71snw/DJ6E8zN/gh9ri+KH5IY20XwiJ3qAkJ0XCEr4EGqMmF/sHktyi43juFnZARCsU
zRh179crbeUgWo/HcuoDypPI4nSRjuco5zxImxIspStK8gQZwRm/TZ1gHOxbyeDbq+ag0tzE8Lxl
A789oGC6htbOTKhXZQey8XtRRw6vG5ripCAIPFxvQGvrOFav+Um8sehYeqfxOUHnyN+zSMEPMHOB
nlxpKpUrCji9AEvqNjtVohpmqGMxVgKnC0Yd/+yk/VVAIrsSxpp57k8XsRxa6M86L5rdU17mPVs5
DhEah4CE1jO3taLIbr78SwvdoV6F0e3w8/O/MJfjLTMfvDKZlmwr2pB6DGcWO4lqML6D5O4BBBHJ
XVJrX4Kbv567+eE2BRHx/iklKAtjqTeY+ZSaIoGVgWIpinYJzYPHOEdwGPcI/kecwoh8sI+3Jdh5
ir6GPBdan+WdCAp16wP0fFtyA+pdPKoZjbTBcZcsUqbshotqNzmYqHJPz4S2vB7q1DTNLq7YHEpx
/5+Il2xrYR62+fWzDIcrfYqRf4zDydekLzRYTQ37tN6YS6haOnx2wrgaQZCumZdFbVO3V2ZeXxbE
Bgm0cB4vtqGF5FUQlM6cl7MGMy23Hda4UZ4y4PA2C/kEP7af5krS226ArzuI/dcJ5ZfTZhLriE8C
AQqtztAHcUEYmOh3/GLaURjodMicZeor5J53tPC/FolevgyKH9yC+jFw591R3MMjQwvPGhS7iGcB
/frlGi6c2yKPKHmxS8iPTF6SOV/lmUMpA5q/26MrmDNDRW3m/BFl88t0RAOexZfohUomRF25oF3M
N2eG9moaIWYuLNXbvsBPw073oQ0xjslzjEWWvzh6Te1KZWo993eFdPnApqn1IExVw+oc/8xkSHos
bsWVYt7LoVqudm/mt3Zum7GeecxWuYtQThb7ZdhQ/NGOU4kp8+YntLIOGqEQLdk/i5C3X3aH0r/w
lyux4JCSVCr0Thoi6fhQxOk9NSudyVetmrl0qIm8GChrtnVktspP0RtLpEOPGzhoXuFPsZghN3aQ
Lz9tc9XttEbEJPLrLnK4GSUuRQ6HBk+mCTB8MKnwFXwrTpTtdsWjUETjF1GPTRHc4i8UbgNG1Ol5
d1TE7vz4RTF7UcZiLIafSptoR2r+85fYIdeMeWzh/jx1zIA81gWZ+c9KjVCPOs7/79171M8HKClo
Dtp2EXpScAibApf/TvYC1vuylSx5nq9lmfQOxdL4IECR2tAdawQje+7b/onvDnLj/S1LB3lHJdeY
oXj6L7nR4wDTN7ifSl0rqv64MAwlRy3S+/BaKQdhGbfWGn8V9t8xU8lsMwiZelzrQbPvQ85vVyw1
/LVmqn3HaXYky5GsLnmEwu8LBQ0BUjpHbeAg9P1zagwcCKHLKXgjkQ8j+sgP4CrRDdzVkgj0Dqsk
ojgcH4aZv1htnRSe78OgahU2caXY8rQkl2yQf9tLa7b72sgEVWNF8IIX4j15YQLcj6Y8tetUvyD2
ge3JMvDxb0jbZwv4cfhMzt7qrev0gY2o5EnxRoEpUIh8dlEbKBxp8mHykCf3iyyuVE6z2O4ZAVAR
TP68W5qPjLChuR3SJWjTtsGBzdDgw999aAasAzZVI1tgw0cLPA6sV6EhfmBG/S5/R/DC5+N2382B
xYvVPxxw7WIgUXYcr8AsscnM2I8gOXQHhfxJBAdJfT875o+0USwQdS3+OSsSrT6conn680yn3Vpq
Ml6nOi6gFOCXzmxhW2a7M7VLD77HRCHcDZbX2iDPJAe1pAOs4Td3ft+A6GCiFggwm49hjRIR9vGF
UH8HuX0O9WTK4hQLnOSLfDxp6peMZ/a4IjIynFzhgaDlhShS9EjrdgQ959bxXGp3f95c5o1dqfMh
2/QX4ulWtQudj91kINcSND4mMagmWSrYkcBczxY773Pqtzjd6SGmH9gyyls8fPKJn6sZxRpoRo5V
Od0+Irf3h83YNIoeIkM7zZlvxI66dCQzwYUSdo4a6WXwYgzUZuDvhc7R4HuGhAlDq5De61FuPQQs
XdPJTK8xofbS5HOtzuuUhRz+w2LoTZ3wOeM1T73VrreTDnKL/huy1RsDWNUAlNmsvuBxw3y0zCza
YQjewJZAU6XBPXT13GwLv8I6id1nSHlFqpZSQuHCCGThS4CE9eJqpYLW6ZPH6/Vw73f2ZTdlPeEl
KGeJMwBsV6geJSb/Q2UnPQinN3cyUy5glMBVBjrPCKWuN1mcpUCRd1gbidOv0cO5AkgphmMy/fxQ
l1xNEuTgfyBNlAwMwnQleK7q6xkOluSlpYDf4vxeWL6YLx/reHYKfmmLpT8274fhgWwWpJ8V7g8v
JF3crL4tOk6JwJib8KGiPRGe6dhwt9bZ6uswMOKleKqZZBesr6FMGA5eXfVzmzCYNDQSor2i2fcc
vdh951oNAEyU36w8WANj8r21aGJiqmcEwRVH8JjyGfmgFFfmdcKoL0JF8Is1dUrT3G5yil8lDe6x
eTlMxes877Cn3abb5Qpi/z9OjZXTT4rHYoCHl+23/JuUbjt/RJFUHzD4KP+EL8K7Mp3l3NmmvzaY
yTSCFmiXCjHLrIB+9pzBQ0tVcgdhYdszxYOyhYPLTtCn/aksVcok7ta4JRXlJrLZ1OB4szyKXa7C
UT9L2aIh1rPJvY25j0A7nXrNn6IvAXzEiUz1Rv3mCYIYYUPZI6f/f9vxrTFJFK1jPq9ermEhb+6T
X1Mx/BCaio22MnIX1GaPGAc9S7svuNDP1g4uAU3qaCafCXxWoG5Oo+D3MLu22ebZzJ/z8EwkK82f
jyNYec+IkrzrvsVIQUyM/9HPDS6Ekxpg+sQmnYgd4ujFflhDO4fUb/eKNMNFTvdUuTIEMZiX1oYN
zvv0QoqhQ1OiN54hSgz/x5WDw2U2vTF6unbKtAe9wN13dIZa57thdW2lmLPNvewqjBir8jtVpUH9
uOD19n0e0ozUQ447vG0xiwiOFLCSEdARHtsWpQL5uDGvLZ1DExiV3mpNgi2+Igv+cy6vXG8N83hl
i8oG8tRX5DmB+5iITTsKQ2LUcPcCFbv3tLRtV1LXMgtUc7PYxV/VvBYrvG2cK+Y6HlSGZYP0jNy1
Mo3X9rPcXIlUUnXIh5xjpDB/OSbHFOJ8a/Bqd4i3WzDFpMDVHgrcfu5fjJtXxgcKsdS+kqmvwzX+
q3WTvi6ZZtvMTJ+cnOtePA1YhQUWDT8+zArPLpj0lSzI+VUhFF30xZt3bdjSMgymMQ7esI7BpEhF
li7Hj7lBQybtnJtO013aqiS98K6+vaPqQmi7nABpP9PoCoLdSZ6DUBeT3eAqVwh8OBEFEY8qXPy/
Rz3H8dpP3sLWff7B55BP7s8UHI1FuoG98mTma5Ty0B7ulOtPPMy8e2awZQ94/ZloRXnBtup5Paz8
oxuNaHcj8NV0vjpLUUEmwdMxOo0EiXAiHqRMGM3ku+UnWGDlNkloC/AmlujFdv5j+tsbJKlrL1bL
MeKDdJKXKHwI2TRiQYH2kbzxtoR8pqaJU2Q963yx2V38uSBE/Ib3f4p4/NKFydEu+ZKRPM3l3uS9
7e1e5tBl8zDYA4v7O2NlaPN3CMytmCBSIRkNasjTKC7RbYzyAbJvtzPdUnyKIUVAKn5s6C+7fsl8
UKUVegHjAicPB+H/6Ljgago8RSf1K4sGQN+QgDPQBg9WiB/i51yM5txCd4gvkiN56RPewmwnaPnJ
Nf1iWUHGdNwIdg8EWQujW+2zJgo900GeSSAy99zjlJwP3Vtrp4EduzQ7rxjQkND1MO7zdgMbE6nV
2ZwXcqDwS9nz857A9qitOccSkdBYm2KSdyhCszaoMq1AtFa3yE5skxlxDhOHKoQlglbX43FP01PK
2ZlmJ7MkNG1tYZYKD6XUMAFnpgdRy+/5G0ZXy9rUCvE7FlSqWbj1nLjVZdADAVs+UFezNb6YVeea
tf9gbxcri4TzCnQDfYFTVV/pKmY5z1Q0r9pRyxqejgWMtUB4nORlLSOcsJkeXKUR1CvnAma0/yZL
eFHIahRgFItu5yR6LHyHiJooTWKVkaWOnoW4hVWPv03uFCMhK/VDttZqd/KzXK7b4Nbc4hfrldHd
orwtUJBp0d/wiv9bu116lGCr28YqC9sCPCz6KplBPszjzmGKfXDdz8jfAaNGm/6N4pR2dYB7m7oT
dBkDOIayY0CSypZ52HL7tohR+UG66+0P7ZtDdjW8SxmJ6fhUfVsgUWO33G1Cs1FJtPDjYFsodcqr
WtyWjXnyvbLFAYQAMBsqbaxBLCMwA8w7u6WTKLn0M9vs4kHSJFAQCugcJv+NwZO9sz6bfbD0oQuE
wmAKI8Ufs4iDmDzvPqjLLkxGsRVGbybBoeb96p7k1s32gbC1Mi4RKIdW1onalUQJPr6ncshQcgm5
aRpMG/gkWJ7QIBVxInfUnyN3X+UIgr4Hx6n/bAvv/ccmdCnP2M7NvqaDLXjNzeHhUTTISAsHc6ml
Q4ivPg6azqZa2UzYAD+etTHGP4iUwbSUbJl1pxZ7J6qD3VLPotxodWSpSdsMKl7MCUZZg8KeFfQT
z9Pm6ANXiP/lMclvJBppizJok/XtJIDAn8o/W4KH6leH7VpUtJnUwNpnmNdL8uIx4F7Q+vKyrHNm
t6dmGjGx/kICOyNgudmDfxSP7Oxs/L9QEWT+GrmY9KThv/nld74K5yz77yVvaHhL4gALpUjFF0Gc
ORif9V+lk1zBGiyov1ZkpZK1WwD2p6tjFkI45HDF4q+Nr19ClHCfUUeJA6coeWAliqPDbwmEJxtW
y/ydqzCujUzcjrrwzRQ7vU5QfBwhaLc7CNlDC4b9gC4KSFCyQ/i9dOFRkvGNoLwzRPcJKvVYNxwc
mYKEZYwpuOq9tiYTsohpTuJptLOVhpbT7wThWzge8w2BYFlMIglwmXcFP8FvcVdz9vMbblQ7TvnC
wj24QpZVXDBnJZXl0nBu/M+8iPPbjZEP6yHSNjDi+jikGGX8djTiO9T0AkqJ1NwylDdZlysLgnM7
unX0yIbHXmcNDfSm1dc/sRNNwLbeVix8DkxKCXPwxTQWOMAdJo7ljJGpMiz4tTDq0FEeK6nzRdfe
7Hn7cdlYHbJI8sqBnPtGh2mndSNtz3B/jui/EadAXhOQzHtFl3sNkG7vUkiVQIUZQqTSqC4s3v3k
GQVdBPFM93yoCqboqzCs516TOKbjc9gXgBKkBxuiPzuNK2ue287rytztwMkwS1FWuTBHaRbbifF4
FdHvDbaoBkL8mGcfYwCN1Srn/L8EHHamJApwrHf3+R5DHgHxOoFcvO20sofXAhl8QDCmN7Wanu82
BVtPupkvn9UtF37Hp0ZBvAkfRm6qVs0MyRuyob11B6qdFBiSmCzq9uWEdxFS/I+cqikk7oA0zBlv
L9T9+g0oKD4WX0MmSjMSeDE/8arJuLgXXzP3ZVae8QPn73kQxUXQSZ4ERNv7d23lpqehQXpdkdTz
yvdDbqWUsvmjMHnk26kYx6PfPrVX2k4L43fcUdscGKzKcGa8cII4OqPh7C1lJBDqnGqU8zQYVxpT
w4CuSAjiNgzuo7x9Don9KwrIRE+xFP2ZwWq4af9C24mIlFq5vfnNNpRG5dynh8sv5W2fXajVw2tu
SE2osnV0gPMZ5MWyyOhpMyNgEKpVCpaRYCANwdqqqljK0pzZKCULyfltel+hQC8d6qJ8O6+oiRNz
nYOkz5Z3M+wNNGG6bqrNG0NHhr6w0+7xB1Um4IDMJlqIkm0WXAOT1OQzAJXHyjZYydGqs/nRKsfN
jnD5lDEHnFORdJxcdzjErGzloRndvs2xEntVmBMxL8Ort0pwESeEbfifgxg7+79w2zxJ5LCiQzqG
qGuCy/tSSlf/e8kbVwRPlHgIDLcG3X9u9raGWpI1VKUpWYPOm1GX141n5zvwM6D56qiW/GmszDuH
+rgkeltBLBEujeRDzIt/AcAsNcvnraSTLaxkVl+6Sg3G2z3/3BI1It4l7hyW8qEkqgeTqB3iKuHj
DAkjqzPCU3dlgv7LXy3+uW6ARtMlYG9qDRc6reWMMcbl4IIApFyfe1jIyTyHKIkP7J11iaYrwPQN
wzThdfmb9Y0IrbfM4TXfLw2xuU4AITCPvsOChAf/NNfzr7GkGRqVfd2hcIyhnK0hATI5T5ALoLnA
bmrEa20vMeQ02KUxd/sWuF7oNbPA3FH1Jp0pNpJXXIH/AroyPxEoNA5KpM0uHMMUaoWIq0O+s/Un
6LxtJ5YVK7EFoEOZSWdWGzUMZuFfCr3My96O28hQKd+0w7o7Dzn9uWGJOZZ9mvb8AD0zg3MNZSiI
qIoJxkI8WJXvMTQL0LsACCtwzRq0mQHw+LI7p5q3DR0B7kuNDQDPn3xnY7V5U2k0Lj5Qvy/VWy8y
UYt036+EQF8HngrsYwlLj1xQnmdhBmNG3lxDyxOJyrYW8v37FUzhlDqfGEg1rAWAIX810JLnv521
UrpqP+3ImOUlZkGRcicftZcaOD08TnJLJtL4dPp/c2TqHwjbNBjq1vuH5uPlNFRp3ovuKEahGBwd
ZpxIAOfLLHZrQb+6ZxRINS7SkPzVOXAsP14Pgfi2DuiQBn4prX/Pch01WHB31xAJoPd715bHQjbZ
nMmyRZ0h8uAh28/4dTE9nLuCdCdpX56VGqfsi5/jA63EfCyyUbNmh+uEgkNB6/gqG9w+G18nIgVX
t3A+/ktYXPI8Z6H4tq4yHQJtnj2+gYWhBIsLQQhLAmjsRndHuX3odm2ooGkXfaFN7fCIurTuHl2p
l3Nv4sFAMkLtGUlM4K5XlNnRQXcdLD7ztZncmwSztiQu3xIFLDyn28beJPlGSU8BRdYnqXrFAd4s
BQIaa1VM7FJz3MWO0zC9CilH/1koBEbn5KuZVbZEsJzwbhSUuvhmCQxhYZq6nzhefnuPX7LoP8Ay
7wXOOteHUEF5EZcFqVQ37lowZBxbFXz0xrx2ELHaNapYgipr6lkK969uaAszSUN2JJr37X+Uz4Cz
//YVSUlNWagojIZMvxUvDMx82DYdt9sumkpeFbpPvgjRXLwd3pDVLMClzrGOgpaj/sdwQDhYSA3N
dgRITevqn+a3YLXLDo4Xw8xrhjfIXtqfjKZw016fgzIqC0vYgmEmLxikQBaX+eTKdzcAOuGZ4Eoz
7J/YVN8uwc7Pe6nCbM0wuk2lGoWSk8AI6RMrgqiC0zpP8wrZncO0gcxyVi2INJJrwJZTkM/yktnZ
E1HvK+vzVlxGem9j2jl1wzksFgz2xbwPEf4sRpMD03yDWIv60qo7cEHtsz3NYlmJu2SNmuY+r4xY
WcDqfeokkRISWacYkrWx7F4iR6dD3TjkR+pbh2l6gyL7tr8GxyjcMCauHXbJw2c6xiRvM15QGAZZ
1NIPZoozf0fdY/AdmURMhB1Y1ZAtmSRiIO9PR9EoRSTGDQZUIcAso/1S+OsUX5OhTkYip7d89jwf
N6VWRTtwE0XYD6i+3307pOFsTIzLywsyL36tJ8aeB+JMMPYIF560Buj9ayYP3aQoJW+mY/TiIaKx
Iz0Uk9+ETYKhBXtqum/tMW+CPn7gPDn7g/aN/MP/Fxkfl4ZV2q/k1bQoP25CdMUweYseBHrpxsle
2oANujbXfsCJ5Bj/vFfgOfRAov0n7BG1JV/SOKHpS2YJEx+4JQwFtIprwWzVSp05zLlrTUshKuVd
sFFfqQ6Ed441QeE8Pg3m3+oqKqxqNI9OxLY+pN/kkuEdXLfJTvmIEJbZd4BT+yEOITXL6/pg7MdB
gC8RxTV6ehmPDKe2nf5dhoOio47lJ0hXwXHwcRAQb8stiTQUevwdHvQhBO/064ru4JVcxdR6Jfox
6S19NTUQW+7QX5FRFk6zCfmjjSgjzflQ8nhrlNOUMEwRXNZAiivqinUUaEzzYFpCxMCmVj/AfoyP
tnXjc8FcgSQLsHjSa4LO1bUXR0IQb9ipWyg8XznsHbFiDQzDhT2ifP+Bwy3AsxiibBnLPPvTFzmK
brQYKb8of2f/fw9pOt8y6xVnpIR1pP+B22Dz6fwBShgZsADXC2ipFhonuVNyiKAFAtTOn3HmGb1A
dZl7cwtmzgiwl3A/ytENJtaoaL8Hc+wlyUL1HRh7GVD5hELD768eoHXIvELjYbnotCM3ItTP90E5
tGJd5m9zbLWs1MeCMkD9JwxRA409pgnGknybUlm5TmQeiUOx6pvSz78X+i7B8CkVu6CX23OpDghJ
bQUnSqK+06M+Gz+7/iNeU/a45eiZ3Zd+mKnfwvvw0qnmJRuMUC6dAKaPpUmnfI12WrAZCVyIEZ5U
XrxMeb2ABxGMAEsJLk3sMvjs91LmC5efhMZB7LSlSWonzAJbIXNOQxQ2pPDsHzkioxJvEylcdqjZ
lLBhgkhQJYI9zhBG0Ujep7l8O71CwDSop8IxOQvCdV6MF/OXBJe+g39njPOJA4RgCG/sCdojlIUt
Dl1xgfHqZQStSVWMJRWPDA+eyl932R9g0AaHCLg2aFbO73f+uTnorOGiYrUdZu95AtlDqgnnlSDz
+Y1SsaQUHRAacAOKCdGw5ZpV77ufKMjcvgZd7077YJ/bk7h7+W60DLBzLgGF9G5GDrj7LiNc2PhT
AozGv2lLmKsPweHli2GgPvU5vkHtOg9x4tmw6dx2aGM0+XZfqySl1RfyJ6Ac4ac3WswOM+HSG1e1
9V9u4FNWygd+fA3FN8ZcgmW7VveV/j4uTVGq4F/FzvDY9zrLhOQJh3SI4tQP/AyljiNFkMEhhMDe
tm7AnfAY4mXOTAK35O2RvYbM/7at4GufBXg0Jv6/fgbLduKlALhYDVSBJzD7MrHJKph428YmKOb/
mlVQD6gq5Snosi8ep5EQN38YoRL8TxPEN9wof0mkjsNz16MlVynPDa+oL1X/J/xCYMwRYlxgsnUR
Ct4WAwNg15ncPbG9eZ/qCCRibtb0wvdCIzLxe5A+BGg7/ghH6ixRSLi2e8Zks1pqIMarsA5s+rlG
ElqLME/WqFS97CTCyIvcwgBTUS9oy9xsd8mnCLkv1U0HX8lcVW9ZFlF+WGWDdX61UeFL9qLY7IGv
hmLW+XS//6WS9gilLikVK0b5tXuc8A7i0DNO24yI0Gpr/E27m/bSgkAHieSLCu2o3UBnJVyzIeIN
aZfSiSVDUzFqqcLAnc/IxPowz3fpy0WuP5oMiPg1YJ6moezGy8maataygxcEUIP1SG8fUdXMUYZ1
Pt3gxwn3yiZbyv7vNEh+6UEqC9AdtSN9EcnAV0FgBaEI7/CMFv49fRIjXULAZiodSUIOjJ5K9G9C
dOybDugRfGh02O/0pqa7mQ3SrcPuROAa2LOCZ1x/MRYpshIXAMWUTNrKlXPrMejkSfxhlPUsHjuP
xS6br4SbkFsQbf+6qXy0aGN/BLUgzeAS331/Q2eLdjDQP27rff+REPaWG5WCOAkCqxbw+HHiBxti
VIodjpSdkzVSllLDfA4lwDn7qr4QvvEtP7J8FrzcMn1aeUvZqQUSyNRcwQeaW3827dFdPXAshF+6
CnN/PK++GG9GDVoMn7sN8qozX668NwS+PdqWxEni+uMBDJKHsd7wcq+S1gXu3Z9z4W5+6hwXtqnp
yLoi3apO5YItQh4U9K1Fotof5e+5G2tyzbOjMjGWXUJrK6b0vDormNhUY0FrY9MRxda7rvSo/l23
fhIS9LwUWyQgw5AgItm80XQA8UizKyKqlLHTx228FbVoi+XeN1WOFYZNC+X2fr7iLajaR0IB2Ora
QA7vDaTkzLkKKPHxR7pqZp9wOWcbKZWSzb2CXpYr3pAsJ8nmd6tAEcJHQlJc+Iwgc4rCMKy1gbCi
cImyshubJoCRfV0rjDk+/afMILdhapbwOcTFTNzd5b776mO06ZSqH/3yiJtprStwGadV1RGlpZyW
Lg3Bd1IcCF9FRtpRrsvphTbUB0nPjWty28Czpqv1EfgzcfCKVitpAfk9sjLPqLw1DkzPhrhon96y
dkE1mHu51Ya+2SVf+J+BRHamxGN8tiD680tKUhIeDpCBrKazST4fSV4xQQMPaDUUyPnp/fWn0w5D
LSsV3OEVNgGECwwSiXFWlm4jbeWkeBZTLAeUnggNQsVJQTqmF2ZFL0Mc6IHlA40hfQYYeIyGTuS0
gzuClcZ89LK21CKFXcy1qxsmil15gx7CHoOyh1jrzUNbs00dMJ4eCL6VdA7SGYMqTD/PTRYM9pwc
ALEhGHkFWtFBgfzOyf1d/xXajJUA1R/9frIS5yVESZhuq2/WrWn+IOZ5EqWP13+8TjTfUoZJpZpU
P45dNPUx7B7iVK4Bpv+TBZ6Uj5K3/2EuvNz3piwIirw9IH2ueItGTVkh5FNualsEF0oxMTYhuv0B
xPcewpy7q2Ca130QgxXPISx3dbweo2FmlxVpmG63W6Genela9sDCz2zvPRVzdS9kCNky5paApvF8
KegF7V6c7tBzCgS8+SVGQOdDKalS47ZEzAFvGl+RqHfpW2try5qVXu8C505eKp/ySBPwMGRsu7Jx
NWCpftUDnD1U+r4EzCKBsfwIL+Vv4qzke7k0Rqyd2Zb0pEmtokESz2pPKsRfyy7kTF+gAFa2LdCZ
di4OKYo7ZzB0zQvz/7alHXBYVI2tSRBxxFtBIbwGJY0ntMgnwxvOl5E4DY3wYRQBoTagsyfjKlNO
NlcJlU8AaRXu9FK+L9gqE+AkKeJ2abFMlHHP0zCJEWTYNhZ14jX+RbUkfYx5j/tPDVmtnl+Pnzo3
aSVR40GUGKsPt5lCXwD57f3i3qWYFNC1ZdpfAHVhn7LDOD+0Vw7QoI/xSdzvADHgOJNdt/eW4+ET
ZtzV/tiQBfZ122MqbZLh4c9V+SU9OzSPpSYBwMEtiF4z9qL5MTa40nLjjEuz+IYqRUhRodvK5uTC
Ynmyh5pk4DSV/jP4u/AH7q1M0AIGrUnTuonPkyR714xpapsE97S0l85x0ukQQsXlZyCh0NKAT0Gf
QPoWU40zGUH+DmriNZl6kcucwvck4bby4oxbGPs5RYgp4fFI2o/urBDJpJCnxWKdnGbOv+THo18i
dUYM94VE8wxvaP9Ski7PLr1v1YBvEh1b+DGjQQkm5MxrLVJEZvTJ8ICSvO1TEo0kxuQAVArusG5e
hSc+mn9HY0UQNBd4op7oKaYjJUrtaif8MGG7bxfyH0Ls219Ei3vwYxhGZJXKENPNM/ya+X4NH+Qb
3wgAOJMhKCnjBOL6w+oCHXrRTmE1wTVQ5yyBzKm6qEpGJNf1P6rQCMmH8ZIB5bHtKDNKvzUv2JJV
owvjVPT8F50aLc/gjE7JZByG90HziaeiDGNAWJ1D+MYF7lleLUpgb0HRZ79UkuTNW1w5hvDCN4KU
NooIxv6Fy49TdzHMekIjP4Qc3aPdpNjLqYG/J3FjXRLXMeMM2WqOTqauETHhVNcZjPm+idYmqKcu
5cGqOaTmp4q4jhCSQLhtAcQIo6pi7pYdPjLJ5cF8T19WK3a9XnNTpw8cOlRiDEk72waCqigr1TrJ
XxEZVwXy8bDp3CAKi07IhVs/sFjMMqFNXNqoxfxPsFtKKQMWn+2kfqc4HhZmGSmJMyBsG8EX0mCi
9+U0ynf7b/1fKI7jtz6TjwRs8c1bRvW2CE0eWwGaXsfOThW6tx5kgjt0OcTTxPtqOWP+HHQyox7d
6lp9FqeeNLxUKsji/sOvYtx5lF1lSLO/HHIIzOqLGNHYkCZ/RkCFj0rksGc+Fk0WR3u22tIERsll
fbyZmOsINDtl542PpIHHAdJfiaJtRwciYjjC0AHjWxSOkokBN538DUELq4ipF1Upx+MJW8Mg2Iy4
JnuHhcyET+quga28WTZL+sM71rfSNeHsMwDwC/Qrxeov6DDOCDPfuDQl37VtDTRzyZszkQ4Rld5n
YllMcLyabHe99MrU06rmVWnehCHbdzTagwQ8Vk8QcVGUzQUvBKnZRSjRWRSEbc1oUyZtuQ1HfwSs
csajuL/5MyKRwPLa/vkufu5KPyTkSFkrMAEhbTGUX6W8yE2YQBNUc8mMa8ADQalHU89C8Fw8xuqU
cqn7ZQhImjK+GskO1kFFB9QJv2FMj5s8DDzJ2sygZjCxRA0Oe4z6XvWkIwdREN8/ob9FCetZ+pf3
rfzbKA7DmpzQtUEemqQoczfSyzWaEDsYd1FJz/YHEhMdN7iGqJptmuuRKdpe6+3rXXR1FYNMyt69
J1PMo2h+V9S15Y7VWFdy9gNm8X21/50llK2DgJO0vw2pm+51Q+IOTAiq7QLMeF9U51vJVQVWfN8H
xV8Jo8f2ToytWAAshoz1u5ZbScfNcx1SARglkkjV3TdYxHke0iGCrE/bZdp9mP80IQHg+mOv1LRq
zGcc+p5NV3rMvZg0FzZ1yJPd0kUL5R9GCo9y0ePZdr7EiHh3OqlDDOB9oOIrBGj/Kr0bMD0VfmyU
H/Id5CAqzwsNQar1gsrA+wkUc+NKJbdBQruP8CIJCQmfz0DcdY6IZnijf8u5OlzGV9/dK24lfF3H
NPvxMTNKzIGjATLDDdRQgY4fgswS40m0wnAYd+pHFYIezkf5PV8K8peSfgOov8+mHjIHW7ZSRMy6
WI1f97N9JO1Sf2E18YVM0d9rYU4+hYvsAQzb0BpNdESW3diruOHvZtLlukPMaXYcKI1Xwa0cgjM1
XxEBGZiHpdBvKRsEIQB8A3arhO9KFVfo7JH5MCwBYSU8hM0KgVsel0pxFhneZgOlDK9HCeWPPI2/
50va9BE8Mrrvy3ZlcNXpC2n0vnsT7x5FVYdIyJ+Lkh4ijv1/Y0M4Nw2Vn0OF133Ka9JFjwoC4LeL
iYasVAN5nCx2Co8CLbEn3kpfPJFLYrmcHZc6PXianGSZFgYYSIZQ+dwfRN6U56wvsM05LHPdCj1U
fgwBmwcacQrknIoNyrA9C/FpmK70PvrEmFrMsmpsOi4TnqGzIWT09XUHW/1i7ev/fjKRttE3H0Mn
A6Kysd7HOOXkNL4bnBHM93AwOCvYJ8yI6U6Z/kiFu6FJ/fsRBiQ8CPmJgLfz9Z6lcPQoxbpXwr11
7ZM39gy7FGbZxgnbvDwcbffREIQo0AoI4fqNSzqfr6N0sE9X67knpVuf2KrWXUkal24HENrkdhCU
xdwNbHfh/0LcVw7TFjSKdJIO8UPzsn9I19j6YBBBjzmPB6qlvoDidPyPXWtnDRRHvRyLSwgaC8cQ
hZHy//I6hyTwx1cfaTRvwY5wKEf6Oi/G4ZNazTOcB/k4wrr5/PAW3GXZyBGulnRjnQQ0tWrFD0EV
vcHIW03HoU6f3LlGBYlU/0XcuvqcyuWd3S6suprWMjacb1sS2L3h+v1fJi4OQCGZO05H27hfZomp
Qgjr9ZAw93ZljVWoWVNN9xcOTD0XnXZDRiQyzDJDYAX2m1v+UaNNZ1eLtXCPtVLXjFFPvCb2sfoI
OIakNqiEBQGH/rFBG0wjd6gb6wn368dzI+brxnqgUamqQXHLff7RK/wRluWfgCZrFilE9Y6mB59d
BtcH986YZ2P5jWjXtqLRa5A2i7JusEBlXgyBvqJ4tfo4A6hsECNUMRLL1Bq8yZOyN3vxfAp0mNDZ
VTTI0QxvmIcZUaWMTYo4J2iWe7nLDf7pMl4YLo05gd+3+T3QeNVekh4v69bQoHM8P+oaQDbYaQK2
BnZJns6LWEr0DKtfu9FN83vjmmbrKOPgare0KDJYD6iVlpME+5RHZTF02h1maRRc13WyG1CyQ//6
4AIgzc8QzzojklULnOBtHe3Xv00vZejHD5y95jUlQ9bvihsviDe/Pg5BRGmEuF0+L3O+fZ7RChSd
hRdcXTBlXrR4tWrZyYNLQQeluOIZ28JupAVIt2W0b/dO0NeOBrD2qt3E2yyafmqyciPdk47UOamC
KBmb/VV3Arcw+TGTXxWhtDEUW0suuMDpMUzNY/fMSO0V8SAWT9rxJ7jALbgzUgI6gUs6/0Hs3Ut1
vDkfw6mNUl6/r//NaPHfV33TApo7sOysE9GSMfsVoxJyKg8SJdH+0kgfvwNtLrcqYBTazTp0sGcB
Xf2YHhjiPdkrQJZePlOJW5TOulo2x+y8fMAiARRVoJ+oaUUhRdLY3Zvntu4rcXhLVAhAs92CNe80
qx/7FDwdOq8lTHlKiYa7v0p1tcp8Mm9b3CYl9yzPNM7f3cjwrgCfpBvAvDByHgTTEQeoQHgqgXNR
RMi6dKcn9EZuouYY1eQdCnEuLijG5HQfqC3VHDL+FX6mgdoHV9uwvUf4fGrRPEyLf8W2U6L7pwFs
QwAzncpG33EnAgVillhVvpf71QXwXyaE674U8SSpyv0eYOWgN3zE9IpOYyV9THR7cUzL8yxGssul
ycw5aEzoqrkS2Cq2ZQ6+/PTGp6uB2YAA0y62wYZqIIphZWBbMxA1brjvduwedjNjCUp4Cd2c2b8d
4etq4APVMUGBLeM5pukXrhzKLFQU33vOn2BSRlFjxYJvOn0nX+9pcySXEbZoMekEOFwkONC9v9U0
0GvFidF9RAjew2P9NFEDy/h2f/2xUlzocK5fmom5FpSTHZPPsPW2h6oqBZJfs+ZwxFGhUPKECwvx
Y8NGvMHrskwfX69w8UWw72kbvXlVggYbSYL4bBsqjXJ5QfMWpsRC0fVCVi4f3HmRxu1BerY0jQxi
PSH1UIDPpw4dNaQD/9DmU3CPgfW/9odgW2h360d8lIvxZcPay2Yl7vO9EjjITYtn7C6PB/Ra0C98
aDi1b+48AP4mfzonQn4e+SFMYNKJFcFIbg4UUM6Sh3X55RFHsRtrSPPIPCQODp/DlzR3BFg9TX7P
3J0lMZvsdihOWGrXsVoP/k5fAhcbPlth6Bo2za1gu21bvxHoUIamYEHOjq0irdGX/aW+zdM8D132
hGkqFVeD4hqXMFEm0N1s5/2KNPbvbNBbR/KSfVNRwGE7VV3EPlgfy8521+ZhtonRcI3bYeaj4tUp
wg7VHBVeDMRzfTuKWg8CAbT6rvClHvIVfSb2Dc5x/Tdddl3lXjBRIR/qE8weK3ImuiU5hGmunwl5
I0skxN9Jdn8xNwUft2J/O9e5ICci9pk2VX8kkRQKHlXQSIgYMuT8aRhh4aqQv+sE+/+1Xwsh6Lhg
Cmtcc83fAylKkujAmE8OH9WVSr+nDFKNrEgRB+kghwxR+pL6U4BQ9iZtbEO0Tduo0z+U+tnGNQ/w
6WUz+a2FCJMmNXGtzqbP/9Xol6I+4Tq/KMuVR5EwK1IL6gsynEyFYRk1tCn38zAIOfoBV5kzoZW4
Yf2CuP76P3QzdncPX7UrkuZRfuqA4Gj19aEDJUPL289ZyQYyomyMsQ08jIvGFFTUUaYcRSEvANwL
U8iFh/9tm6KWfVwJ6dM6J+A2EGJ+AjrQ8Imj5DZjOd2p+oxb8DUoMhWnS8wUgu5pfq9AqIiMvppK
un6ZM9EYMwQI1rTXVCdoIGhBAdvlzmd6zP22xFudpXufO1m9Uy7VD1k/+XX8ip6NARR/UJ4SRHYA
UNTVvdaNb/Ggr+G+hZPA4VYEHDuzu7TOr5x49TYP/Q7tmGbW/EwMxjpVUr+x4et8uoGk1xPSMCwn
+5CIJNiJKJ0L48H3354YTSKYSTbJPr/sALOLrjhh5Xci1SIf9clx3HIxG5+iKJ/AruSeRPeKYcvR
sASjxzzXYGqa7hsYq+e0qK1PJ9OEzNfsNdqd6lIijH1kxgiJuISoCn/Vplh12rBkndPyZ86XCb1N
xzD26/XxBijm813kYphboIfyQwHFJiKNPkTv73kaJ6I2y7rxwBgx/RS4XxRdcNsgEpOnr4xsy2++
uRL4ooS3tUMjiaPdxBh/v2mU1DlEoyulRHtt9l99FTTThuYeAou0KvOmby5odjU9xOhSSnuRG3MW
QZLuD3zQnlRkXst/d9Woq4qf5v9VlDXP0YQeCW41FyMhi/7ziAySAULKMelvI+FNI43QHR+XhFLO
9/SmzKDMXjGqGwnYkny07yQSCOrAjiNhT9elgutpqVYs9ifDJuuLIgvSFICeRTG/mjf6lUX+a9+6
dESdosK9QzA2b+3b2Pn5t2JgIAzGoiLjpLPbsRpiUaU1OlzvDiz1stRXvcgAxO6uuosnnpIr6H+k
tA/bsJZWDCf63kFb9YDEt96hzGvvYDjmESXl9Zuj5z1kP6ORVB4lRI7vvgsQp6nUZeTMWZlLz5Mq
M0P6XQIQPbtvZ6eM3rtXJJedfhTGwfOJu/JA+VrF1n0W+wvRVmJgnlF7GAZz+SPhNTwGFYlz10u7
M+hZ3OBKyRxMS5Fs7+iLYx+7+Ou4h29UIhMZgKir6T9Kuq8GO2VTPJIZ22v8H+e/XliQ1lKSrTEz
GULN8cfv1oZACZCpYor06uKZf0N7gpYZw2NM7S2qruvmxp/cVkbembJNCfTo4IBqC/8pay+vlx3e
q/sHyqgY/0Ht5cVOqU6kimdd2wENq87MN8bduSIEVpOzwKexMnSAG5kw5hgADLWeuxT4ZX9zwU4d
LvXmEApnPv/3FEF7yHtKiDrzI9n9SMOqJTf7z/z9PyZfBPPFi7bqtpM/nGRjcRIFQsyxnTYE5jVJ
EDSw+dYHrRotvlBOyVb18JyIVbtvp53zCDDrFNJGwVX92Knn2f8fULWe9nDEUidj2Xd6NKUknfmo
nT6aCxd76i7+yhZShl3yTV+soB4oLaurJnJNQxwz1vFSI4gOBrjsPi0wZ9mMvsG357QcZrou3o4Z
QE+q6GWGgHNWt20hygtV8+2kF1clgkIS3nlWyCFfV7KSujiGq92JlEoB28Zn/EeoW++RkWncJdqq
9hLzo1g8MdsjB0JkVhFo/CFQ5FILz2TXJVikN4LRnDqb7vxi9tKM8IU++pgwVWrSV4htHFQOeNuh
91dhXV/fwP0x9k+NgKC/kJtzcMdsUPrsysC5VQPaQ7QAaKXibboRNcUyvSovu8OAzrC5x0L4BOXM
rWMydWlfR+7p0AKWixWrm+BF08oSkadTk8XH81jWvb3tpp8QJzQsl1wpvN7tqayMeCxifUZhqA+3
zQBDugW2I0U2QCVZlhrU2K8Xj6W9IuVAp54VL4dFmcTVNqN9AXcvibeOrVLe835w0eeohQGjXQHJ
ppqGTiRQDkpXbQFeR/mwoTf9uY+IHYSRYq2+U+GWJkgBFQlFXvqpg3xYpoSo5UTwu7qewcmfPO3z
cdRVIdzLQqrXq007taYn37Ooc3vYdFAE2j2Ml9NgfNejqC7id0iKEDsaICA7gB/8C9fu7gSxV/iR
p2ZshsSv29Woojq/xm5BEJlOHg8gjwbe8xXNhAXoJk1sW9ml33hxCevqyhECX+aRVQeTjl1JIt5o
8aCj6BGylmd8KQcPcdosB7O4ptWFv4Z9FymiPViQaUqIOQgb1fjDrcmWswKRTFmOIGpmARB4kIFS
AzLpIp7FJhvLig+e0WdcVgn7LFB0YowlF2V4fn6aam3P+6FLvnsqP6AnXWYinXkqgPgDmmyBNlUY
nEzLM4o+I5vCq1WzbHU7XVRaLW7m/UsRNcDmeLNHJ3vwZLEFUJSvDJ2vAAoltK2e/5IHjv1iCT1H
nG64zcTP1GCWYi+foeG6cY2620zOKrpjIJxrzdlY2DakKYOb2ngUXhHav3TkfTo4R2QS3dOrLyQX
UJrmdSaPOU+7ewlBYwX4afklxVRVLe4tMr1QC4mT73stAkINv0liegcCBTSYUhhrFNo7qROI9qJe
4Q8tQrdz/rM0XssUOmXx+pWOYplZblo/FboMxupbDX4u5VOryCL0RtsWR77PYq/e23jzoV+4Za8v
rIXtCRVxS03bCzmV0J44fgE6Ckp093YN/QZ6xjm4ZXSIQ719rmSjEu511U2U857xtqGFJDRM/olB
oQ/VTIp90BjBmxW9X8O9/v1o1dfLXnjQ29VMQr9FwhIyiXjfutvB9aJNUByvpK9x0Tkr5OsNnQeo
75haiWOHxnM/cOZ+W15DUspBp2oxSh2hMH+zPGiuMR4ynWCBjzH03T9AUBOU8m4DYoFH5dniBumW
1O846F9713et6IhDPukDBvVXkKs/zG65og2ntF/QJziE8vDzhtbzF/oAyo6bPEzjD0YBofhR+CBm
CPt8H4h3Aetx/IAQgnn+Q3/y6DTrXsNBTFqI1V0OsiOYcopNgNPeNSC9EYKgdWqEomaKJb20Iuge
qLXj+4WilNASEvnYigrQeswqBEUICy35libh+hyv1bD92Gk6lxjOF40eTgePRmqQG7B8PU6MLHQY
tj67FY6cC5k/QYXyKOXnB6UHBAtDRidGk9frCog5XMHfCvkNRkGoXudQZFqJFa3oq4E9lNj0PO6l
C8Ft1jNlxI8/cSrK1S9r8o2b8KqGLsnUnPTVQ1okZy8AGIZuJsdNXtKM3UMCluMue0WPrcG3buWW
X+UO29I9T7Qx1Rk0wQ34HW5UYbNEg8dpXLNSHlMv/fwjabmNEuP7fhsFRcXwya0gHHxgq5SE1xm1
KwiwnXemX53F4m+vM4coao0buKscvZ3Argi9B/duQ4mfPPYxxm53rWgIXZ6tk7NZESV0eU7Xbvtz
lJvPyUO8A79CDRiVqONmUOmpaO23BdDuY/MaTBbwkAXtLoDyDgYqApYTew0fum+V9Yc+KMymu0yV
o7KiH7yxQ4vKYmRYQOqizBB5c5IWi3Llnj8oPw2OD/FfhUQp1KxsWgYHEucP6L1Lp2jNurX1Busy
8aUWPkbS8aBGwS3EkuyDDsieeDY12dq0XD6NR7U1cymIWDblIEt9ujtLZFLfLrTJzVDWxQq1jOcR
5NcYv6RfIhKn+5iuT2+TppNX3FjxsaDQbVYX6LM2mDlLkEApD70scPWgjKbwLqbK21QRse32tGTM
dTWEeIhxE/OpisOV4yRZoyEEMc440AciZrFy1yvOURNbznOQonFDke41Aiqiyfs7xbBRHcjBjN7z
We1s08lEcFodNG/MoKhNztIZ64PmEdz+dFHtIceyL2Y97X+uhsuLB7u9QiIrQaCgOuQ/vneF2XgW
KhMfAKoNDlTVFTBc7aRwbJuuZdTLwcpZXssQwDX0yf/Pq2lyRobbaZvIei14nxvM/0Yh+vt/ECS1
tR0TJ2VqZgAx98tgqlVUMe4RT8gtwcii7QKplBEqk9c1ruY9BIPSBFwBnpupj49PsJjn5O+yCxmB
xkuebGhSZivrqLzThzG3kD6dJZmWvuTgpM01IyRGyhZkGdFHnnMonehqX6ak/G6KNSwKLeHdqsBA
w172Y/mO6rF+smozMRZPakJhQCaiqtaYw5SqyWKUedfuJECF1Y8d836jGASZw3U1ebkIezBi4S0K
ItotZlKhUb/NjnGo5YKohcsMguB8cnP1GFxs69Zgo9c8tbS1W7uQvRibRR4sydMvImiaKW+qsuRu
awOblz8nUx9w+q28H96fvyNfNKtjEZ89X0IMxGICPUsxerON5Sp4kOxkBB60DCAESOn93nbmpzSu
qComBliEvDd9KpgDmK877O5Ml9TASzX3wPnn7ay3BvVj23bgkXa2h+kfMZ1ritetBe7jm6727VpL
R2VDUXGgGFKf7wAKWrEVnjlD+IRwFpDP0TcpI2MTBZ3JcbaI+sgSUCXa7l8bc71nmxneOvGZXqnI
exjoGIZFLiZ2b4St0/+yWf/4BTtSjv1Froeee/ErDvPpeEkOScZRaqsEbpswKGmGrH+deY49DE6B
RnYcdP1TMnLuxR5r6roavhFbzrlpvPIjwLyruTggyVx281oO2m7eMmsMe6mKsOFjqXYf5i+c1E+e
zkEP8PO+X1j9/ZgN9NgDhSLFB/NcPKAOPwRrVzupgAfoP2UQaBi2KRFjNznpe5IKJ9xtAeobHaDM
Mnoz6zul/i6XakSoPKFujbKU8qtyCUAknzEAHpSJZi5rfmKBZ4wJnJi6VrlvGDQyNT01Qn7Apwt2
S9ZjEKh6AjS3yAUJr/34bFAT6cAaUT3jyBO5DOGbVNU0APAfrp2mGe/8Hu9qQTNITcac15xevqSH
VYFzDcxa/k7JQi8/JwhVRqrmw7p+gp+Ul6m+x56cPiBqWS7leYgQ07c1iY6FqybSWe8d61rcy7o9
1LET9sUoRyTOrUZJimUXwE37tT5nvziicQcH7AtuD66pxjpgo0XEoooWWrdMYWjkIrIx5U8hKWN6
x9Mxl+tK94l3REcva3+Cx3cxcjUm+J068dSob/vKvxZQMcsWWrbjFsoa2ySquQWHFAUKiS4Vput7
wdxnAyCO08Cch6gbQgRx8GAKijkeGpdROGeiyVz7iwN32jwT0MFFuuVmDBVsfF839mS68vGbOH/F
B9DrySMQTznOdkntmPCvEAQ8KcufQisMSPJD4iTiDy8o9Y43VBGYEzCigPwpR3HrCT2kqocpyBkK
tn8+kz4HBXLRsV8P13X0G2FpaigWJC7M0jgILuFOTNBUGnUfGITjSU2XJL7eNZ/ltNtEDOZvre6L
yhoFAzCilqajCeb4LIBy/B4t1sa79E9hkpRJl4Q0xRr/stk/5ZIyqXJ1v5zFbmxL2A89ZrSaun26
/iGqmMfxU9/r8hI9LcY2l2exLAB/Ng9G8PHzQortO5l+2v5KttTm5fCGX5K0qUdKW19qDIxwtK+z
hBJ7vqB2iBeEQv8qT47NEYR3zkfdvWPVa0bCIQ6X3M261ZxZWSMxTMTCzn9CJLG+nXF9jAGKN6U9
XEsTwNKhdkZ/jMcIGfigITfR0h03sn1c9ylWuaenwHM7ay9xMxRt9pMshi5bz7WLleEEhu9zjAUQ
jSdvlY3SSiu9VNRX/pP0KpJ+mvkyxkEhgupE1YVTbokDbnf/zirby7mHsD3mRMCDthptcMAkJeG3
Ye5zXyRvusoExbhkalgBlxeHzbUFI82FmyH0zTWSccUVwHaGskRtYkVcTTLZLEMgBRfL/bT+Gm1U
jasOeZWQv/C2WCXEJRi+UXZsH8kISi3goi/9URuOe4+citUDmidOWfdC+MMbVSsuasimiH0O54It
dLcceKyPefD3j2o1eppoDfzbk76DuABUauRFAvd8HHvCP+/5rH2LXhFK6kGqArJ5dVTklVbVS9XD
w4RC3SxKT8EVHULR06EMMm2eAylYjlZr8pURdxhF4op8GgmWrBbpZSXtd8ylOcr9gGQYANRqsQAj
zyHghVBg3SfJUGPFr8r4SSj/jcWx7kwO9mfnevRx/mxBIqz0umzxI/CViDk2771WMRb/1FBmjGNM
z4F8ILqwp8q2evd3ncF+CtK+WeXw5mPTxcfUjJkBqfAmg4Mjdw9RpFWp5JB1oYusjKFJPDKvilXv
S7Az6lkgBRyxFAhMXpC+MZUAInPODJHm9NoxsO1wli+OZG5WBn6zCXc9f1sZDRrY1d0EpmC9chtF
9vEr77hIA/4xs1VYkLjrRj84a0xgb8f4ObgODscTE++1ar/R09Cg/ZPGabI1ESwwTnR5JBbR4J9J
b3RyIii2RZcisNhK6VffsJMk22h/PWv8Km8gvX7gBraOpki+ZEuCCVD+0ykZ+304pQ8dpSV+T06d
5T9J14CSKrUNvKNFG67NErGDZQBG4jVpLwD6BQlsjDLW029inlwBgGqI1vNxGhmnbGPUtU9ZGImk
+PYY/8yxWEH5rAKvB/aVQaP8b2BC1y3eTIvg4fjA3xkI4wMtThmnYXCjLgzr81Ir21RGxF0YexXB
lmwlwkGEx1Oh4La/eDmLoryJWxsA5WpK5H0nAezP0kzwMuT1J9utaypZFILC9j5HqYfsayEj2YnX
3pmsl7qOM6Pg/d1dqBFJbtcF5oSZUNn4pIwsFcGHPl1TEZmjGbd3B5VeFh7lHd8ArEBSFKZH0iJJ
zEOWeB+PJlybLofdy3zZBqFjCTnxoQkMkrnYH5K3RUGjMMdpXNOswCEugaHEATGsLrtohABtvLUo
EFB0noU9gOxU7l/NFM3mhTMYs66yMasHgTNfyw2v0LfGbuOPMmIPEhkwrUXJy2bn5rEy2JosL6vl
YFsApaXMruVD2yYWJYPvUBNLpAiApyx/J8vcJ8pTQZBrNkSJ2M5vhaFE2FKhqmPDtj5dcYZpVMib
Fnbbtvu8EeFgQ4T6p7SGp8sYrbU1otfuM1CaDvErMKiNCI3vONodY36vLur/LfORibhD5LON9RZZ
x2PASI+WurnU9Fc9f07jB2luR7VSY5lP1cuKh0YjU7rMs/iR42mCZKYcAvDeZmFRhjAYTEeW+QgU
jln0z8RqyFRgvpZtR9C1isajVTUpx/pE5uG88/W0ZLaSwN2+1fqrPy5r20dMYCXInxMFKi1RsW+j
YtOMb/8DRkb8Q2SuVMldTokHM763rIlf6uZ/QMZZZZLd+OPTzzSxKk4raQV8NVDXTitMWERd2uxN
rF+RaRBIZbkiEilzgBAds2IC2XfQavlkgVIaWJEIRQtID4QKSEDUmCn54jJTTZ+/XMHEKXzCiDcJ
+qCw8F/iutzyWwJ1KF/zNTu73bLCFAn/PIAUhCMh3f0QTIoLynrtMBP+OtLFpECgM4nweS5fmiO3
vu1oysYeB2Da770kEbnX2YTggVrth81HAZYIYnZcmZD2aZCy7/mzKnu2L9hD9wA+pYfJw+bE18pP
6x6b+SYwaU4egA1/ltS1rqi1FI5nTc91X+yEiQIl9+oVRNMsI3jseUsV3w9Xgb7412WOJyi+njyc
+zAgZHJmN8hfNCkt09v0yopnFh2ex2TeNlJUrSs3iO7KMuTjMovfRJ6mXCGfkpvcekl9kmsjQZTB
YA8+397qge7fyJQMOI1+Kz2/5JvLmMRp+A0iRdRnXkwzP2NFvQSrMyRFrzxT4NWUUcrG581Cxai1
BJzshJwBk8DYUOreMqZB+qVOLwP45tUpSnH5MIxiZeKm8hnMRZaYrf8nJ98RsPhLEgFnCy6PCfFL
3XOj94Ok2ycV/4HO47CiBK81OPhOl2+XaFimUkb9Z0LRgNGE/BRoDfkW3PJaxOnknuEWsAyOj+d5
7HScidFG4x3TN+qTxEELlR01MR+J/mv0xg0+loNfJ2/jKZHVLy6drmJWTYlKn0DoMd3f6FrxF3HV
brY9TN9+itMnJWMmuB6WD1je+m50vkNBzqbu7jqGDTplUFQkA0kv5bOjO0hiXlp+Y+8u1P2AmxvO
jvaa8z3SLKj7pQYkfH7rrDPcH2/Ko8sC3r/0RiqAYqT3ZwLes6cBVajR8Lz9fJqWLPe8sMDiKwM/
kDlZD8pSPw/z2uWabcG/FjIw739zx87l6NbbVz5reabGEE3h+agZ63x+zf/OOUo96E4fV2S04N0l
xM9bnKLz5VaeZtT6wQFjuo9+RFooS5RChi5ZIFQfE8V9xsjhLNuGMTxeWFWQYcP1Glfwg7Ma4oxr
naf4+VIKDTmf1wO503FnPPriJvgk9iP36/MWthuhaybK6JrNB85eyxjcEB0SM9GnR/OFm+ZS8uDM
Ff4tob6VyUFdaaSNvz+lxbiqJYK9TRtJm44WSDQw0EdLGaejZCaV6hMZgyg4LlRskNpxW1FJ4CoR
4bCxTNlWSBbrnKeS+7DfzBNKgJyEMpJHeyjBJDChifOX024EUDy9oBka1RdVt/Tmb8apPaLQf2ap
NXiDHNND6AadBtLes2/KKFrxNPkuRSJvewDihSAP/SEhJTtTYXAJ3c9IoFOKYrp50XfDeyWbBS52
/cKhFlYJmO90IjpMIFs8YxFlRMj3oEnDgOodhOWt9ZD/blQz/kcIwUwViyV5q3ptSa3HAtCK97sN
G8py8pAdjYPZVI3XW3lf7S/jwN6dXlO9xlLXn6YCDF8TT/xl/KL25GH2YpsjMe0ksFMPxjci58Tt
pomyiLrKVTsZMDtVI7mWheZojAC8LjDOlTNqtPzkix9qnnGae3uADV3/oZbQ7y+9x6eP/OhiYYto
dnZ7l4Yrb2Gc3+4wtwqF1bBB0g9oQQ+o9BZSRCskw1oXIugPISjDg5V/ymjaaps7etUUNZzfALHY
8gBy+VTs8UyvEKeYFCKVtDWhLs4qXK8QAR0VABFEqv0HEq8eMWFEeLW996TqlmYfSuCWGxYErC1F
3NO0hRkHBgk/lQ5UrVRS/AosxfmaAjlcZWtdOf3lP+tTZ6WxlljGTaPeMpoNZgnp0fxsfi9DaUkl
JzAdOQkwQcd+W18XYDNwcfREyFjo+bbbyviT4uG4FVoBMI/x77+HBRI0yzz+mYzyr8VjC1h4eMxU
9onlLkyi4sj9Rkc1rDLyJvaRFb/tUbG4q33xUikhB0z6Lw+juktAiGDbxaTkimH1hSIEfEQVK8Uy
UeelktreYIL+dSTTU718YzPcwTKxWDRYLuZvbgiHYnC9W0eeJs1QK8ZRTt8pD0vs20HwGKB8Etdn
5v0LRVsSm9FjBdQ5GkW9ZR8vD67/5KngBNOdgt0K7vjMGj880zkkeb5GTFbSh4FX+6L0vrEVMjPS
AB12oaApbXIvAX7Yu6TcuBi/E3ucMLMBOKiPWwjqz05nHCemFFP18GNlszMMr13RvELdLIqshCD3
M9JdCS4rd9vcIJuvsXddSOjNZ9OrdGtwa5XQ8Ci6wLlSPjgvlQQh6MnDS8sW6JYhLKbbNmfEljOX
4w8wQmnFbLD+2pXRMCsrL4vGPvuZe4YUhppgaSQYFHdL0niihzFDeOT5KYM5j7aguNqWKngD33zO
Dt9lZ2reNwkzzLAqTgwzU35ie9unEYbZq7TH+8Zmwkk/K6jxkJF8L4H5Ge6I3xlylykMovbe4j8H
ejas3mOL2lW0F0CYKNNQgx7r/g/CAV/NgI3M4J8xqs57feAs5mqnS07x3SfDONb+2hut+nZ5xYLf
hkvR4CqxdwksHLMZcA4fHGEa5/odA0ENIrZrHheTFeoRZtocDtlqgpbTxZIJ0lTNg/Jot3RqfTvx
Ky/26NKTHs3y19Vfb9IpN9EyiyVrK9F0rIZylm6FjkL8qDOtl+DWcX6D1tQ5l/WWK8PY8xl7cUEK
aBdCnqbL+o5KiZ2AJBtav6Kjfyii417TNReUV2rQGx1hoJ1Dk9LPua5RlAyndoOs9c2+PSNsSwJY
18GYDDtjdcRzUh5yXkulT5nbwFn3j1Y0sPwjeg2mKJLGNl6mDLb9LUqfrmZG6GJuYP8GVZGPFFgb
OudnnXyQNJVcDqGTeODGcUPRjXFGlYItNOCApchAwxT14AaIjSxOJCHzT7D4AA8xFhJriI7E7Q45
loVM1c+NC/py6zguUuOKQu9JSNAKLFo23go7vUUstOKrHV1fYPu3qauQUvd64w0wC7slWtd+/8iS
MOcDEKI7uCV0KACA7yfrBAbMjSVraeFrMGWwCdGjpXsS5X4oCYE1ngvy6Rhgs4WMtnUNnno4YywH
31esgE09m+CdkV8NCGA5O3IHQq2N9CQMTKdYedHsURZOT33oDUDwj8U7p2aB/LGyNXFFG23xHPRl
uV2VkV3ZV9Yws12s6eYVAatbB9v3SLuCe07nvsVeO2am+zfiL7Mtu4HvnBMp3Co7JqQX+yUZjytp
p/TjmNG1RE4T8DR863pkHh/vQ25+22R3tXv/bVv3G/A34LRrGq7ORlUC9aF7ubt1ojFu7yc1/bM+
evIqvupdO+g4XmLjcnyIrqhuft5H7ECLE7XbAkQM7ifXYlMnp+k7HaypSAjFto0Mi9sIc1EsRDBM
dSb7vlHqYz2oM/fmeDQBgB6uWLZSdQuSe31XTtMtPqeWtmsfX5V7ufPWIzBJLSw645h+MrxHuX03
JCsjjnOYVb1Advwfn0rTROVaNgHVcobjTMBqadVsQnaKR7VmFyReJXU7HcN2K3Ks7e0vyen2psR/
PTaq26w5RTjxbVpkhAVGFHQsHiK8LkgI+UIg2m6iYyaUYRjrP/6wM/Obx0PWaZnQzwIAMbVQcWZO
y3e+3qOl2mRz955aQN5bZy8FNFXSUFaJGtmtd+FylFsqlpVwmu7mXU1RFrkCbIBKJHN5CnIEeCHA
V4ndccveKMD66KKFTxOqDEqb3HD3HfDaEIDsd1HaQAm/wJfxlCvw1MYizXZmbWnzy+w1Mkd7Qf4z
b5S3bd3ikJjlxeZw4acSRA+QqyVQAptsSvUCrAK4RszapjrspJPiL9FGveHKQmnEQugXIS4hCUAd
hbziZTImE7cg2dB4uCyOygAq2oUoUzcc1EAEqnfDA8uOSkG2tYXZmMp0hRArFJ0XlCku0BQiFnxu
AH83EkGdwb0CC9Y9vDGrVd9TXB4Oi2sdK3MGrsRxJf6WKwkYSCZDnmLh/bV2UZ8tXAX+JUKTSUzQ
IBgGQmP8KwmvvS+ZTSSluU7icouFGIENuyQoyl82R8TF7C3Dg0KDOxj7CXMCtzvC5TrBPYfxi5zn
TnosZngFybze7I21VitwCEIo5vD6SLWwIpFxprP7cPI3sKmf0q2RhdoUTTbEsSLBxVr65cdbDI2P
dmC3JhpkZzN7dKfMlFpJ/SJ6rJp8yJBfilMQ9AuxW95zAzWnVk8YBExpl+PxIvWQyqg6ABH20SYg
Y0XBBYaDQ3JPeAn1tQHAK6HFULzgXZRDqVbevACEASHtrL/heuKeVXn/oZzOHhlcdcKjh47P3xtM
7MyVJKpTmvuRUX49+S+oIJdzJtXQCNjQvrEzI0KavYwQB8dAqgQSJk1dH8wv+niWJwpbTRP7z3VE
je2Aahuu/5KcHVGB8jg9KGnlNv7KeNw7Io4pYJdG7xVxkz0WdECHT5CZjz6WLoh9U5TAcviyhc+t
LnH37C+d7UCzl3+ZSeMQUqjPonl/GqpZqhESGPCPIwkHovAKFUD4yYdeOXVw5ZhSjOnW2TAjhoUe
oUM4cW4BrQYVw6nrlue3E8t6yvShyLI0FYmoFjACZc6jc8KGad8l8jhC9qYXnl6GBZbTiRV9E+gc
iuCTzEznfhdLK2sQt5Z2S1xNd5/O8t+9+9nmCqexJW/JGsSPSQ7co0/wCJ5O6Z5xmJReNlp2T0X+
rgJnBgixQ8gRPSHVh4+nbVfCQD6rXfXUNl9QBzEHqMBIXdTcgWL439Jz8Tug3K08w7Asy1yj1xtM
+o3Jecjdq653rNtOVF/B2GBG8owHp7lL9OSeBmHxo9HMr1+gwNSSOjrluj1RKUbT+T6gEh7Ex6pO
Sap8LQ4RzPOPgWpdiytyky47usmYt9C+iksd6MFbTqRh9b0YK/nNkF9nsirUp3hVAk+Oh2Iiu4oS
aDuCEJazAbZNtvtX+ozlCFSVz5Lu9IeEv6VdtpDIQSVqXg2BoWR2W8QUxrH56rAcG9TJ1BpWfqOw
53gA30UFaoKHfwUSMFOVqrhky9tWmB0/u+TGqKv2J6fe/LCicZN3QCGhjpIuHncpza6wrXngVscB
VzmwBKK7Z4O1fvD6+uyzO9+INIszt6HwpCWIjvtZMU9pqaFFUzdO/9ti98jKmWO/29UWyRP8geSS
yn8nSpAjOIQyqJAse81kE96RC6c1fZBP+OCGLdQBhF6yMhEnUP3rO+irqaXncHzia5eg5htJCUQI
LeZaw3Yn8bnwwYZ0JlmYwUFhH0aA7vk4gi0gQ06fK55uC+IQSaMvvlXuIPDeQISuwo7kZgexNhH7
G71qGiMS+xvwwpGdzhE06l/wPnEvwUwljEv2MopFKRal8jeAGBJTGo2Sp23uMl3+TS844BVgehgi
9KwJQP00vyKfRGruvcRSP/QD+1zyxElK8HPA0ECYffNBFOQZs8Vtx5wOBT46WNf7MYFMZvu5iT3/
MvRZNpU33UihTOqaaY1osI7VDGyEuHJGNUkE1E9Qo/4hB9Hm2SOkWOI4znU4l4tZ/bzmNawjZ20X
pcKJOYNXyah3HfowUExUkwqtNZWw1OZA6TfmrY5lDcouQq3P8lYIUh6qa+ZzHlTip9sCCdhN+Kck
oiKdcKGJY2TSl6z9JtA2FDsUotWie7v4QAdirRJmEt+fBRJvFCw00IRVO7scsBAciJj3mynIm8Ac
cZ/9YKz1vDUNsjLo6jHcK5zixV90Eq2Unreag8SA/WwrVHT25WxM2zeba7suKlufc0C40vyhPf65
Fc7Jdvot0CqV7IM3Smb70tcSB5OC6ClUiOr0X6NIiwQ7pZwg+qkT5HQLtbKgRkl6L32DAdEmq3xb
hROMvHoiPAozIbCPfLSP5EB2BNHlfPaZWhS72SePMEjDX1079ZafONmLPVf18Y+Q5KtSkIoQ5unk
c7C1F34jJbN4UNngUWgXl33nuqhbFRKmhgpboe9W/tFo+i98uN06Vtz/xVK3sCGqBLlYqTUxDSLg
+YUVKIhvVXg1aioRDjUFkq8B4LC1RpVkr7BxKkvtyGwCSi9/If6lQuaFZpiTcXJO66xjCqu7WRSn
RpYUCb8QAqaXU/TiBjWUmDjtnzQzAvvo1r4dMgaUHuYsF3z0xqEkcXbrfuTG7T+3JpmdOHq8a1Jg
qACRNTFS9Qpd+ItSpczjgNkPW2q4+Oj0PHo9DupzfAXfDISs7Rv6lag2WEG3i3mq+Zv5oxemySlt
ZzohdpITF24URat/rviu1V8MMGq6UKInNXFVyrKZ6UNJQzVGzWb+qeCIFm44PiJ2y5B0HIEjv35r
87ihApaEx4KO+//GbIT2UwaF1/EhFccwDExifFMQNGKUbJKjBkvfmPqrXLf5HCFn14WXt6FP+ndw
DUzWuPwz8z8x+PymszenUSjwdqaikelvvRpPTYBetLRotNjGzFPP9t0krxTFGIiw5ONj2qVH6Xqk
gD7J4MonQikykOQQeJ3tzSXt6YwdNV5BIjGPPFtBNDKycAH5jqebSrEiRqnxbFfEWGubb8MNZ1oc
eycVHNhIrmB1IiqN7gCbAFDlhLnDYp/+CwwQ9IabndvCnB5rKzwjZ+oRDe24NHf2mU4DfPoN77ID
MN5tziGznVs72w6kSFGaRkkT3NYLkFIX/aPh/QPYAPjXvTn9CwXrehjHi2Evad/Z/rcKxClzhFVI
YXNTPXR+HW5I5g9KkRtXVKydu7u67KMG6ec2Bpe30OyK/5fmRhDimcDmAbjGRBwmsIMjWxFbmEPX
3NI/GH9EOEsl7hqks/cdY/mvgrw4pVL8WrGgYy/VqQWYIlhd6bM0x8dY2MU6J+Zi+2g24UB9JLkw
uzA/NIAFjNrfYSBbHfb4xrdLFXyySCerVy+HEX44Q1p0TN286lroEEsAP3Gsa1RyyCAVjfPQKJa9
V6/AfO8YNSoXe/krdVZNuGDUSn/ESbFJNWG2rjcvf0gFD168aMCBilVH1Sh7Phxp+B6XcQoqHA6b
VIp109iG2KNKKBGg402qSx3hhISyPWZr3576n5+4W9wZFY4R1DXMcFFr7Jp+gH8uv56Kn6tIi/tQ
dBMbW9XdN+WuQTeGO47wyDqC5B7tUnbc4G+bQWHhluY9+bHa1CK+GCiZ1IIQ6VhfrQlJLnvqlAjJ
ym9+8JNqM7QTdmSjVOy56JumcufZv0gMzKIkP+X6+gTJ2kHaPljz4sm0fpgi/nAqYZCphEJ5RM6d
IefH2KyowfbhXe0UltkVc/S7fYRl2mkbOgB8yM0+KIr4HocTTjDKvn6F3TuNLa7AygfdNZoVqJm1
PQQj/YetUXSwAYnLP5p0DTfH4E+pOQDahjWs4UosQA2+s2v5cT164CmsSlB/it0sDG+cG4F7vj3Z
DsrHvKXEynyInYteVm2vqeoOBbr3Y5hxsTh4DaupNyyoyDN1qlPRg4Fj85g8416GfWmN94hOmmES
qhCUEpuV78VqCcLuoBbeznTzUxyT8dgThkFQ9piA1CfFeT0UL9WmjCEEbJD8tPn/A/WqByGhH4v5
GNLwmMSlIm5BU/aNjQuQJ7F9VD/brG+o7ilvSxL1zM7G2sxUI4YYl+715tmzTUauL6yFUQsoPrtO
2oHIryWCTbSqblMGA+ZnTTT7xdFz0vHmAMLgv1Fj13UdHT3EHLTbg4gnzniAfM84wxMf/9BqngbI
avj6VtbiWPhrFvDoYI24sYwk/1OR7e9Tv8f8V5qizGESMESzxj8ZXImuJ65kooAhWe+mcr7Yyl4n
9kYLwEh6hcvmXxPdccW5hG5nfp5p4V6RgWd+n3rSC2EfWT0Gd+BTQMSCwjo+WUgAjZfxXtO5I1o4
u98f0uwQVCFVBdGkEg5A59gw9jQ2ObmyHRTqdt+HS/tF984Uxx3urokGDKA1L4T3les6X8wwTHfv
6zSi8TUx+T4NgxS3yLSWOat8712AiQievXceDAOYYlPIWIn8uN/ulnpaG3CIOBPpC0y8oGGUS6nM
mahufxjO7NF7lPjNGD0XL9HI+ToIA2QlSERf2rpTsQqUSr0MgVsTxibC+kwCbM643JYKsS1OSIhx
KUt/2hFJYT4G3r7tvUpFCjzjspe4wX5j16jUKrmusq0wGogEACQgHv1CaRLJhlLw5oLBIMezBvAA
+ia1wsqpYedIrsEGZaZQ2RRNjAJL129p6u4HK6sdAEopQ10xQiWJENzonPsyQmfUh0Jg8L48YcdY
gtITwx9LoEH5BBCAuwkZPZ/jQP1PwaymW1K3l5zMHnLockAUAlYtZV2h+xev9syiFCMrbVPz4fmo
cZBPwKroG3mqWoYJ09sT8Lh5S/qlQFfEjMfFZga4rSjLjYF2b10kYZsraKIrFfNiqM4kQR0WWnMO
Q1zkzSAZq4fwRFecBCz7CpbZS+K+OGKnMpN5WLSqMdJD5uEclGarGOUrA1YDUAAinrqGYRuMRBKn
lwnD9F3C9pZJ0NKPdZeCOwcemQ7zbxSMgsezmVTS9KLhVbOSz4WOsVytXRUeT1LuHvqg1+l2RCFw
hW5eB1JFE6ceyQFNIXqxEkJ0WS2un1ZJevTao3ybRRe7j6cnz5kODC9XUx0GvUeRRT57wcTQImNQ
Ga3RjIdgUoGGM+4Ivhs+8KvQc96uWP86opOivq312LnLZlPE7mCfIwNMS69VJSNi0zPTsaM4IKHR
PXCv3Rg3/s6BLPZUvcnd9uYKGCclr4R9M0+q2JcLV6E/w74el7ZVwi45Hh+M50mRstP05UpbKy5X
KT07TIc5LX+oavKwdd4yIMbMfGzQvddQ7loyPcZoYCFoNkGtxKZsD5CDd6TxxhsjfBXAzhnxufm1
cvrSbgKoW9FOncNKMbX64FRxzIKrYONmN1c95da/2x4L3p4OExTPdRBMzY0wB5XHQuwsfr0W9+wZ
nREBhGnHL/LWfSc6Z5z3Xk9TbdCUNsa7pnN+WuGzu7AEFK/yAVZHCW/njzvxmJEUMbPqSBG5onqE
VGoWYQ73TX6FUydMuWUPak/os1q5hz8wCQiPJwq8gQO1LF2cCjH8kxVTrwLwUNBJmSmgMnsgue17
LPjPW5ZWWVn2RAi3OpGAnTWZ+qzugKgTA9rVlKbFLf45eGgdQ04bc2KtKXzQ7v9zEzOc/JwB+6Qs
wTr3T1A5E9tLeCZE3Q16mGqrHuSL17ZxAGBH1PrDnf6PBCTTc/rB7xMMWmo8mRCStBnfUoF+D9e1
PbjxXMeNPAkRSb5fpiES2WBfblBsTagRsiylMEJLrscpxF4J7BUDQvSba2IZMKhw/u6vY+hmWplt
4KDF6XlIRTAWe4uW7PDGW9ilvCUxmMjcYK1cRmC2MSyQUkwSmmg/tGiyX4kgi7iuOEd+rYzPKSZT
OLxtFMr4Hu7f7n3WQ3bbPs+LNIZCaA7ngsA/Y43wqa2juB2urypRnZ1DQtK/5i6hnavGB2lSDfOL
v/pxapDXSnNxIeh3706vQ6GORQx5GjGVzZYtbMN2s2qm/ynuWvahShGvFyVxy/QOYjWNr+Vk7Z45
NlqnHeIq9eeRAVYrgCoqeO0mws2U2ZQmLtdvxAvwgA+aaAjGE++HjXgPQzgzZMo5gYM/oc4+pCRx
M2UpSZyHAXQO/hTegT0AZoH26FVf+TxzWDpCX7Smyb/dLT+wwYEUBm65mSNRlhqBdSg/PBVWXj23
TeMfOYkIrbxZTTcNFcIcBKTc2vPVVDHwiYPeImbsMv2xqCbt2Hx4+bgvsZkfQNz2ovGs2L1OShFp
AQXGE3JZfc1HyAOguFyUWspdUka1jUKh2thrhRsJBNjCD4fq5gUIVv6FnqoUVTKVpFRnsAbUgnDS
QUIkuLUDi5FMXnK6bUh0fqazlvLPXd1ad1A+oiGOF2WBvHpl/6On+tc/Aq/cvCxYwIuDCYKH8YQf
XuzRyoFY0hHWWjxoWJOxHA76ZR6YiKaGF/3UMibgA7eyq5gTzmHdcso/swbCRxts4C8mptUZvrzt
8fPDwde3QtiMN7nzLVEm22P7xV4Rb/8c+oMC7hPvMI2e+1DMXxpzsS8bS1lwKpu34ow4Kue8TwOx
YkAVcTszLW2OVIo2FdfdwQxoM4FKeU9aNSdDNwhR4xhI6CRVPd96mhJi5L1hwTXY3yE475ALpTef
j3WU3eGnWEfMXDHe1ud0OMCfd3nbaZ2LbJ4yIqXIOQEvLbpKA+p4aO3tRZicLgFadMdnJ/mKL4JT
W7yghltEPLum4bJmoGBH9XXcMlRMx07LfKg844BmGZLB77qugzDOwwqTwFa5b8aC2e/gDKm1KDeW
QL3oLUUInwfCbJXBYlNl3XliHxoSVwzvwMDC6ey7F2AEJFobDRxJl4Xn5zgTZihtJqyyDM6BeHuY
z2H4UNwjggLQAEPXMCQD11TxqFliGSrd0vEE1J7f32TA1K6q3WkHUAOrFyVmU/cFvcgdRT0U/NAe
s91Hl+4ldbSKAoeHbCn3CnqWgwESSuAFg1hf1QkpIsWGsBj7iSwjUnDoZQq+RWt2ODlSpIFeJjij
ULKow2MfY4TPX040Fm/8s4sjf9hytCe6bj91n2owZeLqOCnwOZXNzg5Y9bRPi+ZtpBaS6O9NXjpI
06eiWtmYbLm7+ZwCDak0vjWrqjayBbSuVhUF2edesvXlFZLf1nNptbZROiR5v5XwgK85KglrCr+1
QIqliDIrk80j6RK9OIJHzMuL615Z9dl2KNt5SD7C1YjU/CzS6AuDnZ8OrJ9gZGfcuUkoIGKFXn4O
lo8TQqc+JYLdCbEocd7AJ6u5olt0t3jEA01iS135YEtSieRLED/CM157gy53Fclsq2a//1Pran3V
3tEp90pius6jaeao71VOnzI74wwJlV9NPIbOEi6jf2GY4i71mUGYtEoso8z7o7xnT7W+ZDelvMJQ
i1rjXLCziRoeAfSHICYrIDJ9xkQOwm20k9vyNyXLG8lLZJXu4R7E7IluhK6X9ISp+mfiDcuG2moO
AFG9YIjFUhBHa3P8lstLcfXcxI/qClYQBUJ2vG2XmtcVnkpIvovnTtr4rAOVm0MoHJ5ik20/8MHt
SF1qPSJsLhtr0OTrZRrTrQNL8nB5T1Xrf2NXpzf9hwCzf43JbdLkGZ6z6f7MVCZjtsACBed2JH1q
ZTOYQTSDzXCPYuxJ+yhvXzBqBuQDTH7oWQp9O9cdiPjhA94uLqK9gT4ShDxMOONEhyHAVFGv39S2
wcov1otn7JFEo4MQDJ9YV4Ng/DZop4Do7kjOGpRszwnemSMNAYKfUzel1uydO/9caKZDBRooTRXF
npbH6K3yVskPu12SuFz+tWpQadfuVs1dXW8h9GlWdTcrF8TSGjAe8SEkQnMCYiw6ftRUqGbqEW+b
YFBkc+94Mrp2L1gRLIwZjo80iFPZ/Mvmf1MZ4ng0fYee5Jg18/VqxW1Gbz3a+CQLqymKRvOYgBga
SPHjXKYpnyd7gxoCcZfi1JV8I/SwJURhxDioLhbT7+XV+sIM7CsZxRcAzx9CJ0vglDBUojfCxXRo
0TwzlAr13yNq1kNW29U8zMGN9nGMtQS70jm8+ZJG0ydFUA26/GXX7aB1+TmcPgJ56mX8eHmIgVUG
v/eRXE5B1F0VmZ3ZLROxoVeeiu+PetGCfnHUL0LDMEBijTvkxbWbo5HHQz/n+SuAnKdJqVYHbgl6
tWxKNJT2cEcXObVw6HV/IFtcxGhT7wVGMkyPEnUFTiAy/z8LT6KjPRlU7pCZr3AqkOXXAlPXIhDJ
0iaHqt0MfbBVz8SLOcuPWeHWtzVeS1aXCFyIGd7stMtJrlZztrHnmJlIpaEMMz2HIa6U1TSXLLpq
VFfSXCiv8qWNE0R3Wr3rlO4f5xZTJtp4FuZaeLKwo+WxMVKvoO88YjkZXqFlhcJ1BFb7dCISjdjM
pnj2c7OzEV2HwA0kyjmXlYcYYIlwAzFJGxzQTUxjNe0uQimc0erxFX3Icw3gAK7BhRRPX0VWR9LD
r1+QFDhXIAH5WywbN9wVw2XV45tWteMR+vABYgwgt0ZM2sMFK8P/sK2fkEHNsu54KNv8PImt6l7d
t+g8jpcmGRWcrjqALrxkT+6TtMqcX6sdvDYmCCkhTsLi3D3vDpAJ8F/0PZY2mkfXAAACQWZvRHcE
IGoV6fLMMNZfjcQOL69LChneWiv/mxkGIeuV1Lz5p6auO+aeJLYWTuKYswGQkqiKZEIsWa1LiIkx
ALuqyS2JeXkGeRY8qWGeENfjK/UsnavTA8HmcEv1XKLB0PaVsIV3+Rl+JJv26WTKGCWK9S2FHMaa
0x4KrvggvFe/gLiriYrB04QVcfiuQqd1DokyyyfPGyOmVUZpahRIN0obHOvOJpuDBvGBIoK45tTa
aMT5KGQk9Bv5WPy3bu9say+tFK1bXyBeEdSL0q5MnbJ/OQC4QyRJqSM1Qh3a2h07Hf8eKu+A6aNr
uAbFp7Smr4803kmSx11H0yTpdXVLWBHgM6unilNm/gCUfi3L5yoYgebVExolMDZfAodrJtX+tj+a
kRpTfkdIw7P7Gndce8w/srEntvLoqwMweqiwllVdKq+oS6YAroyTU+JkXunAq+uk1yH2b2HS0HMg
AJUJVNZ0v6akyayrMhSU2rcqdkXzFmVYNQ3o/RHASJCHngDXQIDRWhoGyWoyLJNYqym4268Zp/42
GDQ3Miwi6l8tJxxmj0J0X+g/qbWnX5ODlJgWVJAGx0xkJh4bnZ26trHMK5jMwGLB5M/XQXZpur26
hQ0SruzGWPf94RuZHnN4DC/Km2b1No0Uh692UgLD7Q+NE4soHTBW/elUNdsGtW83Mmj7cg8XI8F/
JEtqsipooG6cPTdrGDMj32wsa2LdLxbnn+dOdnwTZ0XvQ3gH9gFubBLZsqrzGKUwdHdUxKvrqaL/
1ytO7c2mMuiYfSJOPjll9258EkJVte1+J5KixLo1kbh22MmOV0Xf4FDf4/ptvsUuIWjRl7E8N92o
+b/tRG5UQYwcPjUVM9bTkDYHOfASm+/AssaZD/0H7THec+s3bo4kayIJGXhV7gJdY018vXDNIqIi
3nNCfNS1KVrEJ0/wHaw3TZ2f4Ku8BiFJ4bpYr3vv2YMK4JVOPcSX9xYmr8VqaMRQFommAw7LoRGY
GwgEP9W4B3PtWVdDHFz3X+UW3rtMqZpBkwTRQYvf3/kA40mQi7OO+exsvMKfsE+/Mt0efcX5y+bU
Fjp4xkjUYsznDvj4kzUvM43GItz7NZoL/G/aFqfKMUlOQH0HS6D73Z4Vex5uZYwQCSiFVC8qAh9B
E3xwUauF3jhbPLONJdnIG+CCpT7UkrV9d8rlQfvwntpnhtT0pNSu7r4pLqRE4T1DvX791325X8QV
VwyUKCvfceWMuJf1W3ATRgXmD8rXgmBD/WrkKYyR3GR9rVEi1o0Uq1SXM64vqfYu+6AZ21TbZWYN
F6rGQ/KvvfPTTQIbAPmNm7IQc0VpR7/HEAbdHNA1FDlGaW78Z4mYSW5kfOVBtlqGqjx3jY5+dsv8
1LyIMWMHQjwBqjUP+OA32DIMml4shYymeJVmLndXAhv+UpHwI7TIDQiBfUuyIcIYXUxzVOlQgJJ5
SO7X4JkWSkbB6K4oE1gOb+pfT9rNYspmz8e0sqNRRIj7GPPCe6RFJC5DTWoPvM0TqQZtUcng55Zr
dYIlOKEQSrViU4nTsTdRXxrTNRsCNnbNhjPMqH4stwml4jnwk6vuzNHcIr5VzdlpnW1UvzCO0V1L
rwkPxST/Hcs0DFITSdBsvJtozVW4yhMjeKxEni4okA5odujmPLdWNvSqyJ61GKyFNCDIS0aBDvyR
ES0cfoUHTeBkNq4W8TsVH4rRLYzA+RQBOuxcQsfKjCZgo9ZoNWrEuGopCHu4/ZrOxhADgOACIJRJ
RpQPZ0Z0D8rXLZkIiKNBiPz3rPTDWbAjhZOxWF9ztOV9zornyZZk774QcoQbcLaH6aiOVLTE/liy
U7rIcpNog4NkPzZ35PkLxufpCF57kfTGH7RIQbbXoykWsfu7fk9rKWdVPMxmcoPoxEe2qm4gcV1c
fR2EI25JEmjbfEPbBMylT8NmeyhqqsJ+Fb3rdQfgxBl2dkPfFCyeqLwupDvsP9wR3DNR/WUMLzR5
Dsi0Q9NY+2l7gX/0jZrHz66JyHPZ4izV4YycBRpFkk5jBSN3vN4jm9yGWSu4rtZAoqBK70Mrm/fI
ll3rcxTCkq4mf+o5ZQSM38ICQge5cRh7ggQMJgcTd/KgnO9j75FijUG2NuBfsJZM49z3jGjKjjAU
hYLMJVWTgj8O3cCBT9XMToJA8WiTpyj9Dq7YgI48ckBPK66Nw8UPo2jz57j04OOk2WjDUvpPie3C
qhZ1gOvU4X3bzPE7D4I6uSEWc4Ny/wRVd9VU7qKbiTh41NTEUVmGgN3M/RkWB66UhGmpzDD7iPmd
7owdOMtRumbDt8tdl2SN9DM+Rp5QDrzHR6+n10+nEL65DsMIIw1QyA3nazLJw9WD6HzCv1DHMQBq
I0dFLPy5MZzZfprR0S8jGV75LpQEEBBFH36sD9x0If6sRwJp+HZ6hYmtwD2+dVtkxisrS0/3f2kS
slqBI81op5VeXcdk4xhDIrg0a1UfibJZn5/ScIklPLgqCJPl9/PYuC076L6hApQaQapzNNLeCp2c
6udCPHdY8DhlOIKq0dpDEdplNp+vBM1L24oieMGKHHnlDYx8/c2cWQpeNa53RCFVOjYVKxmDyaWd
C66jKZNLatwGZDEgb/RPkBcEq5c+fDsEcSL+PkSIuDMNvcWhwqJS3u+KGARhAweaApFL1vLeflbA
XU2Efaua/Uylcd3I45ioHp6RtJe+kf4C2BZrhzlz00xbxER4JHi32XbkfRvGm72yWgg5SkwA2zrX
BH7TX32H+Ykeyuxpf4hCQ/duF1uZIDD/tpON+r6rYMyJT7mjrUL6Wpl6DTrLkzGG/ingQz0rDc/E
XvpC1DNZJBZJDuMUzLaHV6tNynmtBNxR5EBthsz0DmwUIGTtnhKhc9Rs8pxhs/v/0+2LKucvBNS1
fLmNqMDymZ9eLHLs/8K3OZmyZ1eWcp/C3WYDEFHT95ZWKz1iCFQnNx8/j/g0z26Y2thjsSYZ1eR9
e6zKB6citm6PgHj6QE0wmAqcvO1dZeFjnF/KxEkWcZEgtjeKXTBtpQKwx9RcQHr+l9C3GZj+xIGo
kNWkedCmGkq3YJmS39f10LlHfszSnPXkDbItGMjDXiCLFcBokmlzi6LIp+CbuTaiaOwZVv2l1dWf
7mN3PcQ//kUGh8UGrE282aj2Qws9z90EF0h06AFlyDeAykDIKlgJCXqKUwnHW7vQ6rClwPqNO759
xm4GdjU5npQPJEaoAo5d77HStSli+CaQY8SmtZr61eqUhAZzWqsAfi4pfRwbCT2eO2YNCQYyzges
dtO9SoI6Yhx9WHZjDTcvMatYaEKu4ojlbeYPyJAhtJVBNEQ+ZtwtPA8FhMCaV5VQPixmfaNTOT+j
KYpaKMdSIH1478hjW+AipzjLuDACOBw5W2TSastU39VmS64J9Sf1UGgw/62X3ujgkiOr0EBiPDM2
oBj2hOo0IAra2FdG9D7TZ3SU2BjYNN2XYPJG3iI6AX7ht3hqV6yoDQopihe68sxZIjFHHrHQfAUK
N/pSmmZAvfdC7M8++frMIGLdtecxwaPP0vJqtO/g/h/Pm3ZIFjMc1N/AuQD80DbUtuIiR7hcqDDe
QuOcUOGJwSEp4lAG/srA6nZikg01PrVNuSbrYITU1xLjwG40C1C2htX7ozmkaokrL/dd7ZHJko1x
EteR5h3zbJClJxi8cenxGb18dZ2KQF5yZ3Mkk6AEiKcYU4p7KPbJOfTj4Lg2DzXSBLe9HTdRTypu
eyXdrgykovzQtMD5AMG3OYxOSGaS6QdqZuuZ5uBvTDnM8WHdYzBGPWpCHbVa6LrigEAk3Ij7hncp
0vRlarq4r7Yy0n91gJ3UZLBUJ9WWVM61UvSYSHzx7RnCYfFi22N4BTOAhRZfgnVjVhE1pskLtGGa
kl6oMsMsKiiGlNiVIemv8SuWDl/Ih9V4MEqPeZsH7fnT8BCQBbBU1/OySos9Wo4JMhnE9xo1v35P
zGxfeAg/7AEGxdyVGl7COzxHd31AiIeqghr1ys92y3t/GQMzpOso59H1GLHNPi5mnclVdljRC7iH
vSZk42J391N5QWkoP7OykoCT61DQmINr4/J2JpzmJUphGNJ6m1aWsTS56WdhKLX7yc712IFztNOa
i4k8Ij20tfhZfd77HqclbIWz2XrsLscGMG/XlsRPHxLPrz0JlSWYYQ78YLdudGzIrqWH1p/xkCEO
BQjC7FR9y2fRwFPYRJMuDk/SQGwCp5TbIRMoYVUkTR9I9eVvGySn5Ahjf9hAZZTWTUDfk966BBd9
EtRjcqKzE1AaTfpOAuotOg1YhUPk9u9SlraocUWH/FevxyhfzfhsuAHJGeFfq18ay+YVJRczip52
xo9z3IlztzAsGbLTdU8/jfHjPAKobxplXsnKc1y+pOOFtrvFcmj9zV6/Z8oG/iOHFmZja91i1MAo
VUZXBubQzg5/9g7dH/dlEUjtL14/F6y2PMpBtrOkX87EOL9LeiCLPIT9Goh8Ylj9Ksvk9g2vis5E
msMXDuzzdFzg8e7eLJjyMfcrGWRYpFigG6mmLGkXj4v3qbRIhtMaE3Sg/GTcH9kJLO+Js73VlOZH
Fp1MbS2ZkfG8pT5qBxkPs7gbOppDqVL09wRYyaFnspyu8xC60vYijgqbR/311UGOxDJ5eI/XFAnG
kzLT/vs8IkECnPe4eThZYiLtGSiRiHqaN25RgjIfnVu06OZ1Ltugc/wdUojx17fy4g1Tsmkm49tW
t9TtFJpm/EsF7zo7sVjF+pWXcugqbUuO0F67BSrifedw77RrcMY34+OyCA5NoZB2l18v+ytIYBhL
IFqn1GNUFlooth/oCAIbTTFMkxerwOuIqDUtW5X8laV0I5Y+gwfKDubMDB2R/Jl1Y4BBg5dOagC5
G29X+nP4kfqY3NtU99xrqhw3TGjV3QF9gzYRIeNdF0FCUYFJTLgUJJ5RD+RsS0CpOkHB2VBHOOSv
e6vzFhVMZuNPmZ70oi8UNdNHXSOfSNhifl2cahWqb4oLjrvtfjUT7ruNuE9HY2w7yF+pWVXDDOGN
d5yrCs5wPiMlggzdeqGhwTuozb5LuMX+emWit9NqyzZeil+0epBfVCwukg73PHYZfMu3c0qO/t15
zvJqzEcIoekCKAqJEKyzFe1kmSZTX8E9e6hW9yYzngmMFjIyy2yBEZGEDg/PP73y9B178pQVe/4o
i5Wh+MGJTGml7MlcZmBdYQnd9q9zs8DPA42dQMgjBoJ917LDvc0EGZpNm6iOBP//5Tg4GV2v44+Q
FapmCIcH2Tm1Toh4Vd6H4IMo2X/GC2SHSzbGl63OeWIHi/Sc+tEMFSsUo8KOBVRJ9ihM15v/bxi+
GZMssAdk/WIzbId4s4mhRT3hnf5DLUNDmF+M9kzHDk/qADMxvUHJLtgpnte3Js1dct4yX7DrbJq8
SFPE8bahEC7x6os92sNo5DWWDb8OaEeo0QQjMyAPqOXm54x3SHnDcRS2YwWLNvqSpB26zSenmAlA
8lIwyM5OWYdEz/E7iiRPDxMwSLolVpDcWUQeyZGl5740UNaqKkg/E0NtPJ6DNLhEC6phgPLGSobf
DH5yrDcpEVelUNHOHB+Di43aQ5ZkOQVnaTrHtFRF3gtPMh5E61rTIY9+hCk6gAAZkva8l3Og4jO1
+U3E3Js39NglIrBTTncs/enmMI2t9r6r3OR1FBVP+bGuJulGkHxmmyNbNQbn8hd/IMMUhg4Tq9U0
04vWkEGkWf0WaChOigkfcFg8NJDjkKvK2uF0l6YG4pr/iwxN2/jsBElQvvctK07NlCy3Y+HjS3fD
gRU3p/+Y1OOXx8LhvVdr3Xea8cwQpu1VT6ea0o4TroeCY5CoGvxGycDo+9OpDfsq8z5uAyD5G33i
XldPG/AbSOyFPszhmaF7c6H9esCIdoFwY3oNagrjWeB/bCoD3ws+fY1uuw/KFhbP9wlmq5B76bqY
3s+MfsrD+WdDzTP+Q3SwI/yXd8pyOe5x0azZLgemVnH2fypqptFW1UxUM5OdpyjvoCRvZJVu+tlm
R9OlWykE35yDx7Zjjc/tC021F7pyaXqCwigWs93son4UzYDOM2KDhhAJHyveaGIKhtktIzvV6K9C
CERuEQckZpYEPYjrAsnoLdKn5fcWMTr42n6dKrXaQZpTgsT+D+leuB0dXr907dLN+qu4IizZqDcj
70qmnvS8WluqJl/TY9yh7jKlzz9q/SZ+30cC4uCDQEWO88zF1J2IrMy0BpHABStbrodJH0Y8Hcqv
kHgfoJEBzUzwMWgDYWl7AtU83wyGT6b6QSiJbiKU7t3kK+w/NUYO/hdGKTVKDokZ/emBW98mLRun
guxXsAHHrI3XAvr0gfHNHlcDBCT13f81rBPAlE50sGoPUd1lW1K1SvPr95BZbaH+CUh/o6fakzRG
8a27WritKreJPQiI7L6/O8lJ7d4xsFK6fTk5B3LdpGI3DFR8M86r/uFe1OPHJwldSBL9FWIG5xm0
8Tb2Fg3Ges+tVt/f+JbxmivsIOPNmyZoH4Ncndkrir6SnV+xhALZqdwIvz/twmAsMNK1vOs6Ktrw
cUU9mjsYiPCIJNPH/jbppnKwxlJYSj1ObqHGwzyoqfIWyaMe3XIkU+rK43QmjCouLpMeKl36f5HO
qLm+dpwbBORnVbav2wXoh/NI8/6z1lHvsYUlnsK/nMJO9IqDSMtjlPrLw15Lhjc0OLS35JJe9GYF
qKqjNtbhdnpL7nJxdhTA1Vjnx1s3MWAqjD03pp/SeKigMNo2cZBnd43yoD8mRdQQBQ9hDCf5oswk
7Uzxw+I0SY8zr2waCony5Rqe4k4VHbl/t5h4M/GgDpE2z4rqJ0vm38VEElfIsOJYKXBPn3/0hz+V
GuKsV6TCAd5NLgJaycoBjo0fpVx+4BA70/iocUQ0J4mXi037CXTSKPMxo/HOCP962qemPrY5g1Lq
qezlp604KpjVGTLhI1USpHhPXi7n6tVXgOUsZRYL+EXgqHfDUtzGG9inY2w4UWnxFrktGgZMc0VM
X3IkijDxAh/S5a1oLF8DGVsOixZmjASMtVvW7p6QQGUXC6rkyaaR0v6/V9/4WBLNydxnw74qs5gH
p7pE026YfIy3Mkidcju6yWwtEqe+lWvze6EDYNJurrME+vfxp4M9K/0pBL1vDKCJW07HsfdY6ZUY
K3HUfPsfW7QghI7/8QEvyyc0O52ieVi9ISUiqkqhW8k+7cr1p9JVuKuTcnGOTd6Qvyn22x06fLod
IQhkw2F6+txglf2NLx0rQgU5SquQytSY7JY1UWMbBcuWssV9R+kq7yktqwfTADbI9/pH8i4ZrAcW
4QNu/gVHlabDShx7R1VGA0Q6OVm+SpARzni5zToRs3eT55PwVnaHXPoJfesd7VNJV2cuhENsKT0n
CvB4pP1sLj5zSJjv+vJuUtWuBvaLrKQz92WysBddmq8BDIIXp+RiNC5gl1xxvYivq2Xh6+EXuUxL
MhKAbnStgCtlAgplgqLApKeGMHHzaS94Zsce/RTmO/EgqyVHNms4MCDNnHGMl8hrcx20LZzNXwje
FZb/buozBjP6/HJlXYl5pP6o5J/ANibpAd+EGPvC9zPs0cxO+OiBCl46tQ5zIgIlpcTBVeZcTmxe
3LG6C2kGC6XB4jdW0sNaj4oDYROX4WTmFc14Wesu1rDPxemNiAQ4rm4WLs830KOZKIVtcgnGbcHy
JHLIBUUU/5Xwv6vG39l6fXrMEWNMG7n8cC6/r3ObPpzHucbrxbldWR5MXoDl1abd9d7q/GUW2pP0
xC5xXXTfn9a78agYLQ1G8RnvnpD8knC33RnvO/iqw9dqMK89XviqSIq3ngpraKHnjJZUpQ14bWfc
qrLqkiTooKPPiTqd3kjvYRuk3eKSWOd6iOqnIzA5mOG+hui7BsBmNwrSRMn09KEQpVGwr8C74Xed
4YEAzv7KHFDirodBS29/jwnnSgUdzzCYwUCr8m5urwHRbuxWJWnpYJt3d8mDgfA2vsQhdMbpz0S8
ipSWSw6176HrnPuXzBPaTaTAjDH+TNFyeakSYAS0coSBciq9i6Xg54qHjkyqL8sVVMuUDwPY561B
bFX1oltGkRn6O2JjQ4K2F71x1q9qMClSMOzoHK32kCBai+KFPGRpemX1exlj2Dd3vGnp/MKAHbJC
l/nlvw5wLIB0ggNItFGn6TH9mjWgB38pkeMewZDLEfzP+Grli9dA4RSEbDQN0K8MIGjSpEv5v6yr
yo72Bb2E6hapjdGogu6eftjWoB+uq1+iWiXRNtgCJUbkt6/K7DUMgeOto0PFSBNGsZ9P8/DAj5uQ
Wbyuoop+pjgtc5WYsvdU10bQM0+kEJuJfXC+bfrHf2wsz7my6C/IhmktaWYneJlkkRh3vm16qKII
YnjuDfnzyP67YnTaGUlgsob6G0uiX6Thv8N5lhkDvMRziH2ICuUc/EvtQ/GIFBzX8iZDbmEv39Dt
S+23xbtk+rEKnKtmaVQfA7f0gVvs7f1Y+wgXhr3G5XXwQ+FkhT2gcNK5m/7+6hMCmQmaeDbkkrfT
lfeOdVCgcBD7Tse+Nk7HNRSn0cX3/HGVwYRLeqkeSSfRui+7TaB+53OqH19yx9kWFFKlEgPuNo4F
+yYi8jpd//3qn16XTVlR7a10qYu8X2+B/+z4jhI+Xj2WsbtvmOcc8Pb+tJH43mKjLpOQRqssSA5L
qkzjlZmOG4vpZDHbg05GW2XxBtAaJPiJKAmu4Ys1OlHb2/N0bvMdA+ZD30GdNhF9EMMiV8gJ/oFa
qu3hEpjzyD8ppG2NVtDlsjVAdy+RpA3GX+U5grzwoID4F/esc5HkBxkpIxuJkdOdywiauWqjFqIb
nbvEzQS1d0wPsOKH+KZETqY6yGTLf6IPmBn8aMUuIjoN/HC7C4EovtA+rLwVWe7B1hNQ7+5/48p2
lZKNd22emGZiI76v2+9oKiVtZ6j3MI+/sOqgfG7woDkE8+7gCOyO+9HpAF4ihq3inVsk5vlphNsx
FsPicxm52Br/tACqbGX5YKua4wy3xlb//tFoDgT2tVLsErBrkU9gupwGY/vtDYvliOYbDz98YlPa
JdkbKtZHhGiy2SIVc/YxFJCBpQ/+P4tX0vZy8wykSuKMOsWGLlI/FePU3mrBXeGta5RHMP+y/l2x
pJBSMvDgQcECgzLZqk7MKefcNsS4yd3nY4RJk7BROjvpLCDGN/4GjajXE3TIhwPGvrunQIaqjn/W
c4bqBC2a/DM/AnrZkwf9NloB0p+MxbWh0B9HzZpfPy/sY998ZrjTqi7QqIarywcn8DFRInJOIkI8
S6vV03kL7XEpQ9xZ/wy8fyDArsxAsB3k+tJS3LGHoFrUye5dfJ6+ECWPi1whQ/GpT+nV0xLfZpi6
2AJtXdd6KQQmBGTjUFCVEGDLBVq43oqH5L+c/JqXFZWXHXWVM4r34XhQB69kvj80+rNe1e0IDD/W
0csBxbl4V1ECWVXwgIOsacsOcl7yKcFGy+1yRk8AjwCMJatIYm0z0sjlVbsVDIWV0xJVJlOpmXer
fJX7BeZKAnooPbefzHUFgv88NbepuX4AUzfyFgad6AZkGEPg2YJSOwN8EIzFWSAJfiksP/i13tCg
KYk6zgfrHgDTL4fjZjLAgExP+I/rKQVbKZrsxRt7xXThIPjhNVdEeX7LPpKC3r5b1woDNeE5cHb6
WcIY9reAWe1cYpyfbVWbOVKbtM77XJ5M43ppCKvveNCfjmBuFfDmsxL1jINBeP+DCVCVgTLSLRX2
aLKeQv37Q2WG3pw1Crs8VaFN22/Lf6kKb3H1x5miNvpfyJvvFti+8vtuwHa5jpCiy7ZcJ9VPmDFx
+M6pxJY75rlsHVAzqkzJpb9JCkVwCjhAWALwlfp65EL0I0MeeeDXubHP/zRkk+y8xQlUcPbSIiNv
rONrqKab/kyHhJVkbLaNpQLxCy8+jhWxRHweDqS1hS+dbszSaX0ra4JxbQRGxT9MzlfLloNFLzzM
phmOfkxtDICmYOuoC3lAWp4EnW38PhAWcVYrILJkMC8cCYZFSM9eksSlm/amGa6toOOmR99s3mau
NWqStT7ndagARgyToTXnPRwxubWUkyM8Tmpt2Q1QmjYZDFQ6Ut3kmxqCMURAf6IAnR/vpnRxeOMg
180CUuA9d2jow9c+20DcorQyFmdc8EneI8dCGyfixQu+AQIDxVzNKOdR4mWWcRtn7l7M3iB+QNLI
qvHMBx71+vCViEftlwUGgxaEvkKliFVfgEFEn8HNYVDFsZf0vmO12Hr3wka4+5pYVi1PnzW463xU
is03bRRlprV3WPx1VLqbKb6fza85u7LIypZABlkP+hZyiCamvo7ky9x1Ul6GHK4IVVtM8v+rMZFJ
b84deIJPQFIMOh3mzM07SdJ6/AoqOCXddw3mfL52dn8mrAyYJ42UWuA2/97E7TyPR4LiGSCsyBJ1
eoEd5J7or3Gf4/XAHkj86+jw/paELcxFQbUNAtuzbSyMWnthv+RBxUOWtw7u0eOiAqGvu1lgQaQM
dEl4ll+egKHZowEuFnZ44GCbqf1X2aX4OmWPjJH6A1vMuR7KjQNIiD3yfISeMHehALPfhh4Y1kUQ
J9Jx8OiQ8f0JGL/rPEzJgTAQRAwYoy2b0a3+3a1/yoEHYIYQhA2GUl/w9UwDUGyHwwAWNrT1ME+b
jeZA2QLGBzMo1tnsZqDkPnE0uLVHHw5N52zY424TCae/I4jj3ENiZwIczgYyu5A96JAG8Jyg6wkN
z61TXhs83IRIvH20iG4QxfyX4RqHDfcYCUG3DEfm4MvGK8V0l0lsnhKCGQ5ne2ksinB1XvpgZov0
PtBj51rC5Jl37hbWRJiVTJoaJNJfJIp77PV1haBw9coFFkJgLS3hbZCIoN5kcCqnXlF5AHmA5N8A
j2IJQwdY/tiVuWKCmMwp0Hgh9Mlz1g+Eoefn58RiB2HvZV1IjoVOhpbdUsuTfs3OcBdLPcEehkPc
H4RIzbOsDD8Q3iXR3xAdo1hJI5AteXoqs1v0lw0Khl6P6EO7yKwqE+oLtIhUxffoyysjbTVl2ozu
qLrpOnWgpwxthLC/fMGwMEGH5AotrJnSa+UQV25jsOBAdMmpmuCOJt0RJwrIWSAg1oQxvuexLnNW
geAotZD+EtIllCDe4Th/PoBH+/Phfr8qmmiM0eV2o6zC/LVtZ7W6lirvavnOljAhsAli/TRJQQN1
lWmHLtZNwaJputtXL/QZci4qbDoHWsgpM57aX6Bi8uro8KUFolz2QNokyOUKxq7RaPAliGmJG7EX
8yJDmAt4bv267h8Y15rxPbzJz90lDIBch4EgK9U4KEKZU9uWGkUUeNEUo9nTU81FMTPqbbT1R5r7
wzwRnJ+EK41WjK7eelz7CN+iNqGcBfNcHY9ZoUStzqeynlc8/TAOv3V83oAmQB1YZfbrh+Et+4H+
iwELMA1AM2YYwG10z5OAjHILFBJi7NO6FXrNusnm3cYNyB3EMOuRWoEtGnTOM5Px2FSLikwC4sHu
WfjlBuPbbRt6q994nqPpC077VPcOM2jeg3qocnllrxYq/kUQ7lWuli5jMNNevGLGPdnnm9oGLnLg
XH5bVcvd3pFWowXlkwFErHwO4aIzwgTbwkh3zGOQPpIZxf+FwuqrVZM9Zkw8ARsEE/3g9Kfbi7h/
ymjhdzRAoWjKIAEH7rcws+JHCNAIFwbZ2QecF0udeXsBKbMhMCRLWeMMaSGpEpHBqZI71G9/yawu
nGUcdtWKhO7pqdnYWl+cLPA6GTmhSijCM6Rgq4IixPKgkEi87sWMLj6JywO5jJCtuNdYVYNCWYwe
fzS/8fG0GUbj2U7Xuo+jlGZqEruSsLIP84o8o4Dw0XxFpfhRVLq1UXbA3akvmsLNMfuAy6G+MUZ2
ZCnThm+Qlp4KzebvDyXE1DzrH8vSTV3KS8fVJdfq0oOMpBycvJ7nwZtEUZBow5LGgmsaYa5EMLRL
ZgqeC7nG5tydJmEpEsQ0tZm9KIcCGRqmpoDndsmgCPeZ5tiHnEvmEwzojVJAIEmelsUqhw1NhMwK
bv+x5nUy9rgM3hXO5aVGsG0yui2fSpSJ7me9ffJDnRrbfEC1Pq8ukOCV0nySBzcJHYevPltVKNwY
I69wKzEQK8wGPNI6FtBMEGWObSL0pKHfZwtnohYNh/xmbRjlGnwzKaS0XK6ACT949SEfYi6HVg8S
35voVBk8P49gDd9o5BqEUFToLwhleLH/GhA/xmXhgOvyPjr8NkKGiorIe2rGIsN8cVm8akKOfYk6
FdKMFuqum5o8870O0tmp0nh9KXkJBHRpkFtEHo3FTpWi7TkThPt2xDHbAszRr8HRd1RvH7YNvp5P
j4T09P+lbR/Vfi1sUf0NrztSpvHyw2pIPSYef59hUaCR2CAMy8Bq2Q1hnbgbji1/UEfRkDD95V1/
FygYMR9Pi30bU3mTSlLL+IXBKo3HpT5rN2D0p8BCVAOtd3yfLrR/IDXm7lBwjLLRY+Y9asI4fc1n
29d44OfcRxve3teiMYW8mztn6UGi+xhn6wYjwzvUpPN/QTfY6seKnFBpbTXQq2f4KsMp2ZsDTDuE
KG8k5u0cj/gza5G8pZjAgXXWn4aulklC55/nkTFRiLewWvzo2y7HTU/Aoy/zQvEiskM84Nu86f4z
KxgSkjcoXRYbeORzJ6NicKQ9y6ES89BycS4TpZsGRjsEnEiJrQcMQLfLdtSzUVOBSMmoSEDMdJgO
kobcxasOPelL9rn0VyJgabU7aDOkr3/KPraQmYM7xOPVEsnVN3k6JSNkTaWq8Jx/GESrwBSryA6h
BQcXE6OjLoXk+WsD33EP8pfenk2Gsr4WvWCetzpTCPSm9f4Yilvtr5V8GWKtXp9N7tNAI+0xyHnL
1LRj4f511KuXVUoqxX4m5gfie5ZUOrrZ7snIb07titvOAxt9ule0UOyvoqgFxjPFT1xHrahrCw+Y
FZTvrhsWLpZpRaZbdeJD354S4rdt3Mu8VzM55UzZR1Ct2tW3hFFi7fDu8rTOYZ5QX29zUXfI5LhK
Zp+Yghzvh83MTHcI+nQOzOqYpN3YtnUV9BRsPRDc3mn4q2sxcjr7GQM88+977KJHqKGXkmz3eQB2
otpUO/D/ORVyWr+XI/D70iOvv3XhYVCFiENo6bHedn+KTIBupu0UGVKUt9jack0g/VX7TeN/aWT2
Kwxey6/1b0PlMI3vTxRsC9AoPf8RosUyGWa9CV9ZPDdsVQOqH+orijxToZHMQkukhZi4cZ7oQ0Vj
WyRQ3x/fXd6sFTfDNoLfAYFJJB5qNRjsMHF0D97B+rLBN5+fPaybY+57KllU+ANDMvdQzmoGqcS8
ZkbNnylLd63o6fibf71nPa55O77ToHO5cMpbCjyU0OXjRC4943sNhZDYcfR0814n+taikrk0ghnC
Qxg40XJClPBrtPt63hbFverQekyD/HcjkpSA0snGrb08cTyW8ygLTG1C7t/Yj8875CfT1mWUxWms
PlombQahf7LGANwCY7MYcO69vBRd+q8mx51kuaEzwxPm7xuYQGYHhmAbenso2Pt76a2LW6lfOZfi
lNic7DsudCtC3VOG6hBKBLpq3X5EPodKZXgVG3VrluGEHLrtDtvGgPyO+lV3YKO2py76Bw7y+E+z
SwTIFQ8Kkf40pWaY5GgQvuhzxITavcERfB/rx8cfdPRRIm1bcLexFEuMzW9zJ2nSq/KwrBKiGTSy
+3ZHxPFePrzskhL1u3/yrIH+nGYzwoAFY+Xxqm2ZA7edNidEVGQNP+mokHjxKwks3DLcIz4wv+PG
9/6wQxk1JuK4QrhZNTGcamTJADZvt9fs2KTC1xcYssFybKGI7OaYMr7NZhZNcyItodhOvefg2wk2
hbfBGoxhY4Uldgo3PigkzK33jOJ2iNcm73ZO8wQ5H4DL17Zw16F1c7Z1l6XqUCa+DyQzGZr720nG
5hPJy2EoUlrW7amPd/n5R3CKFaWoxlyXFwexEhgnNtP8So8Zy+iDDt4Rl9cAPqITHYAAwXoUHSN3
jGnzTufDCLDVmI5ojTLzkZLSkyCO8cHnpjdXeno3b2nmmf0x6dX/QyzfRsCDuCV8RQCMUm23rVkf
TBd86/Vc+QnnN1+bLIcyaMvdaI62ohsWW9E+JhdIxKmWKhasJPXtcwRSb/z7DpZTrpenZITF9T8R
bmhSAxki5oxxbCpjLC+92HtD6VukIOl/WGQyGmII/y2b8QaBmeo/juYQ1UCTcgCyT+4XbI8Baspd
Oz5dcpefjnQV/Jo81hfIPIfX8SNIIcutU5rYstcFaT6NmO5BzLI/bQdhCdDgw9kuNxZSEBtb7wVE
jsr4VRg3a2qbIKUlsrdi64YDikdjjMAdftWUDRExYgDVasZZTUwAgN3Rng4iI5NZZefU0qlkAdig
7s8RjPhtUdbuLk8XdRxPofL46w3xRq2dw4JsLlVqAo0bzaWcl4i8DyiSY7D1NahkF4D1iRdU7OSL
q8XV/2fod5QknhwUwHW4Sm0qV6rTE4/Wgruf2qKwLBwdmZ2ts1F5DG3WPy5Yv3saJY+V2UM9Z4+r
aPciQVwABElF70WSP21FiLbUBKkyNH1n2Sfntl2TKLdrnAsUIssnflDnsR16MzmkbMBHpP/mxPps
GK24w5BuoWa1QhPZ3fqwzpEP/W8/AfHebNLLB/WlEpdWCo2Ry/66B4lFiJ5tEztWZOD/bxZtZxn7
ObrV7/uz/PwkNgsaNvLKx61Ik5bFxE+nujuPZgdIFi5tnm9o3YSh23pYJDc/tQyvv+cR7agD8r/d
68zoynlbHGcq3hu22SAuWlY2I5V+uhWa/zyuu6rbJzLVEtRADGGpFbslOk3HnNTsSJQ/boxCuZNE
Es1S74T8CU4jub0DyqyprMccKW+dTtb8xjG8wFKmnIdnGvck7qnOTQefVhHAKgi5hXWX46FaUp3j
qjIHX7b0DJfZX42wQwY3DohGG9MDobXgKQrRfnu6zIIA+ocnH4f8uuGjJXGQxttzhlg3Jy7GrV9R
X1FR5ZAhhxSazJAgG6i9K3wPsczZOnLtUkiOf+T8P/wVbpHgEZ+HxbKW+okEwXHEotPU0BxDP25n
eg6PMsDg4bLFQg2UWCqqRgBS1Yo9bKT3ZMSY4vaSsVK4pGnbj1zt4rAtKzauAvc9N08wEgwJaSYK
wmZashYooPVWXgop8PomCB0XZ/N5dSVaxhD2UslpsGlPGS8YItE+U5l19gF2XG70xXkaErDGnKWy
ijqS2YFzHzjY1wAxqkkp8rSs+NUJRC5KK0eiZm1Swa6PrrtBOFtWRgjDVQiBt4STTKePxGdVa7q6
V1T7P5wy8ewRJgfySXpSIS/Divw9UUS5HgdrKe+RyULImskBcQVXcX2VrWH5v/kvA8T0r24VqClJ
IGbsVsO3t6IiY7QsrQv7qfmn2nRYYxwtBDP722qrU1vrGXTgzq57qRs9UCSsdKToPo45HJxKMi53
SxhL6gKXx3z9jVTAQQOo89CjjHQpHe3ks2WO/t0ch3M8syR8ZzUEO+vhEWgCAS/fhMilgpVx+cWm
sqVZiRnd1veQb0HlrbYXR2T7O8j1qevebzI85RhpUfWi5WKmxI/VNXOqXDRj7O/3UvvB1PfvSGyK
HmFGQbyouFrI6P9Z0f4hT4kTLp9J8AlP5AobH7FGPPCoe1fx6Xtd2i+hzyII9SCKhuucWNP+/UmT
eD32whOxQ4BN3JGFcjjXHbP8eoMVZKl6y3l+e1srbDI2UxBwJdRvSyWQ3KkW0M0Cpctnwd/NfYZi
bBNC4vPyVaw9mYqhp/0QRX3AqdjjyssGIllescQsUd99iW7OjioIom3xYmmV5Oka0YNx8S8guzX1
v9WM4LdhNWROlzc4UDViQo6/P+DzFyGCXk8z2yHWtLEfWQ+IDn7gXxrBLpDqSeKuv6EC498Fp3N5
IVDWAmd6E9nVKeLi/wvAxGZ8uEAo/LrUtER/ziErZNgKl4Kvee2kJsImjC9dYg46eb+504qFeMiu
KfeYZazfIPQ3P1UZXmbG+er0EaBnn1MJK5Ir18BJEmhNkcXe7mexvGiOAJc5IFU88LPGNUlc+e87
2XRiHxayrJM6XlUpdscxfAAxBocx8o8JhcZgnd6IKjlXvcTlLKNpsZVrmpEEn64jZIRx5bNwDyxw
czRqEIOOTPAiggS8Dyca8aWWeV/Gh2+YzWeWPZGJhSdgzO3CRPXy18iRyNpYqPh6L0vV+iLdgVDJ
QC3VAL9K8a7gh4k7Brs+WjGloiTDhvp4e7tIygqRA+Y8b3w+H88lU8g34QIO0VbQlnpHNIn6IAtY
MuC1qpaguawDj7/HzjyGt7E1Seci9Oii+f31llehaJbC4cTi2jIJPUZxxKDyNzBf3iIYlDrrw8/O
qkMzCe8tFqi6a0AMqPLA/fyBzlQbNn8ftD9O/ykZKRFLm9LOfDbhWxmesc3LAAVPH+Ajn3/Vfaux
nSwOeJEyysA1BZVGFkah+u3V8JK+cCN+B3/JaH+L511Rj6YlNMhdKBPFjvDU+KORr3eWLTYtFNLq
GWb6cbrC5m8cuqrtf0+BCM0MgL8PyTuhQeQ9e2YCSsNVnVvlf2YLhImN8c7qdn6ESX2WSGZijzDK
RIQd9/JObqhHvWRcXvWShE4sgylppKNirC/Q/rGVzvaJveqwJd4BZg3ayZ5hIsVxBpjvg5GJnYru
kXeXsDmz7s/Ig7Z+NJE04P5OBUFnK1GR+vLIjUNr7BV21k7L7gLTjeKz/uUdR3P/o6EQbcWhVzmY
95X4QAIPPU3rziN357c+PBBh5ng5/wg6tBE84ur17fDTI/gbaD4y8CDAEmmNjq6EdSMqIWVGRMTC
KH0wncDqaq0rzNtwzFck8TgBmfJzkBMSnznMAqg24kA9diWylAyfuRCDPrfuAItbryBu0QD1DPah
qne9BN355YqwTTPbhfzSLVLfNbtMD1P3CH6ep1q5lmA4yhTj+yxK8tDxGkEAI12vEHw1y/z8gASn
YHD1j55ElwFjxnmmFUIl5/SMmq9lbT4j9Iv9FCrCf5T469W3X7agqftxojJYgmtOnQNapHweMykH
Mr1GbEa4H6g6yJJnWLeFFsAeAXpUH8p6Qm+UfpmjQkC+TDbelCkDXywnIKYi0DWSY8oSfAWxgD3R
peu4ZwmBskzQbao17sjp2raaAZKaLiysbmJmrjvCX9WMFC+KM23YIUJ9CKR69s4elfxO8wkOUZwU
Ll70jaMlPU8rcKOcJ2LGlrYUa31K+oanNvIIg6PK4VAXP8S+xNsGFkAB2aOk0Hbm74CfKS4lRAQ2
fPapzPCyGy4ztWPZYhSQ8h4eubjqsX1oYEbZJixf4F2yGekS/1bcodDD7PVwigYCbR/5hSRbMuqe
t+T8cnpFPJYAB766ksj69p6U0VVUKn+xUHFxxmY72pi2qRGigURaLrl+/uz4eUHC4sxs/Rv82ZIh
hI/WrU3EmLDAuamgTO+17MSN3QP8doqfe4Ib6ilJaS8c8R8TKy0VoPUn/unV5vWY9k/ouhIFRQdx
k3aj9zi5vh7Kezpx78awmIupoHWf+gwyqUP6FYQU1IJ6QxG7znrb7eWxQrdf8eZs1Rh5Lkb4s4yP
kXFAbmibyvmR4UKspaKPtAqQyHMO3P3jdeyUND6TmiPsOYAmZ5GR5ZO8p4sNc2Pq3SuQ2cKQVDEm
1iShd3c69T0VwC5YT1Aj/laEmWPH3uwAd0tdOvP2L6GfjhEvgzUB2QUpvShNovsk1ypDIGZEpT1F
4+94d4ijfC+TXCHfvyrT7LQQNK+IGcqGZ8J1sHHRA8Qw296dKZKiywCLh2Oru6sZ+0bOM7RF4pC+
6G70AzYzTNQmH1ZJLVz3mNvjhy3k+ixi8I5KjOa4I/ef1dr8MuIk1Jy6yfxb5Nrzq2nrfdL5Ch5H
CXx03e0YWzHt/JkCWLOTfrIv4YSWeFXE2fY1Dt0hOr2QSq2YjydIk3RcKBF7uDv04na2+iE9Gwiu
4kWV4lNH2U/kXAlg91cNGGZ/GbHudQfcan7LK+0UX3U24r27xSXy+8tqe9a35h2yuptaNEH0m7rZ
Wwe5khW1rZR9MzdnSGdT7njdXm86IpuKK7leIlZqfFNqudnheNHusepGLA3chisyUZbDP1CvxM8U
5Nk8cfe4FQDqcFx3vEE1grxPDdlIMOsX8zJfurDGpEn15LJxV5a1p7oaENTiDBMLAqwsdcbPoLqt
WphEf1pDV99Qyde0iEnBsuF2tQeMMQGumVzzyUDvq+rWfVpQpz1mKmJ+DvcPrqBwAi+LVs1nnSix
Of0PpHCrquXnLFua5y4jp/wj6lise5cFNnP4XvrJfRC6XAxPYPGcYJzFr6SOJOBhct0WbiM5+8Wr
+RLfWB/9G+l2lpdaRkm2rEtZuSgWMmP0z2DDHx+ubeb8B7hbDlRaWXgmE7M0QWJsQXZspNiiqTrr
baf6v+eVzqamCaX62fb7AJ9Lgoli/y3erjGOPCifH6xDNUpB4Ep8g+iG6SC+Sy3Ifb8wm+o+ZCyU
AjneM8VdlImFokwDA9QuK98GTgaEx3DM0hx/05EF2bGiydhkQNIhUQD4hjCqUfxarjgDm/WsXWY3
5icbAEj3T3pgPuGVovvXLIpXqjaAx7FYGtkSNUawiiqTkXP3mr47SZYPRRUhFnYvadX+TxGg96sk
YNDHwoN9wlPBBhLJxYAzYYnXRNooYtawXPb8B6UV482bjVTvy8fns2ut0yKycqJ7Y0UoRs60m1/I
cDgd12ukkDaPI1LP7pZUVthTwo00drGpGrEHJXxZ2ff2gdAPQ90iW0Ion2lMNcmw4O8NXv/oGoxM
XU8yTgU3INQ+UJC6tBSQKmVK9DoliEziWla7atW8Jy/lV7yRCYJAWPNx1tu3wXQE2ppUz7Q5MoO/
HZggDTaKkFhHs+VIbgOr+otVTLzU7GIwBbeWZ0scLbqRy/WHgYYvEyN8lXoLwyDv4RFiTJz+64Bi
s2jSwUVOavjcy6stpLxMPXz1/1TLlo37WD/Bmu2NJ0qsYyG5e4+TYmCFXqWnabsu7sR1fntjaniD
o3XMTPIiYNBG/oakV/Aq6nvA1uZKAcFB2GDqYRRFAa20XfEPuL8wlDD1bOvML31ut/CFXhQvGbq8
WwReR9itJYDHfQBPOQoGz54qOmkaWBfYZQq7906O1RhCn9i9IPBLpZq4FfmMeBo7orIZKbuq3Mwg
zHm4OZ6G88Qrw7nliRpKZAReZYsJvK0sDHn3A2y6S4/vCqYvN1QNZS0mq6Lt4mOhY4ziIS/gFhF1
RuFgQeNXcYwrmMhj6ddoJ8Rj0I5+4xpVtJQ5eFQVaDI3rvSz8243PH5jpz09INQgSQ+2XdoQfID+
8DYd7uFmcEng1ELh0GV9S6Te8yusGxrEi0H90B+5HtmYXsHuVhwiOmigXkj7NTo0B4hjgx2GskTK
H1fxcKnjarrToOKdeQ2hxiJCv2mnRJWYSheo5XeLHkrQ2ZCgtFjKZhGV7F5ToOBuCk2KUUJp+v1C
zYWqOcMDdrzMoFcmQ4CXT0kw5f3pcWEA3oGO4a3JXECOHx4mLZcJSQd2btYhVQoD93+cUYEXnNPT
3liKTsD2ND5x1AfWQxRzv3ElQFzDcSRtqXnZ3+2wTILu/1nX8NJIdrxiuCmsl1otYIffiTrMBa7Q
tASFWlQVROw/7wUtB4T9N7ko6K/piB6yvWt714WCor9CoFxzvATkETPL3YhpPZ+7+CTxLW7r4bak
ltp5PhHGLX9clnZ80NbUJ4L4D4g7P/wAPLye35/BI29+MshWPvJ+zKz9OvlChox2++9fB78Ek1DN
fXDW4KN6tfhpRus06LgaF8oAL0hUguFBIXg2xHHEtcdB7s/DqL+JIXanhduu5OGUZOZhUHihXyLr
4WBNe6D5iVP+psbv/PDy8E7wjo2jATswSW3XZybFKKGltz2lfVnP+/q2mYkX5D84cUAnQSmSEtQ8
RmelhYyWiEVKzICiOXv9Iz69izbkRpDCXKsnTmewX3W96tWaFOJhl8Vy4j9Fm1lqSe0FcfjnJpxk
Sw07RtyyefNu4pMKfE+g+L3gUJPcitIM+VGUAV8Y5nK5rsdKP+HzDfawsnjLj2OPVYVaSftjsm3L
sZBAzmpPVZy3KmzCF9/9aByOaHhxa4QAAJF/ybMuMQJ4Ms78QEinU8F8wl9Qan05xF8YhkLtFcji
YYO+EIFLrIzgpCNj6E6mk37ALqLTTt2oV5E1LLUvejNwlDr5Oeh1/4XEQ1SVtfUUjPMLcssDcC+o
b7EuGgxzfqdlqKtiPR3OLb4p4Y9OyJ2oL4zLefStU4hisVG8LJvRWLqDkGKBpCFMF5i2WdQIpALC
lNfzxf7884EDEkn+iMI+BTKnWW4Bz3nIhjKWwZVHKzkMAXHpmcK6bk1EG80MTsmu5YSRuf3TP0Yq
HkGVce/pG/IeLgIrCoay3/zC4vs2jyc0iSg23ZKiYtU60gZExCUARUE/FtAH7dyoS81u6lprIewm
x77P2qykFyvSP2iLUPN+x2EjyTijVnmgj9SnPnUFxZcfzpu5lwZLZFIyMn8vmlqNlZ6A9m76FSJg
t9nEQHZARrLsI2E7Z7KWkgb74NOALSOasmfnR+kM2RiYp5A4baLbsSVo+t1LQfGPcuIdq8JMB+VO
Dq9yZ0NwQxVmGTgwG/LHJBokJu0ybAkxUTqnmNJoBkj52ABjq9GY/cIbtmYcny1VlrCl036bdFds
/b8EEBRwtvu6ywAXI4iOQMOI4owyQGdgktGAqhbzbXexZiSk6VKxFWJ+jNPWgfWSdRGCeGdNjRCP
hkPzcBI9QFdS91tfbu9bFEx6lRrmanDCIRpUlCJIgseNblejPfUyMziiw1jo83Q18U3VTx3CQnGd
BeEfzPYu4dpnmuCr06z3EhxRNaXUgzHhvNFbqagFyL8WBI+cyO+TqLSCYjdsvRdr38n09Hg1m9iy
dfZXhCSm5wXN6ey0CITDwncO6rP+HuVx9WYCaGZttiFtImxi3ab97mUbUHl2mGD3MXE1bEZgBKzG
IWT48YgQl4Sxcd+B2jZ+OOejzri4B7RqKrgLE6DH7KeQc1Bh1gsTxtXJQX5YHocuBKvK4Ze41/vz
NdnfWbCpS6ey9XmxNci/itZ+JEG0BZpklNctpCUiKeNYeZ3U7cE6+idj6wRePMPHXr0J/1KVeTJR
cKAmlyft+01m0g+zVjwLS6koWdqPsUb8atsD08RE7vjMrX1Lb+gi/1BEvU8XYMQm5aTPhAse8eB9
UlZBWDO2gxI95QQGakmqojAkUaIgae8dJlto3eRBzG895ZvMJnMryxIcrEgfDBZHYDULW0s0jQhq
nx51g0UJhs4bXCsOadFIiA6EqT46rqOzB9iLBb/w6fX4MwQExw00DYkHMNkEK2W5O66VzpkRs88A
hfFlAa5inlluXx02VKIh/mQdElGoxD+hZmS/e94ELWiKNY7dK+4V6T3I+qQqdNCYA4pmpGpp+juB
bPAyCPZfq4XDw9N7tQ78kVdXLJD2BI4L75MLal68GdsKfEpqmQYxIDHEq3uLaFfN7rS8YoDAcrua
Yc3SEYc4mr2QS26g35Wm1Ybky35S+DW4cbFvAzfzYk9U6HwXV/Yz61YDJJJDBcc2RzAkDFsgia/h
NLtNJCvMqj+MHepek8Jod6paoTbJCmPjwP3D34rYJzFkfwAPRWYi2LRejDF6JfA3MbxBIN9f6AdB
x+BwWWn5XF3yZc2MNtWrCcET8YMnQG5zX2ch4Ijb1Lg/W8sbZVjxwvj0xx36Xv4oFl5rdh9Wx6Dl
8EV9RtC70dIDLpSv6JUY2x9e69BCQZo5t+5vI4Q4EP/DbEv/ceAZKMCnW96xLnaTvRBmz9EDfAF8
+zmkUdQpcE2n3kFbtbUugvvvb5QfbKZZC2GAlFXOuLgZOeeWSs12Wwez64VRdWqX5gTzq/3GDSqB
HxHaaxwRBrXOI1r2ouK/ekmUwDSb+6fXFqa0GjWWzhOzlg/+BSdmXmo8U08XgVHeiuSUrFGgAi9r
O4HoMyseRnMCgRFWE9gGFnSdjNHDLhqdJXy8Y/szAPqmcYqg/jqw7VhJdAz7WLXjCoerPH+lRXaF
VAKIIY6VlM1ILTzUlOw+XKaI2UV9UTUKr32A0+b1tuIxG2RKu49V1WD9/FhkaCOLn6G2RtlLIsnh
MYf5ZY2QRkv92g5o7bCt2RkVnJctqDx9qaVhF7sctAzZYVfzf4/SusW0h8mwtIBuvI8ET43OrxWd
Eg5xbhCwXThRoPxehql8cmHvz3Vz2Qr3cRA9suVe8oGsS72U3KGpBp5NGVXLFA8Hvg6skua3HVdD
9YmeA9oH8DIDEb3pewicPu9jJfzAMyID6xKMWGWnQPQQl/xdNp8fXYi30/vjqJLiSwG0hCzfpqPZ
P5Hx81V08H4fx+XCL9iGWYCGUw/8cxwXzAYtmE/x/d7jbZEj6dXrOyQ4+k3xeJ0mFEecSBim/ii/
j+iF6QL0s5WSbj+h+qodBXHbyqYULONrbZH8v7AWc9s822J4gquEY6fyzaDlteS36mawjMW/AQHS
gUTnLihH6mQHKWSeg0Cxb4mCKmJir9CARYcffMssR83eOKgTIhVNYrHevkRSuB9I4gyQdaF1hMdY
JM7OtTkzeZInjj/OAmo+8Ns0BecQUSzywS/B9qfCgS9arYXdTaBHL4CpyY514Een8JpA1nN0LpWI
wRl9zTmIOaiUtwK7jwuFa41xVcqPQSEZ4EPg/I/JNE56JrRx6504/FXLj37+UFITt7HSgzpf20MP
NaafgQ5QLYeBJbrS1fSCLeTOq0lTlAmePYz3mloO55oFIf0o89RrsuMt6wMQboKUvzMYhQEn9k58
rL0QPFSncJQz4PjxzEtvFEUjOcvaCMLOQWERbiYkaUj6CZZm5QcLTQY8lCMPqozcfthOUfqEiJ8H
ApatVCWy52zJ+MdZhxIYdpVpNTOuw66eKFNfOKopblfm/Z8QzYSqDGsfQo5sn7a8ofes+Zvlxc2N
T+AUSy0E5JhghQ6UZtRZfnNPXE+y/O+UCYJJNlx9E6/lRRVtALXB6/znbBiFUt5aNVcGxKKMwqej
cuspYJYuW6ZaPv8t+snLnBPrcqUUr6SMvyIMHUdokDWKrKQC5tpGbpq6HyaYYMBI6v5XiLvMtmxd
ENqq1RZxxc5cnvrOL/D7D91pkk0CQlFBrHhEyZxE0d9+KWelUmBpQJkBUdu5mKj7vBt2je8LDj6Z
EC4/PmZPMXyt5wqpP8L0+nrEXXhrZfgSmlR4tvd7e5FjIiIaCgvNppqKH0P5d08S5+qGnxl1LhYR
yY8OQ4bAEOIl9L/4OPEGDyQf4cZEhDSVUKBIxIkodw9/9rIuehSNIVxzcr3waVTyWYNIg6kSppvL
c8+LaFkT2LG/5t+Kkx1XLaKdWozGD9a25JJK1Ive2lwgCV/Mvp06uixGMpIX5xmihwDfgqAnzZzR
tgqS7EoDimqATvK8dRFcXyw9L5O4zC9ryQpImhSMPG3zyWI10oURFRwMCaZfM5w9DYalg3FnWpVb
sgqA8RbjsVI3Qjzvy/Q6qBs8JjeMhUihPi13Y1nDnjfClaY/r17KI5CC0q+yu1c7x4L/b3TI4BaA
uxsKVcMpXgYV03Xar9mQ1I904RmujB9WdXUD09ziUHPKJv6dpsKnljySBLWqr/lAJAlgJdUIj4ys
U280LzIs1JkYWkONr7kAKYK+OstH3ny2AMObbulZyukwZ61YyAtOwqPyhg0ntAU7eTV5vJpGQMVR
JGohq4Dbrc8IUj9BuMUTB4V/UffqqJWfXn5TFnUOdCbHlKBoIY++LrsqESt4IAWttiBxsnKDY9AW
VevztsKuW7uw34ztzgtK8kCgvK7HSGnCw4+VO1V0lUrxg3C0RmCIndlWdlkzwjifs+RfM+Nzc7vI
9BkDn+110hQcSmQEHQr8+oEcrEF5/RgWqMwcMO4mRfQ4QmD8oeVN4Qq8kMDOEwQCxKX3UaSx539U
Q/haCOrINkpNihcFFb6dzQZGXvP6jPVnrQ5+844QyRnbXollyS5GzPBTLItjS0/qpJzcYkjQsNM1
rmpeoB/LtuJVOeKLI34V0dZWlqZmgc5i3gbMY03Dt2W+wDud2Eql9Ci7sH21FKRCp68wZpOrXS3u
uK6zypA7NHf5FQ9NHZ+iLco40UUQx9e9F5zoXMPhmuzL3AJOlZ21yNSvxCNCVDEZMcBs5y1twNGa
pzzPwadX9nYrK1YL3Uaby0hU81wzbpyz60X5vTfLoqMnKla2Hf1tHaJOGby4Jl/fHUi1lthnHAiN
I3aNvx8JmLNVY6FksKGB/DEjuCi83fCIVau40zH//Vv+W5oBFm9g0D7E7FdHMAijhrPDSsZN4cS3
PhlWl1hXDasz/jbFB4y0jcrqciqPKyknsj1jt+fj0u+Zdo+Mh7ahSXZf6494upmq+1QKBB83e6BI
o8uadbfZKhLP2/LYAcODs34pB2Yo81FlUAyf6h42c+qXN5kxd0XLfDuhIBCKChIvfgIPYNpVFozd
yrlxvmdcWw42tNKWfXL3cYGnC5zBxOcwWYPipox3uFCxcsRYSskh5lSLSEygdAIRLjYc9DXEiyci
zfAX9zyn5GLypDstiC8xzjem5l9K6srx0/rJySB575cHLqb5mNKPJIz/q0OfRqOi/yTgb3tLRgal
8LVUskCbLkunbJ+BHfpSaJ8mR071MQTNJPSr4G3moaoBy1rhcEpERjy6ZKTQCh8m+gRC35NjnVsZ
qdPhyaF2sgLYoCOIIAlkiw+vW9fWxr+lOzWuVfrrd7b6et4WlWtKeO0IZ1y3O8jpoS/3kfNnccae
NgZQTSCAAtKKb6c6fy8x/XbMwjOr5orH0NIJB1Mx22zFDX7m5s7W5kbu6FQsJIN2ggOAGvn90kz4
V6RJPPWGyI1m7txVpyfX965mBUe2la4ZT5FL2Mfb2Oc4cZ4RWVUCW+aPP+1TYhbjn+alnQvQrfMm
nPNqk9JWYl3Fyljz92JplOFTyt0Yy6k41E7UyghSZ9pjCFwi4xilgL72bZOtqRxE3GNnS0d/V4o5
2GuF90KQugmLHVzBnwDFFCHb4b4eCG+gMC5BGaLcdFVR/6KYNUN3ReMFGOQaipFCCObmZJ13Ck2E
Q3OwnLV11XTX87ptVMuQNsrV9GKtPPYmrUEgf3ZOJqE1y+PwHJWTvjeaoVVZIOyXHNHxqBuz9S28
efbRBa00kp3wGAzk9y4ovjkisp9m+2e6uICpoMMiu4o4yWQqSH9QtzbXRpz2GDPg1qwvS56EQs82
U7tY9LdaycrxUZYp8yc0Loih3ed0dO2xkWk94pAzX/bNYWpXKFo7p8oXfckM4j7urHZBuz3bl7BU
tQNMgmWPqfuIBgfok8lPm1UAvIbFW+x9RiadukW1iCgKvGlwj5QcW7YZeHn1maFsS9Z+SqMxLwhV
qTh5adVykeBV9X40LypJUjwGbS0SH7YzRZr0mVfGIJLjvY4sa0lZwheX4SR6S4d4Y8vB06R9jkPt
Ee0Tscplqeojib18wqZs5XX32AneLGgRY2Uiq0Hs40Oqwj4xcXCgWzwJL2R7k/WZQoIPgHPJnI+h
/dokXY8fagBxnJAwuAROKy7zA5KbJrSHEBgAgYAHUXUJxG0rYeC52+Y0vH4ymy/gV80RY2kQ2eau
CY+Ob17UaX32/6BYENWMUfJ9ZkgUZbs1zCW8GsKIkROvY+aNEyhzFHDd086T02sDQt8uqLIkqcTw
KzvB1RDevgxdr7/W6Q6WSzEU0siiDUlCwMSJ5r0TtKa2ikIFUSUcOEpiJf05yz2ac28y1W9eSuy3
BjVaVHMMrEoSPSYQJ0vrYty2ZPJ6dlLrByqbOHfPiT/wurnAYDunFInewCHSu5kmNwaF9JbhRar1
pwvYU+u6KcKfQ2pDg0X4PvW73Pwwij8q0NFrSNDbaqoi337mX1h3fTNkNL+/5yl4lgKp+2hQO033
5em41GWEqFilaCGbAevhYh+q64ldeApUleA86GFTbaQD304zmPa+xSmm/ZGnT2geASebTct9ktDJ
cIjXLTm/Za80l99VehqOMwNm4Qb9rjjwzJGQ1lo9TezMYvcZKNJLg+5z+kk5PYK9nN150lGy8IcV
a8N+iALLQsI/vmg8I/749LVcG5dOh6ENsZOF98GDqOC6sjeZfZn4djIZtIrTpNJO+1m4SqfNJ2RS
CV0Z4iC+S8HUtq2HZuVCqwopgDY4MUBnoGrjJai7yR24aAd3mk3HJvt02TeqIDjutNi7c8MfKiFe
OCrP0vk4BIEZyWfB1r7aQSTptUcjeSAlyYpHh3C2+wb/9oxF4nKakLryehePvL5zLKaKKMwrFGik
hH8GdWzBrxe2uYAU2RvULFyH6mb1F0khbjfBNOwfpnNen/vzgq3+eXxy051sZRt6i71SOLwJM/r/
DykYJC1+08vQM+5mu3VtSWBNTZ/wPAiYZS3YdXlZSvGv/zMX3BqZR7HBjN5UjGz9aVtvbxV60U2h
gyhHLPEXKHHDWWnQphk7RPlf2pUGpApmCQFeC1yx3J1MuVYgk2ySqO6Waqy9lMhhpRo2hWIgozt8
MZ0a6gUZoxsU1R++pBk4a7JJHNWZfKxzwmcyBfz0YkGukFqmX9stRNzh501HCsAUEuskR0kLjboM
pZFAMT19ASD72XWdNQyHCj0HV+/h8nTY1Uy+2d17dnRxcrc+sSSkzkARAMcsdVPf0OmiP2X/Grit
kKvIic4qHnYaZhtiR71OO9gCyyV3NwccrUYgPSsQXdVMHYC8YiY97DXMm7FXxdyKQIT2Mtj8iDYv
9dD1bekENRCjbccNPBdBZ1Cl6AGrMygICVUe3DbumtbGur0ia7ViUY2KJg5T+V6+jOlWqCTiQyIs
W0O7Hbd3Nu2qpJZzGlyvG8srlJAeitPrKB3fRFGALT4qEXlllkuQ9OwJKrRG2WZq9fh1ISVRAEXb
0/H2cvL3cbyYRPtSYtEbM/uwNsN7nvOBd1ffxtZ+nh3A3MlLdRoOnHYP4UkanC07MCZBuanaJiXo
JHmJxkegS/vqvoxbiK8dbVpH5TcGLhF/KucnFRPNbiwgntUmmmnp1RjQ8pw7bh8m7Co2RYD88ubj
kfaIVfvafahZc9lnwK4/WbPfQz9oee6KJxTmFAkB4WSuiNwiZc/JqCGtxZiTUq03nL1+sliQIKU7
3+8UZE+KcLnFLH8molCNcQZfClESv8uPe+hbk+OpcR6wQ1vBtK85lNA1PmeLalhpigbjg00jY5FD
KISAlbtIakEIjubFnzpjqH5VsuvJBBFh5IjYO4COqSFDpGD/FeIwuSprOop72YGVPit1zM9ITFgw
TAUu5l8GhmaSPx5CVcbmm2u2eC4VWkbD2H/TWgnZvD7VP1cF2qjuFGkcsXXXWl2ACvfoSxM67Qgr
BcpmxwmeddjjVdQsDjQJmZnAWysiwrAYUgUQANOc0jRE4PP4n5dgl02f+phQMKfMyjVj7zW2V2oS
RNumVyKcgJ0phxcKbgEJN+znFLx5XX1StPJy0v19yUQmmSLczxe/jlBmEFBFuQSXdkN3BMKScMQl
ghKcMWtyn4lcosR3TSURT4pOj6gD/R3TC96OmwmaVNwxdcUQlgkjIBlnrRNG7pbQBEF7z+E/wCcq
P8Gp2WQ5smj3W1DIXQN0IPdqsiqyHHgT1/u2YkLVzCTNBgL3gxGbHlrL6ZWc/qRddZYAWwzbiIXC
THfxXUbSzXxY3gHhKc1Hl4wt5dsMQMrjCmR0re3VdGTqUkvbt9u3M9Y+cycrfB0HtesPm4a3/JtE
yhVOiq7xzJmTRj3TVFI3GSIMFKMZvZ5voZLe/UCU2We/DUM42QxVzcu9zGoLD7N8cu+c409jgNlY
eEEH6a7o2zzOBm4MhL00FDZe8e4GwDVtNzNtkCp211HeMKdgHXpomQX7HUIyXBmPZ+S2KO9jSgl1
eg+6fBjxS1fGUE1BP2LZSuV+35x4DZGs77Ha5ebIxW40Q23fjT9J+uSppgHE9FKYPeFEzCNjv/9h
b23geWshT2fc55Ji4s6iIWC+KnDl4ZAeCojroB8PDPDVXDI/uafDQwv5MkqgV+ufpnAjB77xu4+K
epxJ1SHzoQ6hvb6NeNVvwNLhCN+g6a/R8TXhybDefliCMq4RQ7CVFja9Qd/i2Se4038Ha5GaWwEM
2BYZSsTRDMWy/HreUGP0WAqUjJFtinAy6/zwL9KJI8bDVTA+2qa2UP4L3H6CxD6Ez4KSLoHOavrj
QXK/yhs6Kq1iZYRQWZQiyXe6InkCE5iZYdaX7J266uZ6N3rmkpW3P4UmXCOiwjzHkl7hVivIDcWF
bEjH2djea5yg7FdmjS2CZC+NVr15WbjCAOAGCKIypeofMAydGeVy9K3i/A3kSMNyUxsLb/G4YTOS
X3xrDSkqgipWUgYbaqWrAKJ4n1eIhNjSblFD3JTWhgtEAfGv5UvmGvB/8G6dS+djl8BO1KJAcPxb
xQjR7Tzu6oKdpQzicgrJyut7k8eoC3a2FnSefoqbParFgbJaWFTE4tgWR/JXpDRZp0eXipm+PncC
oYa9zbf0XdP95ka7NG+8NfXABVop6qoIDjctABdDoVAqYUWZtrcRzxsup7piX+AjKlPVBrr19r4x
vnNibv+srpBvEmSwj5GpNdgsHr+oQaMnlGHG/K77VM6Y1W+dhGWLPpkvUKxoqHwHeCI1I9JcGFk7
/w00EcegfT8ul2vegutP7QOl349QNy6KwDnCvmv7taqaSSxQMTIgL4gFzlaf8puOhOx2SKxWvm4b
e5JBEQHhFB7H0Aah0gFu2Nk9rz8BjNu2jTeNTk1nM9XYtFpbEtzU/yxA+g8J4UnTvW49U2MN3lkI
TmA7OtJerOxgpS1+ncZ9BuldMyGeQaCOR1zqrPGwjYI4TEoW9Ko+O8i7z0c0bP2MrmFfH8y9Yq+N
H8+sA6risP/bIHTYlcA1Bhxyn7fK5y3foJqFJwpeCEDYU1JMxurKdz949rOBFo2KZ5yV6bT1wfZJ
VhIKbx+blZf4hY/ickTi6VeLk2I/2D0ErPGQ/Qj/K1p15J1DBy72hjMhJmbG/kB9i785FSCO4CR+
qO64zCuba5OOnzAfk4BXnpGOZMX+LFc3qO6ndu7UJPPuyr/X6BTFldJizuLb15F2rV4wJON5IVm8
UTO8ECIatU0eyW2GSxkC4aMwXRDBg8+YAemUXpYCg9CtgyXGGn3NPTlW1jwvkTl4Ip1cey34SvB/
xBCycicKlIPhun4/B9O0HIBUK5Uplnivi+6bTekOymYQyYT40mREDRdgAMey2n91ctwSYcvXfsvO
LWB2YxTRXD+ZWuFH13W7NBJquqDQEcR3F2IWyKEWPvDhYixJsgqEDXRpmn3l7QyDdOu3JK1AJ7z8
qoR37+fNDjY101lXC85Tb5Kuw+Pjym9xVpdaQxLtPnB1Txkui2PicTvV41mXU8VGDUBk/G3BIbsd
QUCA1SnDEW+NRIrBXFq8+pP/bflyjiiH6jMC/Y0YOSpNQjgK+bhIuEb5BIlzs2GB0bdgSY8FktCa
+KzDDn1hPoOummr4Vkc2erHIK67t6GHVCbFdKxwMnUt/8spyR3ink6gIVlKC0sElYA6h0tnseHZA
RcD82SZ0wl3BCgojgEUeSqUFeVmqVr+AsvtkWVfToqOmc2mHoydbtrMNlQ5XvaKNXhyCXaKAC7WJ
N1oLec7Grk8ojCu9eBb1TudPstnz7B3kwQuxy8FiVPokIa5Aa7lW8o5ysY5lo9gsDBMf4d8rTFPf
e6tzuMb4NC8yRfDEHrLr+Y2Dl2MoOkdcUlr7lp+99GA2wt5+gTm+3iDsCLjwnaQyerwGNvJMHvXl
C602iyH1gRv8Gi/5inCqu5V70AhfikdSnAWUjZszxc8fHSsPPbxsfPZgqUe3eDmJoiauLIbp3hRt
XyIQU3Q/y/OrzKV11AH/zrUHbUdRYenboYkdmZYsnHQ8rRcmaq6fJBtqJPBFRKtdeRV0hHLoBLIn
4ENEfmBkMyxV/mxaqhTmgCFrhULIUw/2pvoFa0bEQb+aEciMhasge8x/HURYdtiotsIPSyTSEz3r
ZH2iOyWtZ/vpHjqB8YQlZJleVElxM+eFajONE0pYP2LQSrhFx6YezY9td6+ER8YwUid/6XRz+Qpt
KbBsKL500tc+5gvFcVg9892tBn1i429uYoQBOUAW7mCzvbL2jHOMfO4W95x+qnQ/ePjXWNC3IuTQ
GsS8UNDS0vhMWCmmheRABzK08nxa5pN4k1mYEJN91Saca9lxYvdBi+dljvPkSagEll2b0/4vok6j
jxoUtMkNm/dKk1RAMNmA6N/7WkoyFX3CONjSUC8uDRFsm7C2WTWduux8fAC+rBuNhLPo7p+5GBT8
iffr9ZtaLygfBIkY0BVFKefpk2Kft15+Nvv9mpwnmJyCHLGvVpVOJqeKiQJ0Uyp4MoncrEQnyThO
IuEisUCH/Nr67MoZJdZFZxa6ZGQzYA2awGEj32VRXyLaM83aLnxf9Zp0/Z187Q30AIluCLBZo7up
5V+ZfgPmechfEQeSIk92Uwe7Gc2O5m9YtXyrdHlN++cIgxJ6ZlQ8RJJNhXhRYZQiclVgQowkQVC0
d6/J775/pobzmdjj3SXakAYtaOORFaxE4NwLZuGl64h+X+hJ0J2NnQ+iHArO1Y+3Zh6KRIL+DPZp
SO1hoSJV2kO83infyYmZB64myVMcH/rtT+YDrsZh3xZ2AS++oq+0Hv0iqA5Bf/GagtPI99AcfYsS
AyyatEpevB6ahMJP1J41YPo1Op6sGuSoYLBwkP8LzvNdjuD+EegMVrdnnIB/+Idkpo0l69GsoQSw
bR/nOLMtKYJ9MUzAQfbBlxFrZRyt0ny50bommUuDnbKXPi2tR7cSOuy8GykUe3+/Q0qPTBxjQWLW
QPK0vxyx/QXkSWPX+s3gXZ8+WsrqSciex/FIl6ZgHyjElChYbKZpQRlI7xBeBaoLkX5TCxz56uyP
RHKmQ+Jiqz3TMe+Blgvr98I7KRppoXoUlj/xc2JhP4agTdyxykooitAsPaWe1HPyh63SUcfcsGSJ
3hObZypNgrVDCijZEAlzmlyI59E8jjSUHg/jLOILkTF7/CDQIEuXKR0YqQbcn/z1OS5nzFA6GCZi
QGtR8iihvKZxUDCM5VyHlAv+RJUfMftYiNEdaFm10dYvOAb8lUzNKnwgDoxSVU2lcJYwfsWF1+uk
amgqkzCyCAjGXtYPIDsaBTeaLyrDsttMQy/pXW36/el6mFynQIFVSGxjZtlhTXvTgv5pubJ10VD4
J102XYTYUZBmjbEY8sdBBqknZ9J8g2D9AWzZ0pUfOvbcajdX9mhcQuBvClpvp0aZWnSI/mSJmA/c
6UdVpjFinhbfPlzL3uBw+2CEjQV2nb0FnR8JhH5aRVZkEtX/4aiMw6DLgHzN8lx2coVNElbkwD5k
ruS80UV4d/xAslOwKxjZOuLIzt+WE2ZqQqdkpUi1pbZ6kCT9RhfMpHbGl4dKJTf15IFcm1yQeghk
+QIEkHjN33N2sQY6hdF1h5EBr34L+7Z6Xo6YKj7Njhog8bNdNhT1Z1XU2MnLFTgzJOAhEIKnxfVD
Egj5U5eaCSwPceIc2zP50/pPjJnUk4dbqmFND9Svqw/jO9Rw9EqMC4EtqrZQfui76936KYMMjlFt
qgIgveHmPSN1gK44BFI0FTCx5rFcCPOJJ0aPF63vnB5LZ3ekkiHJgYNbOO5eNUrhdSOp0GgSKmc2
jaN+sjna60BETmF6XUTtRhXwctZXew48tPL1s9TLtxcRqXQ18inmli/eKawbELi+TFaxHChJZLxu
I7G6iLYsuPBOSsK5Hfsx5eVau83LwTakfejlN4X384G4/FTfJKvW1Bu4uj5s7Muqyri/uYgjpplv
JJGuiE2RQ6zWcXyqqRpLr/PMl76gJDEBwIc6xZcnY4GnWsMoipwoi1GSMDLQEJ2ILJOPeKlFAuSd
oiVWpM/haArG+cuXhAs1fc4+0ASaUqF/AlLbpxc12yTK4kWwuuNR1cRQa0KU4kSQBHPbKTCH0Nf0
o4P6Kjqp4ijvYO9BwbrBLAWyZQaqskGsrUwMJ1N04UWMTNNFnPERpz05QnR9juif+NJpPC9MKIuL
XOtADBOtaZGWwo2D8BmfiLtyCSmX4upa6yAe+b055hhZFLLQm+anTUfZbFrn6q/kkUDGOQoVlP4C
m/OJYtsJ9S6fNZoKUsb7CLyRny7EMkXzOXu0iipwqtv3vbBGIIbet69Xymj9iNH/g/M1D5FftUXv
QM7eikDIpPwTAGefJ5dpKQlNpHzP+Imyn9adEpcmczhwGrwHgz8M8Cg9lxxWLkcP4hG41AHq4gvr
au5prOPe8D+D1mj2cZ6SbfIYBS60VCaI7rIozUN0ccY7roNMj4xXXjaCWmVvxlyQ4yuLAxUOkHWH
iDCPzQ5MWrkEMmiMIH6azPP+T5hXgy8TXyq7eQ+5FrwmzlEFnnpJQ3jCPwN2Y15ihZDYKL5g8edD
a6JZqhkgkzgiTMrxpKPz/fiGVIg9niWiItaN6z2UxOT6rnPYlymbmZ3wwL6z0WgVZOsZO5KvD7P+
I2Y+V+HFw2JF9ac8c7RGkKbHolYwdyXJCyyIbt43zau+cuOJFqrJF957+goRt0VZ073c5S0OzkGb
BtTAd+OdVwjlP1Z+gU5hMJpSGDUMPHPlUUyTkajbZ/B6qfQD+KX+AQ4u/WKQkSQyyDQAimcXAtuu
e5okLuDLgxrOVV2D22fIT1hZAsc8g2hXtyZC7VVkX7jDIvuvwnh2RWSDbsuT3loJRCi7hb8c2Xsg
hwI+T8YQ2+pI0+0yToU6N77Az4KTI1j60P3AwywLCz7WCnldjVZMKw6xpdYkdEWMIk7S+37oypY/
4Q5eoNUyVBxmOBTbFv21wjl3A4PfAk4GgSjQ/RBru4atnM7aVu8VbVBGRkF5lExEtZ2xe86vlPhs
Jt8tsLda8Akm7Ny/YDN9O4vl/oCEbUuymRdK+ERcFdBfz+cH679kTnSzAX3SD1zXrexyMnd/z+Yw
YnS79ueTXM/5Dx3XmUQw6psXvbJWDZnv3M80Ae52JEU6zDntYAHmF3DVBN3SRUyYu+Bu0v82n6Ln
nCaHste+SdL/H9tIVEfsmslriIrWJqAkV/F0mD9uQWdY6t8wtzSGa851VsYTNqCNCqcTuo6I3k+A
6XSS3ZQImIdZYjug6Qp2JC1Hvce3TXg+YOn1sZrgm+WzoUMPYcGqQ/wZIkxPVW8QFBpwU9tut1CM
4WSNaGfuu/eamPRmR+wZTvncgKSs+SUoEJ/GMazgRWrCf0gJBqsuwgz8oYJHfHQVi729pMRGZGjX
d38GF5nVJ7O6gUk/nRHl5nPiebJZPlKlMvUf+y8jzdQQpiKsWcEjUa2WyOO2UHaA5s+tKG/jXlN6
B9JGkYg9lnvDFqMhZ9UJJoFQ7YZZXOMbi8Jw7F5sNEYBiY/+LXBF+dn+wa+4hsEpuoxz2HJd6Yb7
E3XehLYqI2hKFu0e8pGoP/qvmNXie0dAwM9tSp398QpfXWqAtQwnNK4fKtUSfEUZ3NksByCKwUqS
4IlLowzCEC6ZBWjLa68rCE3niTcylHAdRyXXtdUZUE89ylH6AZxXSSizctawyTjkcUzAYLGdC70N
HrHq8PmqmrZKdYsJLzlmPuwgc9hGYleuJzYQu8YGy4fAx+LNhE1P7Cx8uAdlIdQfJlKtpFTksWpl
OYsGOp2ZdzMmj3TbtCpdKJmHwQ5g7kHSEuS6xnNvlTaDrE9LAVvx3dvwS4v24mINYUZva+3LGaTQ
5GW3o7yxtWLj6YLWBJqIe7H5Otlsest/GIJJyVf33aWRe4G/A0/pZzSu92jLPm7bYx1EFR9JF2F5
vBglCh54CvS5F0Qs4MwVGXS8tMSkAa2GHdueN9d02nZp0Wcvs4VjUgdaVk+3ygJ0m+5G8W735SNA
5zvIWNvCX+i8HkCuLXaETJEHPdjtW+iaAK/WE9n07AseEG9PJgszo0MioIBaSQyk6ElIHAx4Tw83
k6PO3MUr/3qU5c5yJYJB6LkwBgiAGQNqp0OyCl6oXQixr/qF1tP5jWNUk53hhAY/u8/PQ07WD/UI
KT2Ey1zrSaF57VYqsNmjfh4A7Bpn4zGCJGlL434MVQJDmLmTuGWh5WAn7xugxLnmCifxVbhWCW3B
Q3L2DE9ng1wnbsSOTVYihDCoiZ6m8qNVaTSQJJMn+RRojQ/iUETDtl89vYVExIXxKRB+jA8SfaJZ
hfe1LWGJRtlMLAncQE8j8ht8ChPn/+aS3JjjDXm6RUQPDqwrRvXKymhDcaS/14ryTzPw2BpCV4jO
klYxJk22FH4fsHumVjGCn2VYMrl7lCVvVWMMxVRQoTKsPA74J5lxuKofMvP/vIdWpfAiS9Dxnl+S
MI9NOU25O1d2BrlYgVOGeDRosEs/WF61Wlc9UToAdbyzNxGq3MHCkP+mnSMgmH1kNb1m8ciW7kuh
p4bjIKkrqhQeIUpvvG4u2t8aG/TX+uO0MCfchO2MugWCaOkfxjtDaEnGUWRDbONpBdQOd2rDQ/lv
JJCNtlS4zafAxGS+ddGJaEZ9I5bBVGMtSbM/llr6+U2nMN1DnUYgLmfgFFmqteoRwtLGb2aBIu1H
UWFRRWH5MguMee/2IJ2JnRqakQ6YlnEbcLCLAzuljFkb9y5vlDX0VsQpXkTZhh4M2PFpnJWdlyRV
gfZUUmZi0cG3S4ExBXoNxgNrXKgxOwMtYRnxNzhfKvMme76pHZzQ7JQj6a1OK2uWUbnwk+HSf6HT
LOmbE7aK09YsbX3pkAtNNR/nTjkE8kC04X3ozxwySUV/EJd1/4cnz8ybjFjdZ7w75Nys0sOigN9y
TcMTuIASGE6b3G53qsQ1YAncH0cnpUwGqsFs9enY2DGUlWVcTqLpeo61InhB/9x7+GPBF78IeZb6
LmtJkAVmN8Kc8opUaCdU/oYj+uWeiNPV1089RuKiTSyvBBiscXGl3Lqdoyfc6qPxSfXRJd6R7dN7
osoV3MCX1/gI4zy2T5fTfVYQlVi9jdkcU8yf41Rr1GtqhkxO5GW1m0fq9JrbV4pequ97JE5IQ7CA
LDYgak7xBDGlorFjWBLsOBp5N6jFtXUJz5+8sOIfL8c5iEAMfLyBF9T6Od5fToHZuXtX+Svhbkbn
/ifdC8xHvzniM5DVoPMC9y4MuPmbYn16h/CM2S/NlAvh7Ch4z559WZ6A8hYn/mcvasw8+QbNMTiw
MvIV7lBaZXiTucj5G6sGRjiOgAQ4BVxkYUxoH4C7YrdWgnwq/dPpfptQbFjsSaoQOkH9JDAsh8fp
aZE1zdUwncj2TqTloDDIW3IYWhKSqecY7cv76JN63jUhevihi6JvNib6lUeOengPd7+oBSCtB9P9
iX1jTrmqNEF6PPspPhV5xXVO1+dRphXO60hyO80sKeSIThDqgfC6wtoZlKAXLAQ9md1J15eSdEyF
85HDFCdzqVIZVi8V8ceDVzfpyvQ7FmS5A69kJ8bhTDM8ftf+znuF+HeSVZnM6Ux+ONwee7AKxHYP
zToOPMA+rLYCJzCXBEiEPbhGNZfHfYyF/1kJCb1iHGtVmHsQINyyzWkZl58hN/ERzOVgPmO7zSp2
WUN0dSjP8H+epgdbsyg/ByjNPryHqZ0wJjM3MRfBra3Y4cm3cKjRpVbJgaG3dNoy+mCJ1v5hEgls
7X84U2tHc83lz3JFETVCW1r+S8f6A39VDKhZqR4tpdjohXsQXffjNT5V1FHROi78COba3aJVYJLS
XnC+xfMc4LDBsfcVzvh8/ImcCDmddRDsAJOKJHMebX49jylLyhhw0GJ0hrSJ54eLQaLOFGMntpM8
anjsOwPNhfTR6X987ViDidXLwrF1KmG+JP3XRtcC/uVazVE/Bn0TSJfJ2A0cB91RjVpQvn+LKjZW
fvBLtLY/DkDxjsiJNvIs7jEDQ7umkp0L2uAqPxCIlyDA8SzXo2ZxaJgw6iqJrU50NYy7IPL91fER
rHLpc47EWt8/OLogba6ROtCo5RLWb4cGIUrdwKqUtuMavY3+TDS3iDlP82FAxKLVS+GeXngoOBqo
vd1RA0xSUB50VESTV3n0lLsq9yP5z+ryXDXPsg6Fuv5OdXkAxzMzzkpKkSKOLqqq7jAaf/iuOVCT
Aa+hGM7ZtIpm6HT+k1bAApCzQ7UxTRdrCOqhUUWbbp1nADk4S9xA0J2A+BshKaNNr7icFtOttXdh
FnXih5ETUOu9oQVsY39CrchWJyRlUBoYPrFQK2S7ANK4NHYI6yek0auU6PA37tb+xaLaqVKEfZsI
aa+YZ+0ZZaUe6TYXDyhwOT93hKX+2Y1RamNCARVMRMNysQxJ4/OWEQmCCTRzCnzqgV+GDbBVMKQl
tHgZJ92C/mbfrVNhdSzy6btWxKKGwPcdfsINWlSwb48kHD+U+xARy3aMI2wSJFhxDWr8Votb1Avv
t0yz/wXZ42hP0IdfVxXfIgg+++DzU0mMGgIyfbzqeY8RfzfWMRE5xia8EoUJ+D7MaSyaZAbVQrvx
fkA6BylqDvPgJ6ajvfSBtfBIznHy2VjS6IRhnq01jhb4NslUIe1aLo+PmE2V6i2HZPHBuA/z3ppY
6utZZrtnGizVP19zUJDT7pJitaAwJYC/APqLKN6nJJzKaqE5L/XzU7IhkEiw3urz89f9WyoxaTkG
JrPDsyy9ixjOjl9Tdt4sdrWFEaIjFAMI128Hr96R1BK0L1VidP38MfbUX+X1ztoYYjvmvAboHRtf
W3l/Lp++dEysJAX11iJZdAZ4XaZhX+z2DI2B3awCuluL0Da+KYWeLF7MbLf1Ef9cqjWGdB5f0jLI
HoU8mFvO1cPht2uYaNMWgM/Mx+8lrEqdWBo7fPz0DB5of/wT1ysR4v6J0RvinM+UO0exxVcr25C5
a9MiHXbEquPdOLCJ7BXEjeNd3z98SzfzZljXn1NFR/HxdH6lZ4bWJpYvLmpRoslinnW1yuXcPOts
tMZCof0dP/4ubj/tFFMblbzb3VoMu67dOg7y89/i06eEM0ccH+Z8P2lA7ZINK6LObO5+qdzTN/aO
F90CdNOEfTFal0e5/ppm5PfHZUkt5sSRJXHEUrlooPoHhZIhPYXxFR+/NkMnAJFzB2M5jaS0EVy1
aOP9CyZyaube3fQ42yd86LhKrZb/1sIlwmF8lI/d9rribEbbn5Azg8ZaqfAAmDbULHPcZ2Hx00Zo
94vjKTuoipcpdDApa3k3nkpTnOiMteGyyYqeFfZbLLNUvLUODNB0qC8abeuXsFpGbt31oAT8PuQe
Y1IVOTaBQL+SRMrtMwpIsJXB47uop3m1gv0EIEGwIJDRza0S3BLavKzPlbrbBoqR4Vx43xGwsUQU
gGRx2nrpEvccKzxgBh8LUIZb93+STAJuy6qMUhUaxGCgB0QnFNBT/N2riYrhxLVLuvsRcEh2LMIS
KsgP7ROVsn6PKPnIjRHsQGCJMLYbC7b6yV+V5JDz2I+Jz6Vuk2C+r46ZA71Kh7C4TWt8+dvw610G
0P8zIv8XM1VPW1gdeJwVLNKL8EyiZ2284aVk667R+tJJ1w4cnZVwuMcdn2k3YHnO6ZTQPcfe8jiM
x5NzQAOu8VV5e7ab5mcPOWoozTV2emyiBOaqQW/DFiUhKb6v/00TnEi7PrFPeWC3ivQDSv5pwr8d
55T1B1s2X3OQaoUDywJoVOZ47sRxj1EBWgqoJorBfZw4pw81KhQFurB+6hTioI7a2UyOlk0VS+l4
rD/NG1RByAtlNOQn4Yz/PCandu3OKxcOte54/H7fedpPrFAoXOWFQcKL169ouMPfA9jS+C/yJIiN
EzkzL+EGj8OudzFlludVoqVa9/daLuZ9pz4xz+45RJjNRI8pUVYtnulAglF2ZdEhFGxcMjdA6XZh
CaSm6+ef6Y9cw3+qJUONuH+zmNh0LoHZtQZxB6RU+hhF4wLzmWPEWcoNHZrfqIXkb6vFSTfOhWnX
yjYgrytKXPqZpTVL/HCwDmgtiDY+CUXSxjkOpfONCLdzYvdK9JNS7dDTA56De3652/WF1Y6V2GdC
KgFiWJvSDDK9UwW8o3kr/JlkqFvcrJC3dFG77cT7W846YPeOQ8h/OHJNmO0GF/GMO7dLGNd40JAJ
XQkbZ2kuglEdZPSVVoYZ0yK0NpfapPwJm2Kkr4kRMsjgi5KLnp7GXPHdHywd8xL0BX7R6KcFwy17
sCDlSnsuU9ZUl5QvvBdNMFNh95USuNVC407fAYWOiP3gxlF2DH1toSd6HhdVqiuAKk+gjzD84gV5
EfOXhyEVg8Uhuy8N27Znhe/t1SkKod/tUwDfJ1zs8/Mf/MRjMB4zIVyh1ZfWVWpr42WQ6n1xCybF
ANIC2F5znw76/RzLnHMnz5QY/tSI32ZqzTo6NM9qQdmCftKD15MK+UzBxB6uoSh24+PCuptLzjhT
PPNXW07CicgT7/r9paKnj0N0dXWpWkPHn/TYLG3ECCrDNZaiIjdLZwTWFbHHZQyZa8J7QSlglq8J
B1beV0Avv4nD5jFMAmidM03kynno7RG6fPkBQBAuIKhjvyP8aoBCjRhvoivq7HHj6wwreUhNZRqR
vUi5eUqjkaXJszmGFuBlK/KfoSYsUaIEUUl9pXpHgll+FV1zZEdFEY1xuiym6sWqq86r7m2XUdrP
cbVfgc5iPf18jDI6FTIGDh+jhExSfSbzjaritQlKW5zvn3tV86HzIFs5NhnK0s5QDNg+JBbnDJmo
todzGPFJyknKdAa6m5nj4te1l+k5Zr48nkoaEMeMDD9O6FTYiAc/TLmQBjDguykze7rPhYfpQThG
a9kydPtiT/kv3jQjHsraYjgB526aCJ2kJYSI8YEjSWT6C6c6nhSX+JlfMF0GtWnUZQ2BU2favPWC
8gjcKq1RlYmtZrcXbyzBFqFrVL+lRE+WzcgtLVW14VWe3583/JV4/6Oa+v86d7BPdfYO+GIu9R4r
qiw9pCWpUkC1ADEtbt7zuM9Tzh4kCh+nWNPhAgLS608c2xfYj/bNM9/NCQtNvXWQDMNHfPht+sTg
iw3NXCSREHFiSVhRware4ze5yVtpZ6jb7K3HQ1tVkN9EOYmKC0TowHdrTGrV01891Cz05dtInozh
DW1coZumLChPFAb/xFrCXZH9bY92BnT2YRW9kMY3Sq4tjDEqlhYKFEv3IpvrNhoHCcj0W3desKji
7O86gRHOwvlwV18j/DMbtJO7hNrRDR24LB061AsoNKpoYVNbSp55EopPpq7kgdC7MwxNn+TVVC+K
jy0uUvRIGpwIgO/vLZgP99i5V70Jx49fYAcaca0qClFqv6lOFoNZ3TBegv//5RCSdzMj4EMXODAo
qycTZgyEixnsX9RaQoVwODMAWaQFlWzHN1XyGQZMN0Hw6mh1caB7dAEgOz0ksqjF0jkGqenUu/5G
aJVJMxyl4y30MRWWX51ClPG81YVDbjLjAc7dvK5hMOUg817p2i7DltWBZaYJIrmwNFkrD0HofNTJ
vEzI/oGAjjF5bOsH+Wl6YsSYv8jWJYjDM4hP86JsOvKV0yVT+ASGF5ESEn2M5FZQuuPbbOBkpSdr
5GmsSDZZM7KfA3WtThmxoi4NtrZJatqr5/W8qPcCpG9KTDfcQuICJDLpaE+8vHLZV5LMkktP1VXn
aul6CKYs/7FHXIGy61fA4X97hXVqlJ0/L9JblRk33EL836Ar1FcaQp3hpeTPA0sXOw9OI+f9sYur
A0Nx8+jfFSRc5H00es5bKByUJFBrMrIFsxBxlbllKYSXdLZdSDnakrzJW6t2fJThrZESGrWyuSW5
/Yt1bIAm8HzY8v/8Y+zvoaPAvZEotIfWW4kMpu1NXfP1EdOQd5emmINe8ADurLZnpTtNFcSK8S8M
Woa+e+zVSR79XNRgC2xhV6uclrIizXR4LTBICiGZXhlYu+F3bKmbonRy1Q9GEgMkA2sl+l44EErY
FqYYpq6uDUoWMxy24BvftkvlusiTIspA5dmYK7SUJ7u42sVsw15MOtNmLt9g8KlyzurY9lOWb3Px
fyR4x8SLhlxOuJ7wsVjWK2F9UBEnmx5pMyf8mlqdJxQ/eoulBlKWG3gQwmkXOUa0vvng0pudm5pd
2T/RBfXmY8ZnUJX5DkSga6W8Gte7HjGFLb0moDORPTNduu5Xi+PAGnb0AvVBPKLbPzWohPKgM/CO
mo75yeyDP1q4TopmSoKnvJ9YVKAAoi7NppOUfvCy/fpfbQOUAL7A0LP1P4u2lrRrLOQeuFXs9a5K
ht03DGubipioFTE/Fr+4KVrJqz6GpO3ulhaViYxB+nDni0XbTkUIywEaZ6Ren9GWEw5xEtILNDSS
FomzQ0YlviqpidMblq25LySYZ/Irsy1ZxjTITWibmzHJ54NAk+JKzQH9940kVrxthQU+hQazSOVs
z0WE/xz7eQTRILiV1DhKdRAWJ2SzjhSTGimDS6hAONTFgWtzBTxaNil/U+8crsEZLH/cKNlDlhZA
U2TrNCMXDi+nZgcGfDOfdHM2Ex/n1bq2IQVKb1UjypXvr0ifNiLBf4EeB6k3f5gNAQUrQ1ufrd5j
QoTCLEIwseguGL3A5KBA1V9fwDp1D4P39ipuqVQO+UeTxelYp43tAviXtpoeS4g1shRxZmf2BVvS
bwbW65aTjrADqGT/rQ59Qcnmg2m3oAKfYqCH8YFoTB9Fc6mLR/r+V/w8lT9CDgSZ3WP+28GoALIB
pSRas3t0CqYPyRsafqf9nd5FogUEJviV0FLd5eYUzT4KuCA/XbKoPf+GcWpJQkRwxnRo5vsxiGTM
SzdrMr8/CZI0dm37o4gqEC0lfuIb5vTEsDCwpb8Qb01C2Kn3WEcABMfYUZdH3oHhtvTZEwnZGoGv
JqkbNaB4nLFP5A7xhPWgFSGxPlmOiiB1PR+b89DsFt6feiruos/Ysp9ODpZBRQ+Q3dDrSX6Kx8zF
sM7b3sXiBGVjLHshkAb9tmk6fixQWlP0v4kb05GiG/V8juyeR/YHZUm3X/iv2SYNgJkpPKvkooc3
ieECRQ8WKwbjpApLoXvJru8S1uXkcvn4t3uAaQuI/77IQFlabJsGtuk5Ep8G4BpBEqEYwqYn3d4G
6mdKvFqcYb/MfwD5rjv61dP/T370VvYpTpV9Slw8nOVLGdjqvgEv7hTPxR2mV5gFyNy77qG59FE2
MjECcLM1H94PPaComMtOTKGIIAD5yUumADsap8OtR+opaK3mUGsN3sdRlDU/0/QhzkQxfZ8tsmWL
0Y/kgNj1eBTxC9dso+ru9tBOYs2a+KnDt1iqts6nDoLhMo5rP+fGheAsUf1oh1dJAiIX9eyyVu9a
cVu3nwUPF7OTH43yrNAG9z6IW4M19XKwt+mbdcABRx6qAiMAdRNKYT68/WtdZ0vsSNiDJd9wa90D
Hzclz+o26feWtWaU2bdQp2J6j718ndohHze/LKbRtiFzdbWqxPBLD9/DA2ODBcOhdz16iNOx7mAI
02CujC74G53aIrI5lLb7TunLzql/Z20PzOdvDOQKQ/MGg2X4aAOF39vSrXU2zblsJcNgD2BTG8jM
XqXU/qFvDma30QjqZvBVy6lcTKxgrxwKTUocJmdCnzU6sgS0MAZBeVSbb46y7njXBEO6Tn+AKnXf
kMuWm7Q2k1TjpL9ZaE2gfJBicuQTs3SN7J87kc3vMEd4CVXa4ZEJJMrkko8ZJgAi8A4QPUiUQs4L
5OnkezIJrXFBc6b/64k5b1IVuRiN35tbav191nd0h7YE9aGlfPvYqloiv5pmUp5QNqc38N18s4Un
qFTrkth6Vl/fem0GYN+je21Eb69Et3n9adnaArBzCQjNwJk6EoiWxuZNm4eYRuvB/JDC98she0bN
Hupz/pGNc2oxYZTTIAZxdRsXsWtTxLC7+mbnETsOrXnfTH2xAXhAGwWhR1HZ6OHXOtlAGSqCEWQV
7FdAIb/CvxTJTOuE24MkMMkglFcwqvdP4oHSJ6aAEA6f6BAmpP1Lxsx9kbBSflsYvW4bluAABIj1
HGzKUtsSSDP0xozaxCRWPX7fz0mNMi3XRcbH6A0n/R6/RzaOTC/7oIdRqWv84jEE6K7jgnAUkxwA
D2b9PHPzThM6WRfaHuEcXGk5ss8riYsSeDkZBzgUWKfaP86nRT4jyN0xvS99tIQZu5ZUK6tNVmXP
YPybN8T3yNBgNAbUAZTMz9hWnMd6MjxXNAFLQ3HrwfbmqwEJIFaOXWrye5BrvA5Ua3rp56QajR3S
Vmyk4uMSDILZza6obsdWzllrsMhqwK1mr4vKOCmIve/yqkpoI5qzE9iF5WtBIdWGN40gzQZ2dOw8
JSRGn35qyO8uqmdfhy/QXgicY1FcFJEe+5cFWYyI5pEvjqTWFOVOj2GcSQZglewr8BIRjIUQSLUr
OqZIGnKuF/709AKyrGYClBcYyhSfupvBInSKH9a5ws1zZQVspid9I9oswE/jEvyZujrcguGVGn0c
kUBOXYRtDZZ7ciTkvRLRXUKTrq2yPFN+83aleWYiwtLttITB+MdI17lxHohQODbJr1kIkWtR5NJD
i4IgNd34VaDmZyF7BYBL/HrGikFiS33X8N+Z79ZuXMUwGwHNoNuE8HHpdefgf/Qbvgzgf0hrxrxZ
EPDsTe4wRlu1unbuq5yK+B6NNQ76/9R9Jv6rXfDUrZ1RrrzxSlUltqk/FG+WsH8Ut84aWddUg5RJ
7xRPBOhzN7vGE5Y0mYpeVpNmuuYZNOMFbCegY5zPJVyg6OOJd4E49d3ZWHjUPSOlVmtR6mxv1wRC
3/qnOzkwb94gAEMdCvKkgEAFRxSFbSsILxfA/57s9G5u73I6gS1QqejFBVJMTKrVC194aB00jgOl
MjfT80RQdgwpk38i/CoEioZuGVjYZD0V7//gspXkGG+D6nuqvagiEgu04Zx2Fhp/1JGUea1dHvRl
aDgzH1GUNEKiIr0FEwcFg1/4CmJvFB5QeCb4ZLHG+ksrq17G7BUxZILAmhZckgNm42Yng4PnW7m5
2BN/YDpg2KlVM5hlfS0sfuFvVuilZqyruLWL8rgdiJXchJwKFIzlDFmM1v9KUxqCQkHDseAKKM5q
1LEw1C4D+KCogZspr9PMEU04aliv/Clx3IAkLB8MlqknMgfHPBxJGo46x5VfUeBP9MVvZjhr/M1G
AZPGOJryap8RtTd7mZmEOpbGPfkmAhs6IW8uroJpG42dVXQZBDbuUbx1tO3uBvCqqMUsgeAicXG/
QmFk2G+1ATDQHb541fMMFY2t2DusQks2xw36mkkPsubWVueueagDbE0s75D1EYGiqeFKujjRqX6L
BdEcGIpkA2SXZWza4sCyWAWrLGjSwqPGO53rM6wJrlLBzS1PCQ7yStpUfc6LE4aMHesdu//bbRHh
GT06gcuUu2RoTZfLLPkjoUYa+fRtXlXLU9a0PX4ft0wRxPcb6mhFiSZDEUos103mXiT1siC5GbnK
Dm3UVyKCWWViuWq00m4Vei+RNvYJgMW+f+x7eZKY8IgjCuPDjOi4xKtK44ZTwkTzTunp0figTfW8
liTTqFm1yZJ8EfJSzBLfmuJGN+z2dY7EcoHu0UqMfFlDroSeiGQrnMpNChKwZswmEponocw4flE4
WB37h+WAziQyn5t2Y/UVbPBREtUF4sD43o6ePGnaxDVmb4MOoPZchmDUVz49vs0b8DQCmNLHq0CE
Di1iZCQb+DRvpJyRPI1GlQ3AnvnEkXzxjPWUaeMPl0Ht6EdRk6ekw17D1tCEt3MF90OreAKxf0ic
jouA3fMjG7+Ekscgg2epAas202YniADlW+WPsnSj4aknADwa1ooimZ2tlV4MeAz2e2dfd0uQxV4i
3xMmxwRpKiLstPHYs2RYdrk/s4ERBRqfVyov1Tj3AVV/lest10YuNO0Su2siZg6YT6L8U507Qqfa
oWWF3MrcIi1/CEf4Pdjq5LI7DuzPJ2p2ogFwOyALolAFJD2Zl+zTXdNSQBsrFHzhIhUT3LWW+NTk
vMOCxFhG0oJrkBnGMAHGvwIbSMQtG+NeCguglaRnYea+nvtGb0yUhWrU7qJstYL7/BWfW1CcWXPd
5XAziOIge1WfFKjqsfOjASlRWqLwLdjUBLJN3AyjvG8Y7SiXPAhpPlzYBw70RNtumldQDgoOO5SO
nkfELDdpO/gxChzu0CGMiJtHXFvvzMz7WqMgYDj2wdWuq9gEdT2t6mQQ6+GOsy3jRHE7gcRHIJwg
pTxjNKJLez4IkDAHfwwbzeXKjZFZ2DSUoewZCrl7gOiqrUZWWvEbIH9PfWvH9bVR8Oob8bs0fdHG
4P+LJok5DHc9bX9dNs4mzPVXeknZg2vm4bVtQxC7UfEzAh7+5XncmlB/nWilIDbBo9VzAkn4+rrs
mlGSM7O3uSVUjxuNjhKGtdy26UbIt6THiBo3oAJP0jSNKy4cBGXnEy425m1PIeJZonXuPhd3jZMk
VUhPXJ61KUjOda65a5KjqdQgLa3kbJud7XXjkfWNAF826Qjmd3H9fqJGmUwF6Rvd0/vqRHg28/Ue
N7ZHExYGzBm8bWsvbJfs1RZ3cyxzUUfPxnam1OhAyMBBssBOuhe+YWPtHmZsAW5J10VpEooVss9x
dySNb5RF4JaPbivFfcW7G7DfQmAjwGXD35JIKGCB+d1JhetvWonA/n3toZX0VAxei/S41FYbYmu9
esicrBDDARnwleUrRDq1fAm5bD8/jiXjTXWbnY2pVWIw2ir3iq9m5DDXMUUwWJjRjQmRnZeG/5Wx
ioKjWZ5C/bhxABBGtF1asutCuAO2wgVgTJSrgDrzGMs+qegw8HVvM/yzC5wzJjt4Hrm947vd6gnR
LoWjC+4TmrphkOTmSzcNYItNH5UGrSu3Iy3ybRAy98pztbr84Dekobjh18BNafvfxnRarekV8WyH
tbNnI6pRn5AFp+ZRTtlVlijl3kw/AcuxyUB0lGhUwykCYRm0k2OD5PfDyzqV59kc52tAlcELRALb
/s0N/EibudIbHq/I1TPXFia/ZixcMzKl22L6OK749KvUfkJoPdTX5YxKXsBy+XGtK5/fMuaSsRc9
oqRseHsyyN6GZGWxlFg4KKmDQVFkDtH8/W9WPN0iYqiGgQg0dZrXn5H5g61xa7/+WVDufm+6IfiW
gcyvxAQoGMmdimkfREmSDoeLWWLY/XFdk4cOgUIaMmfR5D34ezKQJFjFN6Pdunryy5ItAH7Kf1do
yZCfx37jeK9A9nEIqLEmv+t7aJSG0ewbGHX3MHaxRMJIM6K1GN5G7uQajomlTWp5KdHHzNhR4tuE
0vN4rRJhfS1Ay/1/yOWxOh6M+qMWKGjhvJRe0V897niqP50tB+F8XcjmB8jrQxydK90Qt31od1NA
QDkU2dGCt+xYPE5kUEyyC1DUYapKUS/GUN/73lSHY/MSAeghUgok79G622CZYiacUaTky9PC+ztc
RCU3xqcc7fBbQ+kIE+E7ao9TiaHzbuXZCSZ2MJ7mnTAYZSm1A+Zrahx98Q6af6OEn5h6gzMIMcJX
JCh2OVDUvKNV8EmtezHu+vLuR5f106by+wpdIIbn99wpfwVnzT9pviqeJPtesBHBE734qrlqzdbA
W9fRA/vsu1srOq/a3cgrnwKUzu9rOVlMRX4Sl9jZiPUXQ7Anl8eIZkjlQbPfNZQyvE0IKe++Sw9x
uVRbHq1zSS9Q3gR5Ucpczha5NS6V4bSHS8AloxqpLHQF/hT5ZwQJlKMtfN3BMvvDpwKUrwE7YYCt
nViMOQp/Hkl3QVh7wZx7V7Lw5F9zAU9vL6jXJIArWdaQUYyJGewnDgi5Aa0ByJcQpPPv0j4Ajeb8
i+SOrJDP/UJnzUDNYDr77fv3grvVOoBODlBwxAExesoMToYVQjFNicw/YzKr7TgpX1m9hgXHIjVx
ezBotBW6hUTFOppsQtm6RDlTyFG/4fdY/8lt2RqXwSUdEFgzhPXSTYoPenY3Bq48tiMf2L2Vbi4S
yGcUw+YFeHStqIw9MBMYyeBwGPJyVnXMDWHwNQUZA++fWJvahe19CvMJzhgGu7IBn0dXFjtiBAY/
JcUZ/ZT755z/t4510YnY4ZHSBujbKY3YcJHw+oMcDxeKgs1ATmOAidJy3g6eJizjbIt2KEhK7yML
rgNh2hw5MacU7/CpiO22CzC0G0vFgniVy4XkLNv2U9trQmy9gdc10mPJelM3sNZQb6IU1dfspeZe
Rc4tYzx6pmR8POuh3mQdRzjY9LkH8EUo8HU+CsPhUxmtcoveOziD3VIjE7pdvVSkVx80FeeH6A6t
5rfVz8j9A+WSldCLtsWY0mVBQ8dliW1tDCxqZzRm5LBgjVEsylXMtRISYVubzvJGNNNZVhsgwx9S
UCoYeGeV8p35TKe0hL9yvWzOnR972eYrPvTFT9Sj8bXth5+1CbYR7xyjpq1SJv1hxxewkad50aID
19YkbQ59DoTsCisWAn/1TE4zZgh+v6+jsj86zhzPf9I/ZFD+AsqCY3OfV6VXi4BLPFEmjXBxfPRK
KT/E0yW4Q3MbtLwkenwjMRMJzVsgwlOaksRCXJVUY4KJ8ef7aEMazJoEqKjYqhv2t+rKTlghgIn2
c+EkPAYjfygHeJP638b+UIpJhvJwaq7kSdJzO4U7nrJAjx6HU+KUyJzA3L++ti579Ln7odY/blXA
5nU/LL+8Tq4U4trl5tXE4n3xr0xwmYxSuvVgwnTNsbXMt+GrelfDnE6+hoJI4fr9mufigjChQnJa
LIbHRdtS1tJS5vJMzaZx0jP1FligCfTeS7T6zUPqvldbpBUoqRZC1ZpF17dpTewT/W6Wcqu1LPmS
U1rmwRtQ5OSg3BZg6Zf6+DpPVq7k9jvTZBiNWpnJFtPMtfHyVuStCdePTCMAWdrlwLfYAKA5MHaJ
8Poj8dbJscGf3P+tlNsmtGHA8IgaSEl5aKtGgUHnWnB5BBO13ROpuvkObjEc8dhS5p6jOR2avxME
He0pAktx8NvuWJE8h0t/U+5W1R+P9WthyiM86gqx14smcIC+liteffYQv2MWPSQyFmdXqd0V7Wdj
O/S4CPaTJU4NtBbyjmcRvKAxLFkZoH4rPv7TJDhhFuuZqILf9gT/noaBTaPAAcPmhN+FsxP52exX
8CcYpLsUpL7X0lKb0ahhvYLkypPDJ+VrV6XhX3usBvi2Jafuft/YU1jn8p7pGE3HcuciGCBkSrYc
pX0GtI96Pgj+LcknLVFkQtlhej+9sOYl52NihkMkW+o8NnK8HayA0VQ+sWt6gKPKqsZQiqCOlzsT
jftcnBc3BX8HtrPdKWv4+B000QmBCgORKR5BknJH6JxBe+/PeEbMY0t5IcKNAd0+dmpZ7uqPD88D
l8WWwmuqwuqJgkmRQdrzKWtD0/7PR1li01/A8P9ZBVsaviZOfA4RbzrxehMdLtV8OOHQGNBPKz1M
1ADoKgnk8fueGgFf2fxhnbgaBMK1PYqRJrmyIbK6AbzGHLWXWAKt5VC6rYTzkPGOf9HDJoAaKrlP
BAt+xnFziTI7yg5E9lXDS4RG+8AFbg2Iaj4Mx+W2KMntwRkqACq0rL2ib4g96zZD0F84NZqldV5F
xKBVRQ2US0eU20RgAG11Rn7RQM/a0Zah2RymIDF7/p0MOk0GfjN7o4cRbvs+qUeMQhGGYkfjzg3G
7OfHU+XXG+PxXL8uDL/ScpP+4wkmoh8dFIAHC/pkELgjdGr9zOhwEAY4nDxuCd7JhCRh8CBgAr6Z
Xowe2ylWaDCe73CK4d1GtPX4FbMndRxwLXMPMmVPPMvMBSZDF6uCaBfYk1R1M/Y2MqjDF5bfXjdK
OCf68P98r3aNC8JY/HfCz04EDNwxqAmUM6ushjVpetN+nJg5BQOaaxL5pq5tmu8x4F9P/zBMGLdH
bOHVnTTCeF2G7BNJeAX5fTBDFqNdBKcTsG4NJ2gSV9zPd++FnVVxlJNGZu0AysWhUjAO82HeDOZ/
pDIQjh9YohLiVou1HZ9YZDO5XFv/gGkg53WOM147RtXFeBp9inme3pFzBCfzf+HLqiWzsdbf5xkG
8NWSCeGB9T2iAJP46lNCq7E+2MrNegHz8KiMEMz/O4GgzysKfI5pAOZo9H1phnm41LN/NrENq4tM
+xLSS+mcom9IIGhzaSMT7QrEy6mUCnemrlekz3SEg8Uu2o9qmBlIkQYr84JIypgrRdO3vkUGgbq6
Tt1ouow+6GE8sbSbtnDRk8j1C/YA7i+skO4emrZOZntv9fC3sxVdxgR6Zj108RqGLnO+pptgjxkw
s/vdb0c8A/tjWCxeMXnUlwZHHPjvRuZHawOX1jjf1PdezA4MCbDZziX6VM3UypIQ+y7bp4wOIXCj
LNK50+df6uzHsjitBn16wpgvwLTeuKy1XeSC3/Hsy3Z4MK9ixV3ZF7GeJ+wuJQ6qAG/6SaY+8Q1N
SPzV8dDipexWI/cyidYaURAnt1Hc7Z3fLgr4wfPIcTjiGHkt2dITc9/NnJ/f5+7VkYO3Vj2Hov/a
UaOpqFnA81QCF394ng+5nlXJrEawsPojW35IKDLyfqzOBMHK00DehcDus5lQqcTphaaIeMYZ5cb/
Gt/xsS9f2iQlwrFk/w9MH/PBrkYHRP3VUswVeF82AvaChaBT1P9SqcHsasOpKBpVeVlg898FYbgW
NI0gXrT2jYBQC8IAEK80MNv4ecTOwocPoMRkVOIV+lCF+SHm7cIPisDAmPS8A4Qim2VOCWRvuhFp
mAFBYKbGiPixdGPdpjOoqA+x6qAp/VtBcGvm4k9w2qEvVolT2u3RwunRDvoYBGaR5L+Qc4f5z0Zs
8+3B7NugShI5Co9TGhKGw0J+bTklu71ketNQdhGmNgfA8JqoZsdjijmnp5nZjau9Z/WrsgzsQhoh
GoZdz3uuTy9MEaCODPCjR1eWeVbprm3WT0zJnoxc9d7k/jDYmvXiOjLriYgJj82Nbuhae/ywSSs5
7q3hfwH+M8iHgs4CE09PCU5gdhVBGbII4gQmfCAfsds1XYStD9IFv2KESYxsVv20FQmkr2oInYSI
E+CKN6dKZgCECA+/N2hsjTm2W5RjHnjpedGf1tp0MGUNIKYzVKcCohWrgLnYH7bvORMVcMvju2hr
YWb8ND2YQ+u93lrGUTfpPCasfH8ZpSV9ZaGXW0j2T7yRVSilbftBLTtz6aFKXr6VofVhNuyoMiBJ
Tji45E7ZuGoJwATLPmGOg1uYcN4R//cZjBGDFzkEVD3dRElaSqOYhcux6rmz5t+CN9Xen6/SHZfl
AMvelZ9qj8FqSP9JlDdah+hVHkfIxa0Kk9rq8x6gH5LIY+LEhncwQttzo3DB5/0h48t0o6AWtkZ2
E5dlL6y6+bNA2T8NRAhXOplVSXTMn6opJyNALBTXnl903tiFHkxFBTVSa+1DMm4kOCzdQZdZ5jcm
sikJ9koug6IcZLH0eD3e9VobSMLp7A56GSZ98ZtBJqFRdn/TRAQ97LdEgq9jbHKSEyU0Z4tSx7ex
uauW8Z7rIyvu0owZIArHTDvqFCwPG9hJxkCH9PAgLsG5CQPsPlcJp2RS9kbDkahyvnu4VL6rt+5O
UYn+n6sB1OPkiRcM63tybXWdXNUR5cy6jkX+z8zntzt6h5MMS3S1WZB/BSw4CUW9DK1KfpTUNio9
G6DUxnCNQFgxsagt48L188k+DvmfV7qHSq4iTX7IZG3tVC2uSEKcZrPoOqilMmcI7Y+eGcGEcFvp
Jzv8D0yygYXqWVssDEpEkaXE1NNHvY5+3F6dkXwjTOJOQfBMJBq/G5AUTmQ+nvzubFl2SxT5ju3b
SG1RT+L6saHP7OtVo1KSjQV2RaqWdTkBQI8pD52gR4QdZeT65DVMwDIrWN4utiC5R75yevwk+ixU
LGxfsyEkx+MGRvwKOfN+77dSDxvdG+JsgFL2q4RRWTAtrScZEzyoIzMuZal71sUxXWDS97eAnEuV
dkKXWVHLSbCoNlvl387SgheOHME0tq8uA3soBFCLLEeB6ahz2MEDVrRJk/dIVy7WU4l2wKJQVUwq
x3FWE3FeKSUt8+NQylCOguq5mKc5+xRnLH+padd/k7D4lyqSpo7+oK+KK1YAEwFqzNJ4CwHwjgA+
mL1Fr0TlrRU1jDPbeOqion6zt0WGFLRPmdEMi+7SyQ3WOUj6w1RGYzIrOn0wh89ZJnbYnE5gf0Po
WyJBOSOIKk4JB4dw/D2mmKlUilskaQ8Qc2zY5SZcMdDcfI9NQPLgsLI/AY3SzHBt8kS/wkHMFHDd
vbtWGMpT6ZBj9fman7BrmWZhgbiGEU2PGyCyb5Q7Nv5ejOUUFH3yTgdiYm4XIRwQjQVNMTodd9pw
bEGi3blCNnPr4MDkM7mhae6vWbLwUIb/9XMHtpMStmG2gq7UOXlF1Z4QbA07DodOiF1khiie3dSX
72QzYSUNwfdYS+Y9LDlW9cPzmK3i0EKbpPUIpuUzvbe6Zbai7sCn1eAhn232L688SWC3uTAmEstr
HAMYxbfdBCUwgKOyQY23KbsOm2pYBocH3hl9s/fMsFvCD5gLDJLwete1uVbT1CVWBbRXZpUhuTiv
Tmjp6gzQZZhAc5Lr0URkmTVKsoSRAKpkw3u33M3LKt5wZFoWVOaETiVN0tKSLKd9w80IrGDqBTL3
hJphrpr2Xz2VXr8MKsDsrmXXRUW2mpbb6F8eosuZsV3d+OZCVED04u2VxU8LeKO990M8SovNF+Bg
scRpyS5NNB+7GHOqE4s9szQ6YS81AeuQ3AR32olP9nXejuamTU5TVBwy8S76uX7q3kvICCSXHsY/
mOquw1HqIta3PxwFLYJQZKbO0u4gqtz/BfeAGdm19IjCH+5+XVbqayr/n5/U6TiikEZSmd8kLFZT
W8Y0ZpcwkGp9HAVSGDoby/dYyt09DKN6AoKFXhEiVQfyYJGtfFsZOumn03SD9IrJIV+YK4+mbljV
0f+GO+7gWtumr8687FxEQafBntExHm7XRKcAz7470foWZXRH7e7mDHJm06G+rS5yPH8EX6aYqZwB
iHSEu77eR1Lm5Yd37OH+gl8x8xjUjCs/5XWFGeUkRPBcBOzHryo6+ZOW08kgvjAsr0/HtTRhH2sH
+ciVMJY7re4Ow3z/aAYT+UWZDWMXrzXYC3MkqzvBk7In6rOxH7a6P5BQ3hfQ+OEIj3zaFw8160si
Vou+CZqWR+fVD1VdJ7mSrU7BjqIQx/KrRIfxkXqbJ1d/pyChZWR/nfUBuHV5fua7ZNyJneOL/YDp
xe/6VridVEsxIHOX7eh4/ypoaH2b70GzW2aIQ4lycCGWISwJVvTQGcq55afYlVafIi7J6gvclj4r
5wHotuyy+2AvIOj30srrr5C6AkFt2ycTe65xvnXPvJRKv1UtaHtHCiFmuQsSk5jeU+0YRNyOZ3do
huIFpbAW9G/LLZj2LwmbVr8LCIpw40/HenDw2PwqaPmJCudpg/s12+qsC8cLPi9v53AtdbmFtFCa
Nio9LbOQzkEsLkaRB7E6qY8qucSbE0avHUjB/XlivBeO5+DSnwDsI30mxxehPpFDu0JBnouPn2J5
J+Y+WB5QNpxzmamA27nRpp+jIFAwMZiA6jBmTXVeTK3MFugVznArCh5BCcs4s6afiRvL5QvU+myz
T5hACSMnsbUHAUH03TAyUugGUsZZ5oduFTuY+4eR2S44KjGRjqabPW77ZkZ4tZmGUBl+tBXdi5BU
xh5YVSYnvRnu2jf+0vh3QrxWGgKPmQuJ35FBxk2HkVNNAf+wLMStC96lemURXINYsqtB57O0sViL
1T/4FIxIGTuQ3vU7WT4iqMdz+MwlB6nnu/oD6+rrdEGFLuzabMAusSU3kA/18hKhTIZOmmqlpeaU
fxx4X6KxJDcG3Hkro4Fvup7ZKKrQB6MvRAeSBxmi5mS9MfENwU3NildKjsp6JRL+NG7msS+ixKv8
MFDJw65y5DNzE9oX4Sphl7PejfOKpTNRBfn8weQ5aX7uSpgaJTA5E91GCdZaWaq6uaXMxfujPw8S
BYY2+JyXZ2FCKSIS2DNWqB4D8zTuMv+Tesk3bf21tCCJEDcSSPV6iO8aJRlJYAa47UQJd6iU8zY0
DzkNKasvb5Yh6u3z0Fyqs0Qyfx9l50fIgyQzjOx0Ascpk1yPyHgh9a08bzckAhZI3yQDmCxRWHUN
2/orGDvlbBJA/DFV7JlAUAdV6RHsWLVaRratZznVwAU9KMUevmAUvLzZXj+4yRlpwvncWMyMOwk6
nMpj6Yfwu9Llx+BJi8JGlWamIbxdD3ZCy6FkuWSF+yBltrzUkJqdTBbbapzRQN6XKMTU7jiBH8Py
OxBqE04iTez7eEYC8iQ6E5YSCRGEJVPGgMKYAJN47WzWx1R5SISmL+moe1RdQejJRVuMUvloVZWs
UmMxq+DdQEu6DaPdPP2nEsQ6s9CZXVQL4frc2GawrZgP1Zoz52BDW+hdr4fl0YlMjlG1PDMLa5c4
y8tyttz1THTes8IU+Hx8T2XONrx2k506an8iNg+LCG5HXWDi46w81b6wMhA781pCq1yOW+6Tl3QI
0zTH9Lhhpzw1rpZZEWqG8QhxeKTRpw6K3v7Ztr4P4AIHxsgmbPbk6m2jtwCGjVfQWiXrjYdHMg0x
SFuDsGyIihSbhOjpxJKp6mbzZSNETYi6LCKkufkSq5IA43fwSbA+MIbzyE70sb5rJDrDIaS+rFZ0
hComcd4zinuWBz1+MuNV0RJaPfxIyhdHzI/d+UyrzM2SCxoz+mw2RpUUlnfDN/31cG9MDp1Uwqq+
jaqzFA/deDzYOTAE+99RQx5leBmGVbQBzQySVNhTUFkq2vZqNHXoFu7/6jiDo8uSNI1/aae4Jcye
gKLWgjei/KMLVb2GJHcq2n6yHIXAYm8VC8mr8xZOgKXZJvfjtDzt2wZ8yP9UUomlPwnbgDV/pCwW
TtdQgRjHZ7zKbgCmT5rwU4tiUCfN14GZNIm4GeufDK6W9IR17ASHQb7UW5s2WwukUXgX9YB314Ia
RxVg8sXURive/ZsU7sevZikg/kAnJhIJ6J1BF6bBXV3xrS7KWTcbZpGOYmP7oNUKB8lfcPdZiGzr
G9h2L7yzXRR05kykW9kYidoTKHC9r3OYYcH+lVypxOdDBOMYqJb5iS+ZDbrBEsUpjeTBy8oRjvxq
BwLlzd7xmHnlZmRYl5Er02ffDI0gb0WdLzaCoL5cp18ILa83FgmD1jvwc9YIfRTV21yPjtrkpqAo
L8lMOe0VnduSWO38nuD7U05pYwqiAUt0Nxyr3DimbXbLlSXojgte1runFxqPmE602cMd1uDZV2FN
MdxV7bUx6FYwlVl/5rnbpY0Zqdv6xGnR47n0miGnuSal2c0YYzV6v5FsaiHqATg+BXWuZxVCdUhK
jC2oFKCT3pVyH3v4lR6sVqaidiDVF7Vb+/K7CeNvAji7uZp+B4Ayf+cLp7DQM/1w8JmqMPTMdTAn
Da9rf2YPKw1BJFKWmTjCJ5oIE3YlnNwaK0ayW/eCf7fJcKuxO2Y//3zwUlxZQXGyE8X5dAOlgTS2
8rRI/rhJN9sgL80wWS6mgR8Fy3vO46gQIsF1OtQgQeI7pU7dK1tUvtOo2HljXzn+DF842r3Vvc6V
fF5pWzcEMrQUEdasHdNfg5w903gOMuJoaRBt55bt56G669tvsOvcgmyQA+Y0kflBmN0HB4a+Yqqz
JwYXn2DU6RpERNTlZjc7FOydJEdkvVH1Na+td1mE5baS0bcxWG2gv4051aaeJkGKpjUehQExFT2e
3xkomVFW0WSlzlRfFDp4N3uTWRXYtwLuD4HBLai/L6mQQ9Zhh7wEifu0sAwSik2NENse6Y7ERUYE
TMHK0k+MeArPvhWLtxPwY+E2cFziP9BB41sONbYosIFRcnswc9obdQMXKxvHCFERYTDLUVtOpxZn
HY9SvMqrP+mlaAVNuiywdYkh+cOEmboM3EVf+T5lAK5DM9nHGWntO5lGzwgGKtIXrlYYeiW5iUbh
Fe5IvsEXOrdtzmc3Xg+Y8l3HkcJPNmHFuVSDjuIUlasCFLRKqHH8aDd1xWdy5kGjTzZBcFtlGW7U
O2UZ3RkcXFPxX5zZQzgH0LtGyua4HnqHUrPHJ3N2ycOhbFnzJ+LZEY1NE2hH4naDxEW6di72qeCf
Dwl6be9ZKujcpt0HcevLIKw/N9b8qQysl/+Mp+U010W4JfIOtHTiI/R01xNSpNmnhFOEROjN0rUk
hFgqaaSS7kk+gygr/2S4Z2iBUQOF++tYma27IWpljUOK/uw59GhWQftuYJuv2xwU4OsotI/FA2UT
sKNw2rcIxLMvl6NeFUx2OPGZn5Z8ReNfBaOAeeF8cMjTBiBhR6fnXgIBZiQthSZ3X7PKgWr6fvlQ
7wG3dDWij5j40vZ2nHpL9ts+RJ8iL0BRyobTE/nLEzZvQ99plOzVcvC+Vs0DvCnIJahmeUruvdB3
bwUDOtQV4SAuFZSimaOva7pFPsLhSwSOjwHQn67nzYcp8eZKxxsenO7dJh83PxQ78Wa1YzLg8x+H
NZQ2uycSpWS+c/lGM5hgGluYl/pcgrING0p3qwgh8iSDlafLgVzAnQho+Hq0MdIljVenOTje/zbF
oalJnxDM2lA4UfKojdd0AAktBy+jNAMduFc80xDMJi85pRX7CpxSe85t2Ahjf78+H+z6RKME+15l
HpvXP76UgMxShRy+E80NC/FyXwZQNntibP9L4Ue8vm4lD5/pma3x/2AhaRbxT3FpJMbBZjVeoXpX
wmftg31rdZz9sdreCcUi4ecCS9NwstrwDLJ1Nh24ZzUz9D/dQ/7YQlS1kOO/GyY21QiF9esqh/en
ts3U+G8ARG6ZkpwwFmiKyz7dDbLmoKfl1G0aYYIPNH0Be0KHorwF5JXVnr3ruInNU7uYNDUDIGmp
3VE2OufywxzQp5MrXAEc6ryhyLt5Tq75MNbyiqKkDv/VXGfsR0nYp5Xjl/LwomypVoOw2evL6E8t
KY9EhRQKU3K0jQg7wdpyV4/PIisaE3yGxeVNyM8irn+fyulVRcNaKgD9n5BJ8ipJRficutHan/PG
RUfe/D6W5MGfBvZEtzDG/qAKuDR6ecqEW4ZMAypmQsx0zTNa9A3+mk5QlYJlNiThmTJRbsevZcz4
8iet1qgEFONyos43y+xDhy9rURooMoBA5Ukuv7KtXg8dMP+TVnGOvkF2+Acp1GH85cS2AmCvqlP+
A8ar7WCMg9sjC2zirMus8/+p7pfSxniDjOLCuGFWaeHLLgIrRfNAqmKykYnWoH1cOtNSOCEgCR0f
X2fSHeCNV3xaYheCvDyQyd2omo5IAOC8wxx/jZoHYhrtOZR7zf55EZgCnwtB189i7nJRFqOVcsEh
BB0RVIvi/pSWVj9/WJgwb4ixJPvP5FLwtZidzDo83kMLAhKV48SuvEY9cj8ngzkrIgkK4DUC+OGp
QL3aMGf3eUUJQRG4wrU0hnWKip7Woi8rt4hUuKBW2BH5iL2mAEbpnkj14ghC/wDys9Ls+Y3JCVVN
KkFfoJ73sIdHrcWmoP3QfwVxZJgh/vlhLJqL39wGF4cAQR9hw7MGRW/mjUe1vZurAhxO6Sz3CQo2
4gRTWp6DfekMjeu3dVPGlALyXVhTiqlramcfx5oui2p71j31a5OQJJ5NQGr0tcqov4iy7HZCKsRX
p03SwoWtSYxXlf8xH3zkfcT/qdCrTBPCHyhqJSdlzYefm+3z4nYFRRCffhLIHHJg+WFLtIZgdixa
xHNd9EnpCinpUpduBmxqdchcgO/KYx0ZksVKoYTUJsu/jtDd1tAr8hpUeZiHWQnPAdY/ZeIcY6G+
FPK7TQ9wI0WGGxVX7FreleTcTIVR7UXS5Vob1ISZm6gzmcfETGmHYaIDa4i4NPqAeLExDwyC1Ymd
qRG934xuyoRQC9Ibirkas/KQaas5x0gdlmsR4OG7OhvhA2iAlVSIk0Xb/S2QqzGGzQDipQnm2+sI
OZKgT15ihBG3qyGOXlMtR97eifR8pwEIsTGjKvPIP+OlRc9BrcvjPMT9JGOw+NsIZb5qs/E9EDVS
K/E9vCgeG+AfG9sYJTetsvbSTYidQvznff6JCu15F8EsN4d7fyaHcaWpxaWD1MZJFSdTJXB8P39i
gezD0n197CBcyDOamYSNWKARLLsVrytQ8Kw1FJzHTJhpqR6Hc7zi4skz5OahPWcWn9U8T6vJz2sq
Y8UFf4xnSJc2wpN5xtnfvfKpHxF40RcIoTSkesvtpJOOJsK81CvB4l4F5n8ZeK0bjtb9yfizVqrM
/vqhYuCh+5T/qz/wvvLG0lWfnmHY+y+ArwiCk5/86lfB4OD5yay28khDM+eh2qJ5Y/QXV+2JjkZ7
OO+4RQGYz4kq4yMIM17WMflmcicQQvrUsfNKS3KoRvGkJm52KlTBRVkebigbGuHMB5O8zW6xmy+t
Ty9Dof/SXPFwQPP/Xz1DPhsX7w2oKE/9i0Gr1wLuG45Yg7mQw69ek13w3CQGrKRtjVBMDriOpTdM
bgpbWhErRIKcrrZ1h9iff5HLayqdf9UFq0sCUji3+VCRtX8B8bDekGSqhNexejH0ztwIH+JGOQ0q
wStOXH3cPNdmFov0VWLolbienLaRezcFrw1FqRIwCr93ddO8PwutY0k6+FstKkGv49rgJcD1YLVG
d8S/b8a1MJx3fhTGVPocSbSONo7U1Q84fyKm9eYfebw7Oo7OMzCc690Fed46otoNrLzqh76OjZ3+
NqHrS9n4lA0PhE4eVO04yae0YrxMtvf7t0gXkhNOraLQQe4JoJ44LWfU5qwyzlunzjTojJbiHXL8
zZiWEN+4vGzzrgnlWqiq93Zy3lInG9esbbcE62jPEqrLnlzFbBrJcHf9+LU4cLYRWOF27nCvQNgi
ZFrfUgj6ABv5+B7pkp98ucqIq5ZcstTa98PwGM07C1xyvOYXRzVltsKiwxXG4BF+8Gt/abpWZwTS
QJtwuJDEP+3++8cOviuITfnzswR/SiDsRcdszSO0doVI68iVMhcsNyrk6+JxtOOS6cTAPYC6UTe6
bPblDtFpLAj1pFFsrE34nBZyNAAj1tBTm0M7ZibTeTWDp854umupq6ptIYjpRUTYbfPGK+bxGGL2
WTONeUdS1VeVjNj6BslKOY1MXe343AmFCVwU74/JsPQweQjeruIKC8TqbKnXSJgpqef9i7eGBsvI
Z7ujCbPoWcn4Kw77nn6l65y0zZ5VbkiUGCnv31UjUHp/OWCyr6Mj3iAIzrz6GybUTye25XvTXQx+
M8S9OkvhIS3APWBy+w7wYD0JNGJm+eZ3f9N6uY2ZJTJt0vwdKjcRG9OyIiejZEUKv6FyLPgXKfcq
+Y/VCG/CabYtHnS3zx88SfJETZh7nVJXcTcRF1n7QKOqbNJ80mQY3pa3NSuhhBAdQxTXlQgPhmhX
CA3wPmZKY7v+W8jQG6rw1JO+yTybybvZrJ1JSoTikwtHDHnNQLgaxBwTfE/bzDvp6JtXyNWAV6xC
PY5xYBao9KiDO4IXF3q9GOIAmHSihc0vGgoyL//d1awjqzWssaTg40sYbcqeMrjmUV7+pKW8QcCY
SV9hjP7VHZHUua3MlqSDTP9GgSKcN9XNDAnIQDPG1IaRW56a1h0L/z6jlyO3x4gqHJkJjjhKvJDd
Dn7mvTIdbkflLYR935NCezzXr1HK77GyI3FhsYRe57gVuC+0OBdsaU15k1e+ehAifpNZyh7y8AoM
c6nB8uh0bsEJSXdnFwPgyLIBiXUF44LZ3htSo8DipBXtv7+EDF52pRERgiwgihukPIzse8umyup/
PdfK2vspDrpeZj/fCkgDCkDgNR4wwYWpQbkVJctEnMYIEQr0Hbgi6w22kldh3VOjQlx3c0LXu2Ke
rfRrwPanmlKMf0z0KmMWL9qUVzAyhG5WSNzXis8eseovMzU2S2s8hYEJvq2IPYYqxsMl58ha/xKo
Urv5c/5kCBMjbNnnN/03tBgVdXTx46lh6k8VlASeZdRIrECVVRxpbnxO3Yyd9TFKlJ3MDfwClcar
RxX6CFTu1sQjw8ZsHpcfV8k2+3YAE3WkEguxIszDJcszDlxdarvCNmdDWBo7zPZ1/eRBV6L6Gavi
PurmAaxo5IJTNoStpZn8GJr842r3RcXvriRa99krX/3Nh5eZVCHcE2OJucVWng0zqoFzI9iN8QC3
6M2YMLFdS6srOcCCkxI3LOJ5KcNSJd8AYvTf+nvMmbdDu3AmYl3yaEVImdMDzEyJ9NKTdUi03zKf
0kIVa0ZQakGpf1VZZzvHYvzVhXuc2wwZbm1BbalUaRxz/eoCtZgx4+Ut6dMWbttH0F2QhXd6H0Fe
MXguYOdRaYrk0ugVQgnV0xp8kQdwJQmnTDwwbnj/tXhDBE+8n21kiyx3KgbPr8gBhaaWXqyjugtG
T6l/G8B1KUysaZBmpyKkOYa8C+KgkpOzl1IeA13R4g7QFnAn4wkxLpLGMt1UTOZRT+VL8o0hNwWW
rlKpktY712z4N9akL+3FJbqH46cmsTHbi1qrAYxdpb/DpHeVtQyv2xi0Mc0ZYIU2m+fiQ8JwAGIi
yyZPe3WFjxfbePL2B15fH+wuKLLt3jA+eBi5Z2peuWtA/uZls130vRTtmxz/wnSYyT/DT7Wtx0Y9
92j+u2X6psHpKMgo9ILFsXn9tRmEISMH1GBps40I1JEYRPhTHWjq/3wkI4LHytdx2aGb2/FuMbi3
qiZlTim47DKX+NxWWJmkf5ueu6LfcS2xUx+YE7W/YfQuU1UCFJmWBPk0yF0h/dpeN5j+8GxrmGGA
sC1KE4yqqLPmzFDcNJAh1ndJmGzs8lvliFYQBE2JgwhG4Qj6FkjPheh7BY2Mz7fYQ8FVVmjdUtQg
cI8s1RrIgK2FmKsok2UKUWZYZz+R3+Mbd36h1QzEtO9VvOoMjN2Os299gDbXwdm0UQELSdTDpZ1L
Up025RG1KKlmY9QBFsriPWFt/yXag6JK6HuO1s/FoxyUj/N0srJZc7AUL4P7SZ/cXLcowqN3at3D
sq7yWAGan/pzbkuFUwlFiTi+t4uvU1l31lBdaeBX/yAGdtmsf+lTYECbKqyRZge3sfovjHqI+dV4
5Wz844tiv08poDeG1hsEdYoYcgahLrdKYgES1Ib7nNnLpDqe+gFLyGjqFySH8HtsKuGWrWEFxtcs
g2gN8MMkP8tzMJ7cTspfo70Egtty8Yfrc6L+jTMHJssDc8kjufmIIfu9ooyWwNnQabQuy4xjv2nX
xoW+6FIFIr0VDcD5WMLmoqagD35gqea9DLw8Emqd3fNtbCWcZknRz5aWwNKoMrb+qi3gCYhbhPxV
XssWWQLhYAabSHrMeIicdZ3ISVXClZGA2KU2UwwVpH5FANICzb+RPEGkHtyz9NQqbobVpL4UOKh9
g/daZsk/Er83EHwzc/msYbIHX1G7O+dZqcx+5twk4bbUzb9YD+q58EH1dauLf02ABF/BHC+nbzap
RDQ+jjRO4pENDzjLGyxW3BhDz8ZaOT25efGgZrRtkTbto4BF/cpAlcMIpZwPHTM+GCkYUwSO+NxC
ynKsu3HE5WnOroiDSij+Gmb+h+oEbnV9fw5zyGlYKJOy1wNIy7pbm8EWxi41UvZY71gRb77CB+9e
WURHYHR6OhDiIO6KtQFDheRKYXwywElljM3eAJYCw65v63y2xP3W+JhqokdjgEa8ohtnL8Uhbqv/
FJ7Zl/4ZB8N4bFNMcNi3SLjLtSRPDRF4AJnOmc7fMkkYKUAQbkWM5Q5sTWDKWa05AogOuncbBCEf
rdtAM6aR2QxD2XvCjripokwx0R1AbLa34TJveGYC3bAMOy7we6y1RJOza4aX0oPxdbr7cLB3OB/r
A+uXYxpg92dyw1xWDXbEgbvLC+Oqv3IMxAgYuJdARiJhCE9Th9DDsjkmq/4ce/20N2C2U6RtKfsp
X9QdpqlmtbBO2BtxVGVJtJAjAOTh/BM5ARZ98yc3WMai0yR0eVvcjRLPKJZ8l/xwq4cUAgRHjjzC
CumShCpXdGh5O8mI2IO//7rfMq4HPyCvSjEhIMmbm6xueU5d3r62XVu/pDpNGizXhKXVrvZeK5D3
3gu7X8NOoaAeXkojTfaxzXQA9uVUdheWvdkRsF75KP8cuF+l09eQ0ruSAg3ULcolE5E/o9rx7MuR
iHFR1O0tYjKiqB73TQ+pKn0HGZTsSc37qjpFW7Q7TpU0xS27zgwtrH8LrYO03x1PhGAp7i4nz9hw
bBtn0326AGHkiWcrk9w9j/K+Gc6G2NMk+t1YR7XhGklk/vkySAgCKDkFUAcg6NOvFC5xaTCCH7LW
7obrsgjPRxyMafLt44SeGmTnz7U4Je1GN6U5wYRMBVemA8l7hB2XihbbqIPr+sjd8P/mNssCUOOw
IbjZP8wSsJ1mHz4eTFKUj/haVWtfENkI5u8znoqydNX+vvmlj3L9sQ2RIkD/nbFZgj0h+HMEC+Vv
xM6ZlsIPlLunC6jvNRmF77/BYDHmZIWb937+PcjjGtDoWqGw3mc5LSkbx/cYIvB18N5jjLBwdyES
UnqajzuREITKo3EtEpK+HTJa406GUJu2S48HRI/LPbhvIbVs/27HW214nhHAiAQLlMIPISz4EL4p
EoYC4xXBLbUG8+QHRddc3ZhC5pTgQwl8RqRtjVBINuzaCLbWKiix3IKKHFtiiHjOOwa7yW0XsVu2
PbolcvKSg/WOr18XS9vd58uKldMbUxAr9B8qgV1ZF5nbAjGjwtSbj5QFs1VcxhOtDH+CyA8bsfVu
Qgyno2tMDWAU6U16OWkWDwqPtpjjCSkhVx8pFYlhU5OevRaam/Xv1LDr+SlXu3rW3Q5aFwoS5mT7
fJF0Xnwj7vT2DZLtyfoXLZFoJNqfy8rJzbPIyCoj5aDtMd7ql/7Q5YC0R9u8YVnVnYdJK+IHeR5r
DPz1cd1v8EHZu5uNfqml0DxWlqXBAxHr2uyDrvvQQlbInce+bCrwVEeEr589f6o+YeeDyVS8Rfi1
AMHDioNnTqwYIV/oyfj9eG38NyTw63LmBf+/RQwBQkIwPPPCm/f+yTFGlaMxDSazuDI4xcLZU+yh
WX4B3RW7V44QiXW6/F9Ilx9ONpmNVNQvZGxeo1FtpQRwsgKSa7+1JedNoUYo/7PihbbTuHEAFrv9
r6yfpBiiGJuZixKyzGzJ7ygMDZCTKj6blOLpj/pwCBKeL5ocRQQlMZuJ7uofo73OgcL+ZIsGS6X6
PB6e+NGUwcvamrSQfUj5adiQvo3R41XpsNOXfo8JzO9jLZk7OwiVISv9VeQAdbPxyIBQ6hBfxPrc
yAjXCp7/uX6EZ7SPRcQBbl33x91F+7e5gAmmlpGAbEknryQeQkAwxruP5Fn69xGJO1sowtJTryrY
ddaJmkHc1sZXodVgIOlJcn8I2SOgL7ujmSIjEmMIo6fxVZp4uCmOZ5EU3yf98BVJSaSL9t73Xd8b
JDvHzUdo952Iirwo3nXZLwsVrfsHIZzHoZNlQgVGLMBXlrugdrvRbLbNrGzBgrazokpEtC4Yuhmb
zeov0rao6TKoPxFQaR2xcHpIDD4piCrJ8FgtjbeNH5lID3xgPfZgPb8zg1GEH8MesIQUnol+St8u
G8Cgvhx+ktwZe4ClxADtZZB9fxu3dfpvnNq4ZEXxltn9QT7/RZ1CTfii1QuYFrH4mL2QJ5u8TST0
TZNx41IoZ0cDqRRDhgq11Xct2R02TF5T0SAi2HaHCVG901JB+V+EBNJjpMSwE22ZCkAkRU4tzJ/i
sDBMPJXfaCAghPHJ9yswnaMmJoFaIQ3Ol45dKCBazkG6g6JnrAash8taQrWHmi9bjkwvQ5NkdgGb
O00EkDYI3Ww7qCdH4RN9lvlNRwuDJdjmM9YNUV4kYZZBiJuVN3GO5Bh3qZATum4QaVsOrJ8vifqA
B24i46Cr+KrCr3z+7YGSyMzna0zxhhARN21ZbEZkSQBSHOx1zzC5MTazQTY2N3wDS8q2/Uy0IZvw
8ZRJyFqz6IzLzYiX57Cic6TPBCuM6rf2msK1bZvYXH+rFqR9AGPCa4H/i0o/n/9spGDUnE6pRpC5
/qXOZgjKZriaeOPtAGWDMGbZ0A/HFl9xeKv6VlEXFZRE3DQA5S08TFO/01eCuNgBlgCPytyS12i1
gjfSfJ/SLHDL5wuFvEfLD0bKGBRD4Z/ZWiZtggUUAeIBsmNYj7Z7wdgUMFHBQuwYVSuPy6ehYp+C
6T4ZG3ZW2J7MQnX9gnChUP8L7DQmo/1Yn3hBXJKpAOYQ11l6aC6k0Bg3hmWAiH72S7l71TbKypth
jLKTRR2LcfYrmQDrM9jBB0s/h4kY2ToKrMIsdrwp7OMUtB2wqbRY94yDEHaoKIlqOV59gAx7w+BU
GcGHRSHI4WQhA6gZogfDJCGnAxyADN2xFJArfRH/tt4FqBINoMtNikjKFEJaggCe+OZaW8DaV4uA
gZ3n/6TklI8H4/oXZaVC2MZl/xak5HppZlqYkSkPCk7g6fhe3qSaVT7dnJSm+s39CqxvHzJ7Fei3
IgrYoWk74HRkI2bcJ+uuDt5HlOnKH/vXa+HruN1qBQYYMXb1zIAvbzFShgI9hOJSoPEw8nCWGyXG
3FWWn317MB5oSaqMXSpH+6r/dwlbvrBkYnyXC+6HrpZzIZRbCKbbuIu7TgO3z5Pb2uSXAGt4bNuT
qxTMDuaYUq/2QvSLnotwsO0xs8BlDoXYTXkc068+jjEhSPMHKPvd5N/odGeMEXKUkk8xnf1ToAgs
qsU/rsKPWrNT7yOTsFtNXcR7+BJyMSQR+bgurZjgQXCJxZUYt118ZVaMUQZfYA/8H/y/fjq1w4lS
rjijWx6g5IPgYdjEoKgvj0m0RbpCoqLRX9iZh1l1olKWkWYNZmn8vRs2AI1ESVtDK1mqYQE6WF3n
H7hDqSky1mg5Ab8jrHuDEKZBomeZyOXRUrTZV/hFgNk2FMOTBKfNiec+C/RMC6JNEXW0TbapC70k
wMw6ztC8psIYgimIle31f+RVxaBlXkJ6vsbv5ybhT1P5xzljy/NiWDDbOiNFu+HkCBC9/Y+/9kIH
l84LcTAmLzUHgEDoPe+TDAYPPYlDnm0hMYiVUyy2VEU78OOYzZ/GfnfV4iBfSV1KoUGpb+4TkXdH
eNkPuE+ehJTTetawzGgwakc9x39er6jJUQCV9SUo18nIeh5JGteZ+ZsE3W2EjmTe8vEAq0ScmeSX
pCKAzDVP+TZLbNLVMHzXCYpSgb1N2FRgEiNwLi8+YdtskMB1gRN4GCgesJAFCaf1RtPKId6AD7dY
9WbRx/T16r7Jcd+exJ6fGzda6kdK4qJWodWVsz10+mesCHcOg1RE0nOmLQD6POjrDUlsWzdCzDdy
fGAu+AfZHKDXksDZJOG+8SdW6udMOvTg7xr9P3t20QzYTta+5C/mClDfGmpIbWg9cxzRhq5gxDAz
DAeVgDsjv5wN19LxCQbziHyoU2X8PO6AnquFk4DihuNNQDgHO1LAdf5P7YJ1fiNKFk5lpYR8er9C
4vyhW0qH63gl4HAlju7Cias/l5aoNJOU/aajMlZRPtKQQsLlLWRZhDsO52HdhdD8bKJ5NdnDweNo
tNjIH5065eJiYOz6rH0VwlGNOknM9h/2/H/mQv8xhu8coL5lLq+G03gvQRKlaY1xpdJdsqQLfn1e
+qj4sOkjAtkKCrHd4/J3G03x1Zo2qB3L8gh/JkFCfE94fR8slEnAS2XQie+oghRaG1GJtUKngE/f
cMCIXWQ0Bu1RQrlawf74gpt13MfaMRwPzPgatBeQRAcw+Uc0t1Lgmr4cd8hZmnU+6oHB+ZYw87pw
ZXs77tIip346BhaFLP02NRWkD4pA/Z530g6CeAtCoyDXk/FtWmbHeaCoDUjcRzLTCieaSYvHjqCP
YCCSebj7gVHaxJI95TnhsvSFTF9QmcEdvgm+xCCqiPCaV7azayzj3fpCKM+GYZt0oIj7xxVz3ZoT
qNALGuEMPOgxdKY14JOrnBpgVowQuX/1DwW325tqLuwCD4YiVyxVlGFuX+P5CyRaE3fBvNQmByeQ
eytaKfkGbTKVHlijnjdCOg3TXSPT5WnwMQutEPzGxjwKxsKNGfc8Jbs1aG2fF7YjM7FgHORp0z1k
ccgXkjqU9FZvTkfbydJJAl9qyyU0TCWv4HmFcOefu6P4lSisgpKuxJMe7A3HU7DFfzNDf6m49MSC
Tgk9IGdxln5GOR5j8lN2Gfw1kpI11wrzuLuClkErkS3XAThhPSjuWLk9zGeHvLdduZlSHzDTc/BB
axcHzONVHkrKGPRwGURN7nzFI1Idt/lP2NNqkCtO9kngkl7HHDgmR9KrKm6PH+MGYUVU9Lt4kZ1d
bKF5P7Z97fU5jKufqhMBSz5GNTHx8pk77RbhOFPS7z2H8OW2IRwq+/kxGHQ6TpvuWuA0jIUUenx1
prikp+k8jVQpKqRcAs5AK8KRuxiEe8cTHKRe4IyCg0Fbm0/NSsPFwNhpZI3CJA77HzCciCYn7Oss
b/bQeti46KAip/Nt9rxXM68GqNH8ikafTrL6ZBvUextm2S1d24Pb0BHBIheeOCxJZ1GxQ5xx8T1v
EBZxVFyj7WsYycj/6o+JWNGr6NCpbKTxCvihNj0DKWokplAuC64ZPoBXBUBsQbAjwfpDiyWP56dY
6W0sM+EZoSTeaLbso9t6c3Vj4BZWv/Q+XYKQcKUeXBve0DQ6QqAs4sAfUVsZ956/EC1a7H9zuWaD
g6VToFCok2OnRZuV41fsBQZHbsOC0Ec8+kN9srG5K0jGeD8/tTKVZ1UOevftX+P2p2vqxfBLk6y3
k9jTilDdIpyUz2UORZAnokPpfTHKDVSRgn1T0qrGL1DExlAs8VSH8arSNDFtEoousZ/n+sxwWl4P
B4n1NmYSQXjQYb0upGfwYQBdmQHaVC+BbgqS86AYhBbFhWOnbMAkMl9IdSE2iAP6VZVNXX/hP8ad
+msDVwmO7XWjKxzOtxzSH4AkG038aTKIHclJfhSL9x+SjtPpcM890HMeaRkN7HyFMCnbP4pTn30q
fuhi025Pdmwqc1NLPu1yX9MSRHioojYfwDGBV2yorVK5faPkz5xtiWIMikIu/fbnBWyUqMedOtWi
re/xU1uaTVibvD8DCYir/6vqLMkhX1bmQkuAsyJx+aoWGqsBxcspxavDJnfth0uAbkiwOIOLaKxg
+PwpZmCMczyC3rLvTC4NTAqM/CKqOXtbc2aACuPc6lSzo6YcK/X//FyTADGnjEQ4wm68LPKZQAIf
k+rmbpKYBI6sUzdJmCmgzJDmzwJIXTEPOPCt4wQQKHmAgVpL20uPNa974MGh8RNhklgKcswnicp1
hpUdQXpufkGfqlOBDCR/EdSO0ORg8lC1YJRzCMjx1HuqlRy75TPDfJvTcBq9sBpnKMwkS1sFwL2n
xW9ZRyHX37c6oExelyIEGhsy4Fh+Vz1mcr5L2QDqlMO0QMepT4bYW9PAjMZhMFt3qUHmXq4QIzNo
5qCDlMvLbzFpu/MQUDWDa4sZ1WllsLjrt4zK9H1AJOYY2ic9GiP8l5aLDg+i0P4LdpUAkyOoNMqz
bWuT8OWZn1ZpCzVw1eV0H1LMKTxjVnzj3D2tkngTjm4d/0L1ZE/cJ5mnHkdS67R+DFw8AtbWUgxe
tD6Vs0Wn+C/p9h0QQht60NFZEu8kGDX300V6L8znmCEa3/qduRb5n3Gi6ajdURF2bbQo7KNmWEh/
GvdhR33qhIKBxknIdyiQex196wjOxc3cqLekXb/52/6rswHRU5sjdzFE8nG0r+ZMIjlKHrX/YzVo
B0hyZB+/bcmgO+hu8B6v+PUTZDJ88H5blEpPYC3bDEWP+AaLAeNkio29GOH7k3QNwF2lhS504WWj
bjlJ0Q8U08k0tohim8gOppjFBtxjyCkCpwYAZtaR1el/VyOjY4ADousuOmOGO9hmk1vU3/UR5eQo
lCB46HPhpDemjXo5IzfdDxx/kIPp7yv1N0J2eIxhQID7SKQLyOx5aJ7fKoBBD48HLQKM40e+ZlcQ
kCCMIs+qMubWfwnV+3SgiBDGGEA67VhPpOwgoRJ5Tst1maMw94JIlTCP+u9PuknRNumsVhrpmaE8
EI8DbTNlHr5gHq5cvtPjQQPOuv03cGfSBKrvXvyHJQvSRVz2MojENYfgzaKFFiqEZX+qW9YX/0Uu
MASecf/yXrqcLFQIOdcoFHRQES/9rYXOWzasL7+fhz+egJUIfCrreupbVrRTPU09P87szqTVSYpJ
MTqLb11wLKJ421wlUmo1M1UkzPWdCMBXYOdzmh9GLjv8mo8XKAUuVRtzyGdW0Z4EiQZRrAuq5PCb
HDHv15lZUvVw0qz87tPi7C8yxYgN3PHub3G0jSRL7Djxnbiu/c42PTuuyysFsvjNzcxP5o3ftVP7
Js9DOIvzp/MSMXNsqNOlra3SKXHPGWuG3C6GVV0PrPy3Pny6pBjkIIqlQn3PJg0fYEU9bobsxQhe
tZJFt+g8V6wV4ZbHFGfdTvWIrjB6uwEV/6vDujMH4FT5b2tIzExNaJYHClc2fACX76FCpxTT8o22
NHgotsJUmjgDeBQfIIOu6/mdsnMjBdDYb+IZWB0A/nwyBO04jQtq+1G56IW2OT/rbkLRisXXgB4y
ssasf1JO9qMJWKcMhsvWRz8aiH6//iccvJ3zjTwbUtQPDRQAFXMh+YEDYzXs23swcSOxy9/Qte7i
MaTWG9hutmagMlKYWHOGtklMvtyyioWAV2ZRYM2wH55arrYLL8HX2Gr70PcwZn+WSfYwhw97jLhI
RkIPh+uD48Ua7pq58ODO3orqQoJrKXjUM4Mnde1DWIIDNcGW5ZqiWgoVo9hvo7oRaxscx4LTDryz
KS2EHBtQKPbaUVOP2bWuGiFYzssPmRiL7Ebdb19i7NxCE50y6d+43wltSn6+h3dn16wS+k5BHBGS
+BQ7IHGRYxyEeWvzCVZDi79nWULf9jo4X008uGa0P/125WHeWnMMcx/kc3iH829cHqJSgLrjWin6
y1wlJPtzGsNB2RGakehGPQWHr9oqZKj/LAL0RkveeJLpHIlykLQkL82YNxK3wpePVO+1AVjC5afE
wvZvg3PZeWhG6Br1wbV/ox+Wnov9I/XU9gpnvd6NMa2dDnYzoFqsiIfImZ56BKjTiOp3IKKnBaT1
aIWAafc/L1LKJqZOOC8VywBoeBMY19WZkKAL2m7DSOY/K/tMWQ7lG9luGssBby7DwtO8cUdLT2IA
yZP0nQ/YXsBYNey1IXxJhCOP9iAY6nF0OinL154S30dUhMm72dIymzs1cTZTO8zGwoadsROVO1CQ
5fL5SPjFT6FEswBTSAOGWkAAIFAJblHX21/UDaatmfFvEUrAIgen/jcaDlpme99qeOf8gyGu8IN0
T+bIuUBp1r94eZ4LV2OHS+0nk44EUVStnPPW9H19vPYlZuhD+fD/5JFSC6VVlMN7K/VMlzzlxD34
Ul8MRb1BLYI+OmPIyfopcP0x3r3ud2+zYTFKXKVGR8vVKtpeu0J8oUNdixVCccs/c53agNGTLD1+
R6rBjf7UszVhYm/4i4A0IlQp26jvI2+l0Dlybfb+ZV08o1wBamM98Fg+ODLaWaQ0LzXCHd5KUWuh
s/WWLk7xHAfvxHYpTjwkCf/1i7RqWvzRZchKOusTMoxpqhkeiM5lZSvXsHsPvqTd1J1C9O6tDnYe
oPXys8uVZ4zNFf/4kZFRpdFc3lMNw1cFj21unMQhlq0ip4M95uwpUZZckl9/MSc1aUvTyZYB5wvV
akmZgjBxvTKHp5M4voUy0Pp0tZOzCddvSCHqzSQgsSd+o0tvN+W6b9ALyMMZZ4Wa57YJ4SAeBQj/
1ACpiD657j8ltexsgOhDz9eVqG1TsgNtejr/uPnUDg0a3B9fiZu6xIb0B3VdZG7B4R+UYgcKNCvI
pn/RlXRyjnTBMg4CfnCyXCsHdSa93lVrZFwT8jGGxJVYVPXMiI3WBJ5REsplrid8wEeaztG3/Kkm
ha82JsnLnjo1VLJWvNJVZirx7RomlMr9rKoZBqcLjDGZjpfyd391Z6nR8huyuOecauMgr1p0ZGni
7FAIBVndx9hwBIuc25JpY4jT4+8OF0onj9OpECnNo6t7flZ58gQ0dCMfmBRRObwKm8b2EjkjqTLn
+7GEXsqjJdSKiOt77Ps9+gzMd0ZLLcTJiTNvg15SuGFESjZRbUgcxyaWTyivW97Tp+kTh5wVhc1W
prrl1v8+fCvQSBbvVijPImaFrzCwdzRiHmxv31r20jfwCuiMzj6/RC2cRsU4zBm4gQd5/iA8TBAA
HIAFch870uojx6Cq0y3Jy7M/bJhD4WGXfN3xvpUZXfnxClxfZuoBi7YPewT3cMWeFQ7lR0dA7Ric
X8hveQ/sKmYYsh+kjeB4SLayoLfJgV5xPZqa85pp8OESI8J2rfMsByawbP6PYCvrw7gtIiB+t/yO
WgigME+6srKGkLQNBXROlY3cWtRNFktnB8ML/yFtgqPfoy2QBMeLNw7PyD1uJ8fFZx0zsHcESiI9
14CWazeVQH5r+18Ui+iRmi/8IYPnDySo5f5AmD+kPOOAnHwf5O/ORqvhWlIIDNBXIjjdZ6Hat/qh
jITBtvnUcJDLH/rtm+cP2nUvdE44OEYtza9isCwWLl+6yUli/JTHE9SGka8PYJx85jnBiNo/sT+v
v2SLaTi9YXvlsKKmZT0AwaTRgm4hqkNhrkxPnvMVTPakfCLHgcLZbDtFZLNoqf0dkjy973CTvvMT
vNFGsrX+lePeay1Lw7kheoKmuT005lbD4KXBypTMSDnCcHAPruXQaILbj6zbR9Hj5ESBoGkP/Ic/
kgV3AMoAT9YoFvMql9UhQ1swpu2tjf6uopoXiWimCiNhkROagx1kMOvOjF1+rc8p9dHqWv2RZGmU
E115G43Vj997SAYbNzSQ6ONi+TgeRKdm0C2aebxC+FH+q4YmGIruRX1bf7EGaGL1uu44rmrH34Z8
lhkcB+QQ54VRNx/xJM/tfNh1rhWlXqQupAA44aE+UbVh5cQE2bJNZxDrFFnNkt/PFAZrH4Jh9RTY
uIlN/4ZCOaIS+YioFaZ0VTeQbSuCcH93SHPIwpo1l1oQLwVCdua5O0P62cjokffbpWbAs/GYgjNf
BmG3+5uKKBqVq7SOciDsDuf63PeDDfNSAupegVHfnEqkTpWav6kTcjjhXiFDmZBOVFK7ChXbTdDa
Dc60qJwPVMuGOKtK/HC7vQoMA5co3jjCaVtKRlXbEcRNnqFk0y7mtqZQ1+fn+L8wUIa2hpXxyiQa
MBWrsUh/25iFr2Jf20CKEZxdQA9AVZag+3feN2sd4/LWZopjmL3IFFB5gLssTOCNozRri7TTJtbN
S3yoJjj5y7ufkw4RxEQBXXRItsWasaDTR69R40loW5OfvoFLc+a0T01o9hDONJS+2GZ7JgwAQ5Y4
P862iwaLykc5plDmROS5YZYi4/U4NBE82FCXIc7pSGnzV/DBfV3w85H3S7DtVOwIFlm96Z9Pxzq4
mxK9Fl+M11rvDrsUzvbMJzi1S2cZq/e9wbj4KKXbLI3eSlKlL0+9NrBz2L7fMDdmyrXKw0KL7Q9+
oU6al4rRkNuQnEIwClV3yR4mbNzc8hIXA9kWRmeWRPxUPWqXqnqVr3bIbS0ERJ/Fy7KC4fnRUm98
lOhVNeFPLeLiDkeT6XMA3MrzjOyBcdmYIBqrYuFcNGFOYKL/Si8UrZq15ZrZmwsna0fIAUAsDE9P
S7iqHhreaZa527R57eg3/KdVVkJCgq/hXGgIGbq6qViAMy5BpffEUN0SAXAIqO70bEDR7gCktx5p
1GuCZFSdDKpxpCRrlxu8y2aPNyEOk/iFxyy1nAQQg+gPVOFI1gv4pf3CdgOkDHQcfzmkalDtlzGC
aG4egvIXClW9qwJD3ARqFQx75PupPUzRzXThrKq3c3gbrA8yn+sKpwBAka2OwbI8bJnrIMcqGwsI
IihWjZMZVgk6/tdj8W0aYrxeJgdJ7lWmwp1OWeaGyT216Ssj03uiTPUdobdvCqH1zTtIwmz9hzGb
3Vcon95wBGjLPypzJ8HVNQ/3G0mJSLcUNYlbMADPIonYTNjGIx3qMQKsRn3cPgLMddccN6zKXTmV
0iAKH0bwhzRYLOiOc5dY+tkhqodnWvtX4l9TM5jtKUURWY/+Mo1kIO/OCNACApQi74X4JCrO5QGL
RfdT87BEATCprzA0D76/lF0Ifa4Kz+FJth235v1u587ZH0jY9BDTmUFRk2YJCDMfN8hH5pj7QOW8
dZhs6Wy9mg1ajcl2n+594wCRKSI0QqxgGjWWX+MvIdGrFHXMjuucVCqQpFJSVko6PI782WYBHMuF
crQF0dyjE+wl1Qqo7MSN6zi3WvzEHlDvoVf82nGfN6qclnvBxQMq+jgHi5X+vMgxkTG7W4/arQyH
IpF8PtTuOL3KjXiSFyai2RcMC01C5JuEZSnMZMIdzSlWdQWb2j6CyfiM1km4rDISSFHNLptcDHXH
dgwFXPbzKq8LbMpjQKqTQ1xrxGSm6LU/BsU2a2Scb2TrYxnN3zsARMPpOWIY0cjWQX2S3YBNrLxG
h8NfS6AMkJMirVbhmFXFSDB8f9hGvpW0sycOilRWTeF6/k9OCn3xJftHl32j82WQ+dsBWdQc6Zt4
oK3WDGbcyOVp2B5D77TZ09CGaoibpfPduXAAvJCmEzqZjv/qqPiG44HxivYriUCtpQeDDGRRJfQ9
6ime8igWQTQLgMG8ANkbC5acM4Pl69GnyZUeSEgW7dW/xExnHlD6WjvxzyC5bFHX5e6qO/Vbjww6
Z1hjV72D1ubqCbwnRKg1IL1xeWHev2GegM8l03ahmQbIoEWPQOLRhS+8R0xnHoUWpGGccCKhlYKS
wlN+MkCiqn33YtAZ/PNn66D66lWMqxoDM2tUffrN++IwMOMK1rKGZX+0QAZmOxyPPIo8/xH+SQm4
KuzYDB162PWdGkxADT/AqGCoxZ3wZCqTpPVaHj0HU+GNO4zgiLfS9iNreD2X+q1y68pv7NdHadPh
eNry1s6Kg5Obu629cRTC0EeG/XH7dnpECu3eHcDe14sKtgtMLZXOCJIOwNI4v9Me1dEEAJgxNdeB
L4o0AZgqP7EpzP1/gH9qYC/LLqkm4T7iOfE8rbv83QK8p4Psbe5RpsmKnTY/T4mfeAMjT/ZVh437
jCPOWgaKCjY7KIdApUlHWWf8q6DuJ2nQfMxFnHyHlSyeXKb3tDEfzD/S2LDvl8llGUXh7rqYewys
dis2aps2hR2UOsjMLVIkNLFdANrVtrGAiaKsNDtiu73lmN+YgVIvUkqiJMPzd6RZaLeBg4Tv92RF
cHTpmQyvcnr7aJ6CASPREXKi9ls4czRfKuivROEwJ5mEddVo0s+TJZRFich9bc5h5uijn6iw7HVB
dQ0oDCAcGA5fufIHXwz8dZ8cgcVxFKeR+V7o1wvD24m75YF0AhAJoCquVfz/sOUkqgXGUifD59gS
sNhkenHKju5kwyN3caO7YdjepKzfwUNxacuquI8tgMFvUUDrnUynyJAhYxOD3ABS74TGHQuLFqJA
DV6GooEAOJtuBqgl8ACboFaxUIrRpaSgBkjPAMHfvv9HBDs3Jbi5Ne9bUhEre6D85+QqUtuYXmPn
5C+lpbcsMcqONWaYVs2RwH/5aGpUnGURQx/uNaVJztlid/MsrCuEJDDiLfgaUPxx4ezVubiWXo3H
sUwg0yVog0HR5H5tpj8tVoZAzwj081QBaHYU8y/P3eSs3ZcILUAo3Ha9MKw6jmayu+t3adW2RcBq
/EFuPEAERdTnX296VWNPfKcP20rQGahOPijpjuAPXfcxnb6G0CgXgU9AWsDAXLS2TmERiHpzft0x
1QpfIRIFI3K225xoW1yV40Y/5Y5EmMYsOB72FLVl466wM7E6UBeKR4Go4VUGkSL0NSUE2A/huRro
4woexuPzNCqYYCnmr3Sv4p186EhCfkTT2RupfJfOprYVwTeUA/d8J0Hsuw2Da/BHTBMXcAZ3Ijq5
OT++92j8yUUpmdASTqOsdc0vv5GUtgUCUofHm+70asGvtSFj843a7Fu1cxH4eWFiGhOVyPx15ZeI
xgR/EDKXfLeU2P8gZm0SHbP4wLviKZADhu0otaSDPDyrufyRAjU/6XbEo4JhI98GL+6GZ2LrhsY6
LkRhudsUicGRVWocYP/sh9eO5PPxSnOBb/hVt8FXe0MSmnDAb0NoYkSj6zPGYRh1PKSEJGvOysFu
W31SxlwibrumqgJxd2Roe3Y5X8bXofIVc5Ehz0uWS1L75bC5/NB4OT/1viqiRMEjRGq6yMsoNzkL
5PTQRNbsVGWEG6oFnYZBnnMOITOrWPoYKOYCNR7TLUNXn6DWRkrz0SV0eZxFxEHwn+WqqJp31KsV
ilj0xzEl903aH7cHzWA3leBBh+cD7Gtv1M4aAKAMaXxRJb8JtRXXfDonYUPijMram37GfYWXgCFK
Zb74XKSL7YlJoFy00LhNValPFAY9fLQEZI2+MfMx2PPAdGbrZCCGvPgVYj1Gp9buPd4ro5wuAB+y
5GkvGiO3ugOnMaUh7XuY97IGpQ5Bb5zPCcdc3Gzwqa11GesRr4KN8TOVNEwnUiMQ62qiDySHUrkZ
qahJtT1Jv5zeOH6W7Lw2vmjwlRC3Uh7QfqpANdgw/P2Ou3nGkr1maUf+P5SP7QU8ysh3cZVbSOuO
8z9u6D2DoKGtDDnr7XdT2WbmPCw5WNUda4bsqYRERkGaFJT0a+VSV/VV/6ceQU9lfbyIGzJHB79f
GLw310Lo66WYd3uQeumgrcpBQOAd6UR/t1qVDJbr6TvNk6YPAjmhOK13O4n5YqYFk7eY3a9c14ix
WMk3+uNyP905/AEeLgAWWVACID+M/xf1lTfb/Yk9YWUznHNumkuNzherF33AZcVn4Y0sfPOhihQi
xWSshVQ4O+PPPgDm7EuGZBSBi2L+7+NrcX9lWEziinDPqG4gtL3ma6XKSAhXEyIjyDsSWcjKwymY
jyGQGclTlp1YinmMsI5zcOm1pfccs/eWf2hU8vLv8p5fvIpJBnda+2ESwn3fx5CLq9sKORp7IaU3
GCrZVb8JDJo16DUc54Vaxdr99+yG6FHWdMn1EELqr/0AjU3RdPdcjAhNhJFG2PJt/44wAxheveKq
j5HRkTa6PGSZfONiXeIIrY7Ae1Mj5axBMyZfm5qj0P+0KZHWmGIo6wGUxawlwXiSdxpOJcidiD68
DImr2vMMXxoPu52qJFjq12D7hFd7hbw+b2DPLy2Y0lak+G0qim+ORPN60YAWWTSOHY5klK+PJCyj
Vz8ueV1g2jDhzCeBP+EUbp1YNaGTeGjzCmL12G6jXB8IRQCoXcUdhvxXurRq34YGkKSEEEDGeoIE
j5TXSV1tXXZnaHE9rXBT4yn6MxU1woQ3YfgB9sGpChOTxZjZ4rAT+elOl9IcE96afhyUcSjxtu4C
EC8FiOxL7vjjlR28jCv8hnavIZzgqZD14oAhu+/vnoTh+cYBrsnZyFNbnneLmaayozyaIR2X+0Xs
3w0yXAYofXGT5l9Z8e/I5hDltvN5M1QuXhoW/Y2hI2uOuyte6iPIgDzrG0zWn6eAqIJ0JyhZR+Yj
X1LsGU87L6fKL//gaRN65F+ONfGtjFS+hbz8wY1P3x8VKXIIq4Qrhw55NYu3yxbneSLtr7ygMwpr
Oe3NIrNdW0zHzIYCxCA5FMxjw10rsTPMe1hzDn0ITmOoy4YfePmzZo7Kj84pnVkywcKDmTcrZMDI
4EcfpzSuWElQGCC7rgMj0si6/o7RnnagRXKDok3kps0TfTEDj0IsIxqaqjlqgnSOb3SXMOtPAPvd
g4RBSZ2fROGthI0pCz9gXgtMZRN3VP3UtlXm/mE7364EVYYNyv1FEd75rQKKFgWQBjh8Qdpd6WWR
hRrB1E4bVXrz9ZYlvsSTt0ZSkZWaBKsFdMhhUyQmdxALOp+MtFHgjpou6EIQmJ4wlXFzTnhRct/C
B7BykoHs2Wb+uX1YYVo4cJoBWSlw3eMNM2toFxIFVrZKOOprMxx2Yh9osN2nqQ6+UrqEHOwbNlAy
Hi7botUlUujXadvnD7wC5T40J8UQTsAlz0VRWUTV/3YledK8FGErFlE5S8EP0krdRxU/WJoNrjiy
mlBfWn5VcD60cK5HBebQVv6jAPQfTfzZZ8/CBgK0zlJM+Vbq/m+k8SXRxOw6ucggq2FctUT44oPK
yfjqULTJb5NsHX6SPn2c2yq5o8rUfuLW8XIJrGae65pGllZlpGXIPb1qdNnTw7z7mxkt8XHk+LI8
1DSsRr9pUz1MTfh/RBCtN3psOp261qC1OeZAYnf91bb/nMZFb+F0/iaNP6StXJWZ3S4s/IUgKx3d
6hnRBuuzv5XaYgPq8Dfh3Aq+jNIxmuxZY9NAeW3hSLhTnuFcK3ncPybBtaf191FpNHkEYhupT+JH
Py7IznmcwleV3sx9UKnQtB6ayF6xXPxs6Yta3JslIj1o5Xyazy3DnIQzvGwMOPbOJV0lIIRRvUZn
1LjJtpvKqylwB1T81HNN4UeGWPxaacS2tffFg69r2fADqiBgZdeiZPVt4y6kva72hkvDKjItX05H
ih8fJpZEijq3FFdLtsasFoG1idz2phiLBZXpPa6BP74urlXbuU3SwCgRB5dV0AaIfzOaSsk+ytmN
LgjKvHhV28x9gIIwqT/Fw5pysSxO7hFja8wmxWYSWzhUiVrEEn3kcaS46l5bXo3Ep/GDiMYtxRzl
W9+upXs+J5UnwRsq/uMR1IfbEYKs9fk4NOWkVqrtXngE6oDLmN4uripisMzH8kMbLQSPJS9a7pYa
PkyCFCZyyMiuW3YrxUDmXYb55tqIQqpcQ2sy6RGgInrynNQXUdUmWjW9MX6Q1YcHgPndtrOws58+
ylpxfm+VKK/B6MWTBZ4p568XBIqLvGjPwFEgmIy9cNiuUMWdy7XhtfxVPCtCKfXbxrVqXVURoMeG
ldEcddmx5USRZzZSPBKsuw+FXWYEIw4E9CD+SMU9BVk2tD1kWvtYJaGO2ip0vkeynigcI8+PXaz+
OvCCNZZEVtUdMk3AvIhPpe9enVVaNoquuf6RQeuIRXXkkHNrcilDB3MydaozoFo7fn5DvQw/0gvt
9723MrHBt/aju611j7R4J8dsmnSbj1SsverF4zkIeSxhpmwkurjPb6axuPQYEuLkXBCjQ6xngnvW
egF4iUD1M1742vtt662u4yIoCji301PXVzKH9Ivg/lUcPerMSwx65NR2wqEwXJs/a7wwC9XngXCU
RgaGxxdj5OlK7f+RlVd5LDEB2kXRRRQ0PJJmIz3jymTSI65/vwPcETaYHtEilo8MXKV5/h6eCksJ
+nfdriIEM04ZGDU6t+p89mPWqazAhBxW+rZ3asBPxLJKd/omXbfMJtITS8m/10xfIGTbC9X/U9iE
aRnZSNzvK3kw258YbcliDielU12ozfjfhGnthWNcHKCQ9uQgOeMzeeFcYjZldRw2wrQsZAgcOUfF
JlYzxw5vPM9AnJnYcDYBtyHjMs0JYJ4bORzBGuYq126lZjTCb5ckaKC1H4/X0O25SY7+cIxkGczQ
NHRlYIQCU8eyihvtWeV0WLEVx9MO1bYMQ4VlEXqpY3z7FV2YptCsa4EA7FAUQ/Qf0EnS2mmN4WnG
U1v5X9H/ZXhpkN+pzfLGSg9jkzNoh18ixcO8bXU9vGJOCi2dPQWD5R8u44/PtK7dGsjfnAFWTQoD
8Pvb65ociYmWmLohXCBJJcoTCogmNJvJuJxczMnfsPCAayiNhZ4xTdt0OUvk2sWCjWSDdqfdNbDT
2e48h0xkotgG8tBAtXuWeDAQyVljlT9yBzROPEhczCoZ8+zaU+Omv9MEDwz39KNB49Qda4hqpEQN
B+NLSGKhvuIs/ANLC4CjhIFtd3xKAq4wJ1NAtrsgJMPPwxkpH0u55st3GvVdmTL4AwhWbUsC9JDO
CDVxdssakatFN8vSWQreoX8dqHv6RUure3WvATj4/D8gasj+wO/wQsnTce+MCQhvSFFYjRx6W0a8
nSF+mXGUdNfVda7MTPmefz6fuS1LS2pv2wvqBrwb9NcCAxFcNqB4NLsZYteP1zajpkjH4JmlM1QC
1f3Zs1ZGHe7EGxHGoIfp1B78L1O193oO45yk1mclOea6GXPQbtRGBqx4Z5xK1dhgbuaW0ziqOduK
Ac3KCS1hFKOw3af+D/xL/8qCGPiR4lL0EUvTw2C9Zf7zXTEPmabUZ+aWPLRJph0QvmXe1lM5Uo9Y
iaOwPhSxNeTwYvTFT/hrkYWrgXxj6TZA2L7wSDs84RPO9cjyG3t5p+oLu8Od0A59e+RshBu2Dt++
nbHR7EbRPdDuNWde+8DqAHOIX+fn9Qd5r5Tem8QLen4bYGdIUgdcBF2sF+dEAjjXds6fXU2FvDhz
CMchr+jDvvqhS/hWwqa/bW4rSUjUcGXytnimOzX7TGae0S5t6xFi/2gCmE8YXM0ulJd3Sz1u2ehR
5lvowqmIY1hD28wo4z7wg9cibsJ3M/WVVJfm64f5ZR8Za6VD8xkaLADfJISAgfFkiDZsVmj8V3kZ
boOpsYqjkXtMkNeJZdmsGsBYNUDJP6qR8cguEujpbw69Swbs9877m+gpsPjFzDYyPR0lPCo2wq3Z
UFRgGxmIDAMOK/92TRBcqln6cQoqav+7rL0iAyuj5f2yO9MXnaW3NKsiG/W1pZxWjgyPmEhVwefN
MmX64kBAqF8LxHk3dTAJ1/P0PBCO3tAmeogMXeM+u8iYJNI6uSn4Gkmp+n0iG9x6dU8sA/dizMaA
Xj9gWH+8kwn0j78VH4Po7RayYeHai68rQc47KMwr9f7YtqY1CSZg2s70JKjfx6e7g44y7uqM9BOM
AmnPR0ovAcLL3rgJPHY3ybI/7TvU4H3YYaNooDeCLYrX5PJu9gLFSpXudwfGvlvy+2RM0Rcsu1H+
fc4zJCYrG4WjWo1t8IF88UUOrXj49M9WeAvj/tGXpkyQMR5aoJOfEK7N58RTi2ZWsoms5Y7LBCHs
yE4ksx05F8dxTYS9Sh9qJTfT4+YtvcQJn0VRUNn8W8/cWGM4O6ZOs8/P9yM+y9J0JgRffqaSKvbh
d3x4+y9WCiR2XJaKyDWaq+QY1iM3zfjh6UJW5KEYL7zelsVXK7FIlsPf5bsUbmjmYuG0787Ztz+M
JKmh8UihZJgFs1NCe+nyNgrRtqGJ/MqrjaGboXVw3aS6Yjuj8xOQ81jo8/0lVoi+lMisSS/WTJa5
h7bCTA7+imf7h85xifD+0te8iCyRLetH3hGgv/1aGYU1EPc6Lc81Il1PeH+E39gwAmHE3gsGu5XZ
2Hi/Sae3vLj66taNSeHsPNfQC8taqWIB1bbqGqk9giwtRUGhdMAMRSFeS4MceXxCDi5G5DJA12gp
3kHeEiZzPz+iUi4gsJyd6ziuq27JLvj6PgYjnY3pFoMOopEcHn1oTfRF4F0QyQe3WkGK4oSClJnm
bJ7sFnv9uP3G6QVdBMOsvqZ0PdlnIKd0PDq/ahHFFBsnmUT+45lp+OONavpM157S7Jm8gxbYmlAR
PTQALsIh9nXBHH5Q1I6Yep/klMtQJokcPnNPsZ5FaLAAAq2DoX+7H+BKePzLhuQ/IkQhlfcLYF+W
vJqK1Bsok4Rdeu11+nDM7VJ9xuyuEt+eZ6jQfGHn/S7AsZQws98CWe5libz6iM0YylywmbTy0STv
fbHtBm8enw9h3SuDIdPTqmYuJlrSPJsScLscPVdTG0txDw60tLTAqFdCK4L+faIXZ5+3UE38l6G+
RAd+erY5SD/ofR5CPg1d+wDwvg7xtBAfwe+1j6DH8QxEzSmLmvePbx6hn80Im/EZf+807j/dYhe5
7pTdO2Ns9Bkgjwtn/bcnAPG2LUByIt1SQLeDErBoCd3nK481pzPjcPu/SUTSF2OncYNCOtFeraVb
4YheRc5VJB8yeAzHCFdnJd/rrhvOSX3n8fw+cpRQJpBR5VCHfL8XbAtCSh2M7Lr1yixNQVjrkMvH
IBihM5HUGHOlng8zhVcC8XERTNXWd1bZlf9KVt2IdunjRYlo3TUvyrzWN3oXRK0Nni7G+ptdSpQR
A9voqCijz6cLhOqDozodNOkkrnFaCo2y4nXK2s5fQaNvy7O0BrNvvwx6O+35FaqB0UFqX6EsBezU
vVYhx+u7wFBZqatmJxWmvFOOsIodtKAkinQyjXGOwZx5vm9YNfsAusaKep/0/leXVXo+Y12Ix0G4
XG0w/r7liVpBLoZd3iNsUtOXJAu6lr8/4DPdSoNwEx1boODt9vURMWirsSIrn9a4rqWAAiGaIxT6
W4WF7CaZermvsKclxhdZ8uh4RwSBbWy4EbE+bizjruMIrd+1PUz+e1o6KYll0ZfmuMqc3xAfCTwU
ia83MmhO/c86cKakmsYZoPSsWAMIdAhGMjDK3wHOBKlPLiAlCGRrWmynPiQW2hsRWnNuaQz2RYbk
ofhusQNAJjaKCT/Dg+zJvnneDEiLvjZ8tQuDbo4jjxLBq/cl3IipM7VBN6INaPU3+JEN4OC2jZAq
2Q7wS0hGUkW2KuWKb/l9TnHSHv0Prdpt6fx3q8gOqOgAlda50wbmT0VGpuDrvYek0KoOe8OBX4Zz
G5nAKraidj+92uA/hAl4E7D4TAfzflbcPaGO1xy/HYQbQ/GduERbxSM70mu1Ay17uP+jZ/1N7Ymn
KJvwG1z4AA3pdLPoBYDIqn5aaT500fKpftx15bcxlbG08y40y3SS6Hg9xN/gmtTYjYhS2UcSgkgE
31zGhpUXyauqH9Rg2WYzSJqV8tq3dHXET3Anudh0l7mpi9x1VMMxN1hlLhHg5hskrnKBBGvRt4VO
gzBhaY1o8RZ4rbrvv/F2IbnpFDYLneIJu6AAeUguxZxIZ2t5SQEywFE2ipe9ptOjgEoavgj6qWYX
NKJM6Ppf8NcMa0a+3uBhXccfFXjHRbwzCYRJ7LXxbP8WWgMxzN2rNyjdFRooLL3L3aoBxsMHXT/8
6/0GYHvuNojg6n/lyDDkfGxcW0HFYe1/fhJNi+gwbdKtoGWdUk6JOf77LKuujM2yQy+egrxSdgGt
yImPmP9pGSCx0+chVOt5W28qo6x/tFqCSVY5F2L/STQsV1dB6txQwAPvYyASmK019Mmv0DLwDObT
B+ltQLXD6gYCfKLWkgbfeZuFg6WLndPhdIQnLx3dHG6vWFIzp6u36H2Q0huMvwBiAIzya8YvSDE9
YZCe0XJHaSnr0xMgtFDL3cmWQYg3w25s9+Tt7VDSQO61DdqIs/FvA7YNS79XSzlDv9T6SisQTTg9
jE6ixCBKUTF1Lf8sFak2/uw/94TM96lRQJNJ49OfIi49OtsgQauQX7BmqweMSX588j170T/kZYMJ
iqsJTeYLW7iuuoJaiHzBdrLrfEe9H4+646TS/sXk3Ol9sdzAV6vTy/h+JsFNFsS0ETDRvpHXzHZd
s7vUQoIwZpwDIXjuWTpPV+97OuAMGAX5vVQCeghDZuE6I/ukzqvSBVbFFBKdjFY6qyEZ6NDLhUaL
qGneDCYoT6O495m3GqefO2jNlhSy4oLESGq1LQvP7iQPkh5cX2DNgvMxtC3DKJVSUkeeOFJXEo0R
szSfixaZ/gE5hTbTdpWKgQKPAr1bI8Z2GWfXmr/MFOwNfoGCFOHv0zReVUN/fHZCsQIo0ux+uzrz
IfEMk30hFT2K3CSGBxptWjF7171PDt6Rh3Fk2DMi/sE49oDkys7KKEfnM7FgjclcOBhgMvtF9mfa
vNVUq5lY75IksfCRoQC8+MYSe8laJwc89/usQadrom+IrMsfpV4mInus+6kImeMSgixvV48SwJWZ
3LWV/q3RGPKQ9CH8JrPk0ERR/fMJRBM37uAHQXgKRpUKJ867AHYgdMLcKQSbXTRZMq0xVNtN45sW
Dvi//eVlLdOue7u6G0YorruFmfSVZpuEd0VGAu6yhFjUNJEwd4G6K2APzvCvZcVxe4acu4L0fv4/
XBpxne3sU2Mg3ZnaNJX84GnyjMqM1t+AvH7tR0WDclkpaL1vqmZKFGM7lGUZhwSlMFg+0uqIT1DT
p00nMsmUXY7kQOuKwutUxGoiN2+e/cW1s+xNDv49eEKlNR7zlqM1ItFT5lCB7yibVHngGFWh5k9j
eoVrsJbsC97+ap1Fg6pBbL+vNWj+tU8hA6hmzL56jqaHaAEfokJcB2wTly3gUoCIH4h+EfJrf2sL
lijrt74X8AWq1iv84YH7P3IeU0KgruZtkNaBRxcxDyuPmIKeVWfSpWe1syvfvIeBAPmo5/TjFyJj
zsgwhkVCgf/iyByI9ESNrkD/mb4WO6ls7SBlbVdSplEBvS53xgQ6NlT3Y76vvKoHu23j+m5GMRuS
honqueYfAiSk0oTEuas4N9hP4A7yIAQQJTfN3/E0FHJXlh1EGKSCnFPITenC8xrint0DJEu1EHg9
JG+eDd+MseKrY/w00nnYPAv0OUAIc4jLLYw9q8f5M07fGoku0AU8FIY7zXPNbB3CKjGsJgosGIQA
jj2ybl6v3wJ8Ma9L5p5JfSFHL6sm+ssYY/IacwCRP/Jur9aKWY3FaUr2ezFh368a7iEzrPgaqeJ2
pt3fL/I3nekCrcwgA7b9ZU4Bd54tNRzlNduEc6BaYlynnDwq+2EUSrEQWvooKe/5/PbkboNZGEtN
YtOsXJxkaBUN+adKWOfm+7QkKAYkhfO6jxUiJhu3pfqCLY6g0z2Gxdr7HNvHFtz8UZgKPNX4kinC
dFeLWGP3KGYAAfdVmCxXbBccaYVSGKkfLFc0yTVEN+jsiytA/P4kRD0KH9oRrw599jS7kBwOdvKK
c4uYCJH7vygK+9ZH5eBZd+66qudiSwm64xDSbGR/xl/Gt8pSABM/VA/uxKBA9ShMuPIE265JcJdS
w6cFOGPIIRQgH2iFB2jJ55bHNzCig1uP3NYokVBtJxuvBWXJW3ceYPi6RNLw/l0Xi0PgekVT5rpZ
iYSxMEZ2ZcSQuSvD0lTaeU0kL48LoTsoeuxZzm5ruiPBWB2+sfrT4SVpqm6jOM1hZF5c3D9XY5/R
tI0lQEl/Ho039wlTYheMYxC5NuWaJxmRhoYE50/LXRDhPnctroIzVMz57mx/YZ593CZd1uH+1+CJ
CO2QcTZG9UqQycuI8pUZ4v1fFkl37w2wR51CdYtCy6ymjvBbwdI1C12nyEp4DeS7S/74SE7HDUVq
tkTHXmOnVbaitoK9MEwYHzydruf8QnPYiJVDMn8pC0rW4+KxXtcxaAVTGAN3H/1D8uNf1w2e1hDB
9vlxOkFe1Bgb2wkAL6b0IGcmPWCZ3/kz7gz8ZkvJV4lDpwzN+8OEoVA/bHvrBc4zWlAohQTOuWO5
ihCZ1EGlVklLBK3+6q/VtIP6oI8MlFcFXrx57+F9WM4+Rr1XSRigodTvtOVEejNgqkGaiJ4uNgW1
THq3sibayFrErY8RJiVQmdSxa8sOYx1uRDmerAgpiNPPZZHfJoew9Tc8DRayzhL2WpE8q3Fqg5bT
mTKRmQ4oRaoThegOOT4US+1q6IsvwAzMVX1CsQe0BzC4T4ku8Bj0FKrdhk3AoWiAm1ksb4oFKLiK
FNcz3FdemOpDisOhnRR+CAb0FhOZ0AGYTZkSazOZlUlDZbJMvExzlXbjVql8+dM9Ag7S26mwOZcA
lbbM/DXQFKOm53ZxrFSWfTokky4A4cZAE15LP4UGSheVyFQX1oYABXrfJ2goFyQTj5ooBnpXtKrh
FfKa5eTwZtxG/jXVdoxq3kE1r+dqzTx3of4X5Uv0weV+UtP8DxSU1XZNfAk+qg5VCJPIrjlwEV1X
6hMvzfL+CV9uMVQ/liD5vqSzahb8ax3Ozfb8JO/OJLvzZ6xteDCLy7d1rqFpp7ORM1kgaLC5UPSF
23z1Ew/nTysu8iA8oAh20bPT5GD/yfi1fYKb40CgwUSYLYUMCpWno/HKwpB+LULAs0nujTsa0LdG
2eAFdkvLXV6jdO3ciqK5hM+lLAmBx3WjiBM2LEIN5Kc8R+UAEJ9NmrhRHMP52C0EDmDaH+iUkukm
liH1Qw2eBAJ8XNzQAQFV0iuLjHYgnTmQNC9mImhBFgbgzC1B9ixIH5o79G0TSTRZw67sa+c6ED4l
ohgRvf3jZz3K7xPPfBkVnj2nvChOaZAnzNj5LzOlzlYtiYkRB1oZo9sdbTCnnxiDc9Lc0zfdkIGs
JZRiIPaFdJJrSa1TkX3KyloFXZY3SwFpa+LXIAiZsRK49/7qBcnvcgmSniuUGvunXZ7VZdBvXruF
cMEKpMr0jjn3a/LtJmrXyy+tr8IrWIergkb+gXX9e8EO5zotht4IE6mbJc8wUOvz1/9HWYbNhRZm
LS+LFQ/L/I2oLemyHfRl1HOq/gDgcsWNE0ia6DGv5RlsLmkwKBxjTMVe/SaSaLWHxRJ97s5UncGj
yZAlqvnPLnjTKErRe+HLN4FvpsWKIJO/XJv0cHxQXjsutPCoIlHIVp7G4TMnduiyYP/EzB2/S6dk
ksElFgFcfiIiBUcfS/pNzZzOuNWFtivZz2rFW4abo4aqhHFXrvz6tY6zTO4pyv+F3BVSIqEgupTz
OLEQNSfiMejZdAjCkmQpD6SWieb8DVdSakIW2/g9xNCqCBkYo/+T9AkEQVvoAvxB7DaEObba4M87
Fod1f33EDWG2bRrksUUVm4qTaKsT8ZleGgig0j6uES/Vpb2L6W360l41cowytu/G7Bdw5RBisYp1
hEhsaNqY9RS05lpbYxRiWaO5aEHqbhJ6ecwHq9eR4R2TD3f0TyuMSP5yYv8mVnFr4JuIhMRspz7P
q8qLo7RuPII8WASHuOEsddLYchmFAc8wCMYhHXujH1O47EN4ZVUD9mXTpvDsjglpeo9R4j/zWNcL
PA0VzSLlZu/33mCmBThK8jXgqYW2DmtL+JHfBCEWLlzHUU/f3aheOdPmCB+Bxs+DTLlDT8fMCJEv
t5yy/ECNTnKcBA8zv6xleHNXr3ALLB8I+AWTXokFBJ7S1xzufUEwK7na+VBuwwP/pspzJcJN22eW
JLyJKlGeVOtzEL5vbdgRtwGGu7dnwJ4wMRjftC401yf7obXuC2VJu3hkcJQVNRNUjphCPly5n59C
yGc0jjoBZCF6o3/2phGaP0YDxu9W24bBLVaViCGtOhb72puqRbUBsYjCnvEJci44lVNEw6wKG5HX
ji36rR/ekmpDU7TjyapHwX2y8CUcY357Lk7smryggX4CrWORtOEbc9/M3KThDBQdozlooY0rAhWZ
DKlsK/wWV4czNNYZTKyaPCS7QPA4xA4joeVkTrFxwmbG5dy6HaZBZWaTRSAlmN1/QZcHH4Jr89IC
s49jkTGIDLVkcicOW3QFtnATBB8crwMjRRAHzs5fTBx6zER8t+Zqaaq1GlAq/djvvagEj7APdbg+
uM1ReP0Llkz1F/ZBm07ud6+KDbzoBqgum+yFIIztvR+ocjRiL/mTUgJEJcu+NylooEqEwj9pdTGY
6FcvUOLc5kOCO270Tuxs07EVnJU335+Ueou4QvZeGxN+PoRAg5/JBnX9mb6ds+EM+1ERsL1w2AyN
04SCXRcvxxs+Y0247Na4Zm9j9w6JtVVrwqlhzv3hsZHH8IqDi1wfOpSVSyCBU2TB49WAZSnaiaWj
bj/vseeea3y+0OHoZETdEs1hkVPDcIGru+zTubdwEC6JQLVzkZkZZLBIckRk9txDY9YW3BEIl0+7
TkXLXyTW7u5GQYdx8JVJjc0J2yixfeCNgjG4t5IdI/b56Nv87FWwqyG4HJe7Nc1Kc4RY839Bw87P
2edbnVfonmgUaEeQyQskfgJxSbXz4Idp+L7+0yDOzDgjOx/RTBaPxC07GPzUP+aj9n/7TTYnPZ4A
KNP4tnHX9yZtBi3k7ppYLzwIrKaqI/gpotVTrYJ9+5X01+mybXZSm3psbe4pZjxk8i4dY3lf8G4T
3M8LyfmeB3P3MU/9hZinxpZOpWc5baO4aJ2IY2jjrXPTAuudMY9bNR9PPFqRCaOKLd5WMyxDrwwp
+NkCWPQf2K8dZcwthXjfQeAgzlFblxfEAL8tpB7FvpKg70VePRjDspAw1yHOz4F832dFxnQ2tGCH
hkDv0TMBaRn1cf7yR31aAKq2bou9BbMnKYISzy0aw2OhZsqrpIWWYsWq3z6IRpi8tLwjtCRZeSVs
PkozA/rptYrOaNELwqlDp/tIFSuWrvx/sdmbOVYVmoH2VoasS+GNQaoCoq1iPJKW+TwNBWUDt6N/
vnHc2GNPOKTzMmxBl4gBN3+IYwF3ShSw9CrKRR7nFC2K7qnf5bsrA0NVK0RclvB1GrYr4eDkSYUK
0STNtpvkMse1uo44qqtJdrm69M/04jilcRFVYRFr+VuH9okBosyt4dQY/YLELkUXLDzBFGq3Uv10
YE1lbirQdIfcTq4H8COCeMXIbRzezJJ1MKu4Pef7M/UXU4VFKUwNdgHeEkXL1/HvFvI5YgWarhFB
BpA/+iDL4Ema7QIZxiuCJ2NFqRKJ9us5HDd+Mh1bdt2dIpuPYcQAl3186uDEapJyeP9jFsHT+6wF
dGmPWGEi8k8Vyr+lNS731I0aPl1PFNzfsoat3SIkoTcjD1BMWgZtkMb6ShaFBhd9+4x1Daq6144d
j1Dh493IaaCrv4UZj9hVm5rSphZiqM2PmNfy/sCoALhiis9jP5eV39h+Pt91jMW9P/+RYVNNuZw9
XcFd//jUjTl0jie+1LdagFLN8qKyJGBaYTex4WZgZIHzuAsPyR25XpEjs1A2TrlBtkHQcNupV60n
K8qNz2rCE0YfPPVjtoKkdRnDUC82NhSGZYiSuLu2aSlic++XBFARZOylUKTuWlPbn7itUBeMH7aw
BaxIFV4XG+rM9hB8mdJVFOUddoEL7fF0lSH6hVp+IVfgZWtZ21t2zRVI7i64D4G0z5eFoI/EvbYz
lncOERSpr+NggDHZhR0QPPfApfspYCgEAEEfNAl0zd0Dz/u4TT5Ow+Rg/tR2xXFdgijsHyEmr+/e
QXpL4HK8H1vYXVt7dhWVfkhqAJaJTAyydCA2KR3TL5KobmlU9ucKOan1nD0oXc8pgP7qAjXgZmUX
JkOXhj82HmsClLssHMIU15o20WR1N28a1JolXVr8vnLh/lIdQARUWURYcQFz00MLGRX/xg5ViBPK
bExDrVQd/vLDaH9T4WWs3IQbQytjQJbcS/WA5TOmiBDBKDL32m00QUX5qRUcKt7Yu6U8mOfHu7FQ
NZ1v26hzz8YZyTXFDO4SJWgF1kxc21a1xL5B9p5KT4tp7fO36nq3YTBnpcgFBdoy5riYzqiOHTWP
bMhtpn65Nqmrw55262Q9+pZSjkX6vj0XLv+LrY2n5Hv+eSEDcFUyZ6wa56bFu4s3yhGUE2if+JhZ
oGvoe88vNIyaZ7aAB7FqGzY8S8YDrr7ZDVEYbpQoEurbmfJ1no3tjngfHKrEw4LMQiNaTmULUQuB
ZCrAfQfeWBA8la2oiynyzoNvchefCbhLsM5kLpQHtJN4MzlfWibpOFGp7Cj91DrbiJgZ33OaNpUh
ZxdbvlgGFeXKhnpqGfV9CnvK/cwZk7/yVJfQ1aBtyp4PXFMh2gLTMf6t1o3A8fYClIG3MpPLq4/P
h4wML5Ituf3uCUVHzv9vsCEwHileCNgS5gCZrL8Ee6CFi4DZuJmPK8N7fb2GbRT1zEVv4u1XiVQ3
L9Bhp8Avm8ugNS6P4MUBjpkNpLM7xZLaHNOp13MojtU9iUo/TmCr0/vAhAL0fGIGyaP9C/b8d4ba
vKQyfBciDCbisZz+NnLmd9HiOeA+30Nff25S00SlsVyL+MzmB38yMSHURzbIdR0aKkx6ul4OWxHC
IWKh15AS4RE7IGqMuZiG5cyd4Fu7DKhlljzmqbh4Z4Q5AqcWO7Umtz8UWW84+RREEQ/1ft1fU4Xb
JHRMdYRruNyS4/nC0BlqzyQGGvDpXM+RZITaqw0SiwMc+hfE29Iu1JAN9WuSmuBLT/MsXy2ht3lT
ebS//VwdXXx9xEHtelatQeA0xUinjN1ZH7O6tLcdpoKp2X2LG6kbLBMEBKER72fLU0pvLDs2MsRd
PDfCQv/w0V7IqoVD3m0LtZRN7dL/ElHPqEEh+goNOHAeX3Uc/HKUn5UDYdyHMiMIl3DgHA0/Pq3l
/Z4A1yPnxVGdud4KJC5MpC4WqBV52kSf2h62HHqDouTClj21Lf+oRsIiA4F3ucEVu19IwIEdkKnh
Rurb+j8FDPrfeI7sbUIqlb+0ux4mY4j2pAuKeVKeVNB63iaDXz2ZgETM3O1tW42MughUlKKUZusa
GUUunjrbc+jzrNP7ExWd0C39bznt6i8X4RmwdM1u20+Hz9AzWpHYXsLlAfwn/lNqdAujvs+e6Umw
bFFta3p8KqqmcQCWWDNqcCZi0i1necxh4N5AhL/n3dcV/pfgrjweGEKATLwHMxT1PYovSB8nM5oM
/m5DBL8cS+iAeiD43xjx8GuXmkLgkTnN/YCkQDJIA47q7fxaXzTmYLbn6/mTbqAZDUcjTxHf7N3T
GwUClw15q5bBbTWlpL9h+hP8sTjJiGAuU6TyjbHUo0jZsii7gheYLHCmVHZMZ/ygum3nBY2OPL1S
09ujW9vwICHcE0f7Essgvl/f0Td4SBhsk3hwnjTriWx4eS1hl/ic9iNSaBXNEMTvNzxe8fK/xJ1C
KwPBluwZetfttWpCx6kC9quP61MqqKX9YLmPX3vzSmbj0L/egWOq4COrl+UnLSRRD1tPRoia2X/D
4WTW5FIYkk/lbaSvwjTXDxf5ZiQsv78+UXAi/YvF1k+WgYifENABz5Ij0Ws+i/flzyDWPrnIJRWs
uD+FoVBSP/01SnNCI8EhJKhbQUUxXkZLdz9WbvXwE4WSG/Sqkqlx8J4rWCO8LNZ7qOd91P6K0Ojc
mYPUJmwaUcU3KZ2lE9yMoBzaKMqdAt54a1YFvpQRs9M/ghfpkSOQleLssEr30HuXpHeKsZ7zSOrA
9tHSsaZPJIT0eV6M6iQJUI/dJoAkMPFWsR4uifPncyvXUB1srNuOMEMc0JCP7qhYFnC10NsSczCk
r5UlotFYIUipmc9IJY+fhGRJ6Eel4rSpqA//hzaqqgv2fjAszb59eUhghvkGzyBqwBf/84tbL9u9
d5NW1CNwf+vTeIbGCgyVKf2qHqj0az+FiOSvK3oWu/tByyvoQKq0A4hKAf37X/t8cv5+8IdCtjpO
VbWXQMnBlD4OQjgubPmBvfqcVkudjtJtEGBSaDW4MPPvl/mfSOIVQNDnwTmUDWj1EAJobosZP9RU
7BsIum9Jg4FK9Nu0VmAQS0anby/aVodGrWTVhpuekMDhdFTptE3KStLe3h0rAEBUuFL2/jHpUBrB
UO3jT0KUV4pIcHgZTVsjQsS4r5vUt1Tr6gnvDHEZyGdP9dObLDA7696OKAQi3TgeMzRcD1gZezA7
8C7Bjv5Htmta7IN1rRKFXC5UmKnzZHuDxsehTJEHbAS3j3qZKVu5TWqigLYznZsVJSOmk9IUT5LX
1l8N7GPhFx0cKywTkAuEEZ8XB0uWoRjHH6yI8Y87sH0hObEcDKfU3gOGzYMNEAmiCaRTPKo2yhf6
rqbgaAt5I730D4GSIra9OZ6G37hoUwFHKu3oHliuZWyvUqTNoc27R/X7zVyDw7CIfY2+ndmM7bDo
JNnH0Y8AsQp3fqH7bFSAaklFko/bJj7MFQEWzve972bdu0pUHz58fzWxJc9Jn1FfGqvwLcOpA8zs
2RAse/oo1KZFS95Zbj6l3BPAm0LEmmDxSVXup0efflpznnvMCBb5kTIGDF9L3q7mJCC4KbsJ90zp
ZwoftEvNgwWCF6lRfe1bc0WYNajFJUvtCpdkwcEvT2yfBJpUF8MAM/VnwcouN+yFZCL1YuQlW+P1
o8K2T2h1Ftnn2AVAQ7TSP1Q357gFc3dmR4oIZTa9f7tglwNWwp6xqerOg4PKtTFazxUfevTG0Kct
SWTp+0tLyZGuB3Z986sc+VxQ7/NHTLcFpPus5PtlrsEDv8IK3K7yM15JTRqt1/Tc2WUQ10F3Dml4
pUR+55cFTKQ1srYd7KAv8lPmwVDLC39tC8l/ExfAKIOtx0JPRxObIpcIb+Hlgus1TPzmRh2ZJy1H
U5N7/9Fzeu4DFe5gFMKBSc1SHnueSi+jxM1dW1zzoKV6LCWLjFCXsgl/I13/+MiQpxRJGbvO8j6z
S0xIQU+ZFmbe359kCeuAqqT4WnvZX3AfBm9wobaCdrj3IwFVer7BcPkP+xJSdGM9gaRVXNmPEicZ
cbWD0GwVfaRFkBJ0kifB6on/xhWZciKhXvyD4mgqRCogI7qi3yXYG2o03vhZDyLdV4bzFbWG9UDz
OLB3/C3fN8d/HmMB2bYwyD9HKOstJORcjXK3gbP36DE2nrTCeKzu+Z0KvjlsW0Be1k6qTdxg/27T
zAx2taKdj6wXaxELgs8s5O5QfomEHAygIufxwcZV1vSMUl1havt9iVbPmJ1muTeh7gez/cqnAbW4
sZRhfpjCH7GXhW0/MeLD1i2d18TSy9TTks+BGgRT0SfK6/+m5mJ5BhPlF3JkcIfiGutjBIPr4eXd
4oJq2RPXwEIp5HelRzU6fW8gZOjVVVCBEWL2kgaCAaYcwxSAScM7iBrBA7mxm+1JOmggairT1b2O
AjF353flQCXr+6jGGHKdA1IOAKrQ4vY9UVhi2VvMY1DmlwhyUwMVy5WQ5He87Y/ZBjqHzPrK4CXx
JxF1n4+FFenicyxNCDrJMVKZUAl/MTpKd9DnlUEaRqC+x/YAgsaRmSIMwIvFZyYBbaoNJdrleOAL
WWD2KU5fS8lDsCUe2FhFajKbemPcAEK5NlitBju6CyxaYsqKrkG/14yyEpO/A5ECPci8Pr4jqK40
8i+9qCFqFHft3SoaTB/Zdqcq55VN8A6QZJ/ZPwsyxSG3e0a5CIi1/L/1P+4ICk9UPYR6krPT6Uk1
NyBrxPnorKB2zb96TIpzLsygrOukbb5DyVvKw2OXLIkRNxuufbf1+4H9c+PYCYfHUWfJBzz1rp7o
kKQdwRw4/SFU/Lf7lFAflLYglZxuC1x3+jj6HPH1Bm78xxQqEEWyN6iWBPU1XqXWVjwJVZsKMLEH
f8yxXFq8ClTPzFxMKwEhCLMPv0pB0egOMqBOdJMije8H22r6U6BbBvrPECX3WbWJYkooI9gYxW5c
/Zn3RqSaDsKrWrkM1wm1ks6pxrff0CkveRKWC3AqVCQ3NMo8QBvmA9NO8vC8LKf0cPDZVReMyFgW
XqDnAR1bVX3BEgfbKnndwWtVKgQjlCfHbk1kHmsOMudpmO+gjgUnMtJK7A3vbwvRiFlNSC1IkaMD
qa7PulXc3GUYv1fCq48as7LgsP+ZWk2a4zitWA7aWMg7rHZokBBkRVsuxwN6NaOLnRJ1818NfR68
RAhOUv6eIKCGLExIgF7wU5Y3NRk1Um0sGJiEb63Mbu+KsbPdHNu5IkeUXNSER0f1knqEvACXQj2E
6S98huki3geqFNVMG2vjo6/rggm6bqsZjnhAbGaMXn7+S9cIv1xH/mv2ToihlVa2ILrYKIl0j4Ct
rgcDZcnY4WiNosBBlj5oC3QuunKIiczyKdddSfhrA4ZGjFOGKYAJG/Kf2rkrxwBOJazvUNboaCf2
dXGok8x8Jgc3yP4THndu1nmzPzUh+BGVsc78ci/tmBihGu3r6VdOweoSj26LDuPrn55stlRypFWE
qnbSfD5lfjTTQL9ETBNQO65oCHoO9+Kb5YFa2jrX5edRjQ76uY4m+Y+vSxtpPIod72hhdj20skkc
C9WtDFSnOZ1m6oZ+qlOU/WK5OVyHAt6D4dze4pkT15KvMZ8dm53jQCLjrSaqlNQL0tEb1lsMi+fo
IcSYImj+VUnUPsTHItvgy7M1DsVjBf/f/Y7u1YC96d+l1RTsqKVLYxiXpam0MSyCFY4e+LnzgXwG
aJQcGrfhMP3+caMRIBTqVrb9pR8afscX62KUr55otAWtuePjDwJ7GotQm7RWFdyfIrKY5Y1hm040
XpDjrDA16ITAdlPm7chVJCJZ156ITW/YyJDgHE5CLOp1roAli9OoodOu320yRExvMobgjjVeieOv
D6ddnp25AGBfa9ED4nMkAwoAbGncw3gcLUIX3XJV0s6VxzNJ0qG9Cmd6yOgvt6TTMWl6kFym2tAi
WiUmHIdCT7MDi8o0M2ZG/iyjQGcGJIGA3Zr+7arBXesvgH5nmToZrhnckpks9isShOq73u1JFDHm
s7q3VAjeVy8rogUIdijW7IHs8esJ1g2vC/8f7pvoqCdmqC6nDe6R9oqM5ThLlvfzlMO/HDkdtNIy
85gNzebDfI/B/uaGlfOb5GWvBJIVhcY0ljSZOuvarggz9eBa40iTtdrfrL3K8AyVAdxaeOqspKOZ
KMsMs0mu7BZqIMPn8196q1ICoBfOpz69BGEIT3O9aLkjpyVeMW+rkaYTyyhmF7Qyq9EWIuCMBRys
ZI8+d1Nj819q0bWysBVUVhA9tdonSBsHfvCLB43J0WhqwL4FfDaBDFPG2swGLt6jP8To/uHMlc9r
QCeRPlOq1sJrC/Yn3Er6reI1bM+RKg5VkDfeORO0oOenYRGEESfVTk8ke3nZN6OCDGLkkybuoJV0
N3P6qzHYCzGhQvZdTdJhl7WrI5+snYArTy5dK2taVgsNIpcqUvTOT++d7epKfer4rFGxfw/zG3xr
GjOSu8T2HuZek58UhIDip50la57j4csNWD+klwJGZdjRU8nZVupQwSDzyP085WJCFa2MTxbgowYm
lU6f9A+wmkcTAPQ973YKvMyTppsQQ9qqMEuSiTqEkRViycu/x3NAr2u11CQWnexgoqfqlfXOJwqi
iMUMzT1gjNTtDfnzDe+7uvgMDnMe3zsTT2phJVJvR7y0SNymQVTpB3A/UDrBvXWQV8rajxvwAaNi
3ipIFAuCzeQfgsmSySkSVUzWPX/Ml67TS5AoVu7iUu/PBzW/ld4j+0vRMIwrTmvToPono1yUOM0z
aV6VA27aZIK3nNXeuWp2qkrP5UfW0vgQhSwV8T4iLQzjazFy4L0/B3TfzNmhmN9tJ3Za/E+37prK
oZfrsmcEBWrvfO1h94LsDBmTlZ2Ci2dN6qDNDwssHnyY9t3PsyMHXPisjqF7UOBRjsszjJNx/nw6
s4hdmWPbDjN3gPoZsTt22fyjEMdvLd4IlL4bE3RfRxMWpoH8HDHQqjBfyP49xth2N7sVZ3eiFhg/
F06dE15j+H8zIyAQItjgdjziFG/CppcnVnA6uGfB2kuJVUG62inkybToXV1b+vs428pGWPYUHf50
eHdRqQLpFF6pQjIhOnspeZuCKK/aqKDFWR1RTc+HfhkxQO1GSEvbKwmB75UGeJQfxewPZnambZZe
ciMdDk23IhXJTemF1ILoRPYnLRg9zMBwtWtJEjxu1wUXe/FE50BXFphvLmq8B8igayE0xEZNMgGi
D9YuwnFNKCb7YvRa6OkOeoB1goMAU0uPNzig1WkxC6UwTZOOgzAzg8xSeHs/qY1vQWqaEOYi24OF
7HQvkeQtA5rgsrBNF5mAn6/WW3Is9NNTUOv6v/EnN7+Wfkwwad77+IFWD9mfPqmxJYeZ5owgczfl
xgu3TU6GLzNa7SyfCYn1VNdJ/V0N4alr85ooXqU5R8laINkPjKDolhyHPTkLsSLMwMVkunVsL8rn
3WDjK/P03Jkyrh9bem36dGhKqd3S3RS6w6VdqIlMcDgCgDZ0u2q1MF4PBBeOAPJhSIjZps1/vjh1
zQfnQYMXKqV5RrSjmX66+hxNcW4l38HLZ84oJUlZ5MTuVZES2YC9nUoLrRTtJAyjI2dqhsjoF2Qp
Qp833qj0bSKV6IXgRXxJ6EzwctR/9l9W446cn3ZX/yZYbW95shfPMSd4Ms5nIUBRIEraptZ1ww5F
3nPTx/52DubR0fK1RsXpYD7yk278OirDy+cf33+//B9RDx05gQkhH4wTHjEwaI7HU9x2N4mHCLN+
Zgk+zr8r22DQeeerspOJlTEk8ENCNqgVKCzsFu+Y3TbTR6ghqlQj4HD0H7UdMmL1PHFGysR97cK6
m2xKs0kQrZUdsSnRPkPfm0+e9JnyT9KxXJ5VyZhUf6mB7sOdhFRAt08PDDRqoLsIMWmQei3LYG/d
KLQWPjvshvXCvX+6GVpB3osrSP3TQBmG+Hg2AoZD8R8ayHQfmmHsBUdYJJlazWoG1Dxh/g1Cvd3f
wCGHsB8kOM47i3tdOuZ10LuO1gSlJysmnM8AjhgYdCzDQC5TCJY1mp322Pin9/CPCy5sNWqgb859
ojGSx+0LUv3n/DuJSmBCkp7ofYw72HBR4yqzoODxEHjL/AP0z3L3kV0tPmK+I9OZB3HcOoNWMXIY
pLbruFzj0sDSs+J4A+HOknONWcV0c0rCXO9nme5d1TyyARlqY34UYxNidVGS9B10VCDu8xVY7gPl
mloA5cH9MEC9iHryIq+U/oBwH8s/717v9TwYjdlsCmSYdrruFpVEGbWVmu/dRVPD7hXQeXWGO++d
DWqsusCcGHp47b66YgrL68P26MXPMWdn4Xnu9fPToNH71c0+QdGojuVww+pX95tUCMsENvRgPlSQ
gA/WQM4gxUktTd7jdUKE0Ak3Tqk5advOEpH66KAiJFpJa+QM557ejDUz2FJ76NO6c8Po/CRX7Uoh
LhaSnczhcIpkWnnxMhkgD9lPdqsx/XncO+5JTvake5hksmsLrP1lQqnO7wE/h0TRdhI8eR8d8UNu
/HwFUlB97HMYTX3XT06FPuEroTawEiBx61IdNSCpLlVp+Cd1XnPWu06IAqlZhPKhYXkRFZZWgxBX
zgYjsoe+AbSJ2m0TsUpu1JNFjmcc0lx7MjAe22TlGxPEBL9mYFCrvl8vjEJonU6f60Zj/u1yu2Rv
SI5QU/9GCjd5xG4BGkKThILpsYA/oR8v86Z9bidAh6zaFuJVixj/wd947SWkU67GxOcXrNTKLG0k
eHSwtLcEc/YuKyVeOb7J+LwMpAE999wEE6HzYrS2Tnd8vUOjjNn/uHSw3Y5Max2FnuW4XhRJTxHj
ufUpB+GHuCOrV479u5xZ2una0yeNWnCPu44EXtGBjOiuZrlK/DOr3zOg4i4nuqdyVAbV9eSJoDVW
4nrm8o6TLEntlIAH90cUixGMxDOk2kS0r7TGgS0FmUxjCNH86/x3GJCHYIK78hcutLBMY9amP7Qn
ug6sW6gv/DqMqhDmvv5aU1vshaCfhjxiyJqTac0ja8y9km3/UZeEo8mhUmXdOTawgVDsiW81fnah
PNFNrDW/mOz7NX8/xkQ4s8qPq5SkN/zwsJZZI/XcZ/85z2HL0CPN4eRw2ex1Iem2qGRnu0NHw9Ug
ijpQdpTAvWu3zoK1Rbd3xJr12+cNWJLujl+gbiJPLaQie1SS9hVH0nzFbB1W9Ml1GNJO4Slx25rN
rue+7X/eoWlSORjH0qvgvPUTPgqt6xaeonncJLDObGbo09OJhBkeyXUQpu+NN+VbawkyGLisfUnc
Sn2XpSYLURltqQSF6qcpxxVduNtJyCrfbdcsieRrDjo5DI9XRY3C1ke5p3LbcVEaLkZidNs3BGKp
neZj9AI7TvAk9D8QXerd4whTkFCOFjgkoX6V3YPPBNb4ruH5Wf68/bf0FEWd6Bylj7wv78eBZHZ4
QmgMLRm/oL/kf314OafbbpV0T5o2zpqP9j5r85+DmYdFy2C2HPWXY2Z+agaSDRWDi3kp8ZCL55w4
TWGF0cVAgx/1/HESX40VFJU1KtqbhZl5UuCw95bHCCn5/zcr3xLAwcEbvQq7XR3ChueNjJGTpfao
+ekadCQZu+6o8y7tbulr9TCtvLyA70TClns8i7jcdbZahtktYyngSRgGm4HnZ/5Pr1AcneBwrRvi
TG99oLbH4ASBUZ4vPt0LcI+ySIeQ8J7a7UJO7PVjHM2XsF2urD8pEd4S3eOJfMK0YeafjTxnpp0r
IzFnEaMpXWScs3cJCO/D3bmOeVVfGOSrOG1lrvEjc0HjQr+Nkq+y2dVQqXyiFa0VmZhsjTnaNsu2
vVOfubncXDraWIQ5xZKvDsU/n22qUNl5SEEFKc155wAq6zicSXxaRTSUYqMv91cRw+K1fmrI53Gi
/aYl/K3yaWm4ha8lF1nyzDZSmAWwyPK1/JIqJGTmee7wgrrjIR75LtZ7sbUhVBo3b6H4Ap534hMH
99kIJ9kbMWGtfFm3fhVDhB8+hDtc++hlgcVI3wXtp4U4IsGtwLY7NXkdZmZTmAjigMuwdWUTSjoa
iLgOgCowfsdYh0ivOBD7QfIHkJdKbLGOwmLiBUMsDm2BzDFe2NWr0HB+FMtrfnygakXiOcfKE5wv
7t2ATNnUwFZWqGtpgJpTx2Yn05QfXwN0SmasUjjrUDa9y0Mm1ZZKC2+fYlGt4bZ1YV4y+WXFeMAE
F84cLTdBnmZKfPtRpGVbGTd45t/0zlMEE/vLKvloOlu9Avt0sIqJ/42/oMJ0MrmJCKKA9we780eX
7zj4VQxANqmAJISXrXGcduPIEF1YEwFKKpPv5VXgcW0PPUr48iUGBolzHmLli0Msyu8rEqjhRdox
jNOwxhdIOg7G+S1zbe3IGyFnnkaIB8ce8uInEMVic6Ht7i6OIqlov7qn0hmSEeSapLWrQ76GRgLg
2IWyOpLc8PtkTforQGQnL7/Ewa5BRxR2kWVCI2OpUnVETp1sF2TzRHicyZ86ZruRZk5vZCNEcgHL
2Kdc1V4ceWJJn+hJrEIie/QgovXl1yS9Rjqu+YJnr0jrvEupgjf3+seq70Dt5LVTUOJ8Dh8bW2iv
FTrNAVhcSDtdf7abUIj64CRgnMc+AXM0JZ3xfPMTFy55h9N9wVKKRxHz9XdpQUjN6hYQGVf+b6wA
FRQDHhHEVPeHSeT7leixt0WgOdzZStAYyE0yZw5dim146ow+5+V2wjQmUiMHtrLpNNt5G1qZaKAV
bTDdLsoA+0SzGEaF8Q/UWYZkMEs1NlZTXWC0elWi5c38owgpMdQz0O+GJXfuR1xDO7QUt9+Y7idn
6VReq/oJPUDmOcxq19QMX9r+3rUi7iORWmhQk2IKNHpA6qtPKnR3zCjmIAcFmUA8ATjiKPJg+uJp
kA8xqld48gcnC3SkdDh0aHfj87PZezb1F1gpSreZnaz9DwVLjuurPrZF6tzhLBGpVIzb4MxetYr9
IN8BViByvkx4BjS9z5PR0sFRw4toJlVLle308dAMsJgE0vPRhx1F67eQTahq2fiGgpRQbeAkCuY1
9+TjNqaxTpl355RmKZIo3oWb9oAgwBZrkS1KaJWFS/066qVwhfmK5jgxE/tXnHIQkEzAEI/teh9G
7SxEch1s3RQtvVz2QPhBZ3XdacgmgzANqcYSy+0otF55gDRBIHJh5Ku7X+fro9wuWOTRe5EdZthU
mPsBEfbh4CPBmFVQtNwh4+ginDAGb7Nmywf8f+ClojvhezM4b+Y0DEWNzk4QAfk1cCt8FIwRj91i
Oore3U+OdO4hFuEorO65ZbWqr9EMEKXymNGhBGlBIFgAf8rrRYG1beU0/Ec7ye7gt4amdPOAoSah
oPvaO3THirUWaqKkrZYd16Hsg5TMjJl0+7FWa6m0DCRHhdP7aOsoV/Nr2I11/vscrEv/jSVAplhA
aF+RIYhTQr+0lflkGCF+VAgy4ipynDIYC6omkIOEM5pKYdc4L0H2f/p+5MMdo+YaNNgmzGq6m93M
S6RJRpRT82EtaoDmBPJwWDaEAfSm7DhocITx5V1yvy4ovraMWzFqhKJH+rhzuQZfnqQACPnp/PTo
ff1juiiS2BiaSySbDUgBsGG0IH7la2XKp5x9/vtKbBw8fewnEysJYmBGF3zPdWcHCR8h5+9s4/jt
Ixp53+Dfe2cSU7S1EtiHs1ek/lK9PyOrkhqgZbhNww1vFHYIhLCPGrly0fbaW9EwQHZfvfpKhVpR
3bQTBO2hW5FbTreZeqUbPSMUODgIZGkNBAsUgrR9ujpbtvmMAP4mvUbJWHC3u3VQMAcBHG5l54No
/+bjbehXnW77IZmi3Yf62K9k569/s6ZaDuPElgjROw8eeE9v7nh6lRbpXOyG77NoS1XWur2fBd7G
ORfH6WJ8aXII/IMjrQARym1lPAZ2eSuScNWiIg/4uMOd5X1bfizziKW+X9ng8jVomGpIDnGITJVh
sZch5jpQ7sgR8TBFbKWr/ArMrfr0lds1vEZ0qbJ7D/H1ncEJjWlj+7pZt/gsds+SkAjGSheCQIJj
LoHEXR3OcpESSqIU707Y/tW7S9jK13BaNQcnHgSpqp6+j6KQvTmCbT9udtTJZ36kbk+7Qu5VtqFe
ZNx0unHaG+8ukLb5atRhAzg0GwtNgxrwssI+WX941FFxhvuarulXBPC/Uxog84570GbRUAcmvMHU
qXD0R1a4pzk6q6gpBribxWnxpXxu2nJSDPsIwmx+T/BumGFaIfzZIHJrR9kHBU3H0ABL+YV8NEjV
ta/fo6EJzJ4LXL5U8UD/F6hOYd/8B8mzk3dtgWBV1Q3X0G3FssJn2txdqvHF5/Sq7nvNhC7jh3GF
srC4iqngKLQLF8ny0hy/bMyifjPpFSXL5tYX7ydvyPa8lMnaGJCye2zeO4OvwkRUV0oJGNurjrl9
KUDkXwU4pzGUJAz+El4vADyOT7UkNtCnN3sj/kIR3r7YngcSkpNUrWx3auqHk8xl62nqxjPFVbUw
F/Cv0JysRSe1c8hPznnnnXoxo5G41wrWzQLCdMFUzw9IgrMuCbxqu5JJ2SCLWdjEdjyG18PM2QF4
vIilr0N8JTAqSA7Kmgv8C32cDNFgoNO1HIEp2lqmC8A0ETmoT9okmH3Gde9MrbnncWRp+PV5xTlQ
YCyDsKE9hYLSPA65CN6NRMCG1d7d7NjGvnE0rF1YDvHEnAojPfDoixCSYYnZlMmmmkaDgs3kD9Yh
LW67/svgIdz1/1IVfsp27vse4bU+PBfPc8yq5VNPwXN3kyE8yrR4FA/TNMnuGFTHut7fArmFEar4
aqIsII8se3cPdoXA78a+vdOtecDTrKwLIbilS4LSKUpsjEIps/hNM8qNRE+fTvpptSgrH3sKDVCC
DfUjgcmwLgbsPO6WECq2X3UrTyrnMfWPle/JTglJ01oQQ64Bjx93OmuOK6RDb1qjtcGNbo0mC+Ow
hRVFviOwZSfKiKb4ay4Pgj2SCoo57MZYj8zFyF5XrjCE5IKnH//HZgJsg/fhOHuaB4XSAK3Dc/5F
CPVcv5YyTQtArOXamblq29ks1uMwb7J9lCEB92Fc8/wrkafQaE+sb8Ph6Joy7sbYmuyzbRdbAQVp
NrUF8CUHH/wCGt5BDTgsEEssOsG6+9LpOdratBiRXQr6/kfFOoxbjS2ihBZXpweT2GhQWXDlA4Z4
U3Bqtz0TaUZ4Q5B3Wp0CQbQ5OGdzHw0lwuvlkg5vjhvmoybGRoaXZctkI9RP3KEKoRRXXmnCkmok
vsD50bW8wJnhQaf0Llmcy8IDFmpOb86UROaZGv3lTS1nXwJ1I3oPFYIAd3GzCdX0+eh/F10nArdV
1uuGQbfUqEs65SDzR/cszGP1WJ4AgWPI7e1TYIVGMYoE31cFudfYcrwYKdPVNVXsFPqgW3GYBS9u
iQoDQKFnmwhHB7YpH42ao6d+rRbW9FlGQ7CIGUoKS2HC6vNbITKtE94QUzf7RJZiYve/TJUbTpFY
c4wMKvLYeOz+yHWQd3GZrRbAkMLKTD7Jko6vJ4rqccuqx1cQour/oNBXcveT0pkCD/kcbNh76YZl
tDhqunH7nBHesV/zj/c5RdbM+WgD32+Jr9ScBuX9mwgTVE8LC2pFcSXVBk3gtBWg+JDNBzb9MCef
Bb3bBvJ1EdbHS7cO4SUQUu1ftPFMP38R8bQkO3C/4OzRA46D/cp+Mz1QkCLDi4dPs/o5bryd3XuA
4Qfk7ZzNsPzU5nfRADCRX8viGj+qe1xWcjOTsRadNb+CbBZsM0QGLlhJEe8pBz+KITjjbJRsR61F
+1IpHHtWTATgbtZCzbMXc2eHu/dJJQPGCHHQOtYb3B0LWEUiP4OxwXD11lYzdvA5GS02WFoDaCPv
3zAOU+ctbZkFQ+fDZ+Ulsa6JUbgOleg1AqN6JmeGbialBIWo+1FLT0+R2KSvW6IDROKWZ96psYUO
xhBGoHBzy2Z8CtIrV3ds13wfaU6eSFLsk3y8sSPSVAflmmdeitP5j12W2Q1VTRob+yzG33PCKkCe
pL7/QYy4i1GSCQdqy9k9sviRokod1JmOQIhGIVBWsru7OKdEtX6q98e2OnC8+mM0GVNO8b4o75oU
9FpxUQ6a9BKR5n07FTPgTgR0hVOqvw8EJ40ZMUT5XfAjq0Wy1fimWBaRHzq1k8hRp59UcEhhK5Xr
9Ui5YaaDVN/L/82sqB1rHMJG6zP54eJMYIbccsk17a16p9lwUzLcC3Qbf+A1k343BUhj8zsOZS6r
2r6Lo4adh3qCHzF359ESLJUytoq/M2R0A1brUXct7gU2g0bViiExYPS+fWn4q9waNirG/8L60Ob4
FiAHQtrjqMPf2eOAkeNpVjk7oMJEBA+p9rrBy8Tr2cRT5xuCnJsw0Z6eDG8KOUlji7PI/JLHPFgQ
vbJVfi19Tp0D13VV5rQ+Dkp+neT0n3ZNHA4x6aCpgldinUdpPi1pYTMNRx+A5v+QT4O67bfk5zu/
bWcYuGPJoQssHbHUKq8KmYCzT2NZHcYuU4Xi4YmAvtIJ3ngEpyloKCHvARFwTj9u/KS6Orbmxp5P
zdxcn8vH5HgQHrlcV8quXQhK62A4ILdNEqpMo+lAe0GoRmv/9dVVq57rsUSQN8wz0RgLRXvA9nzI
FG9nIUvke4RET6DXJXluUkrlNLMTKLFm23nK8N8CCMwETfHCLC44FbG8apggVoq3uTeWVQZfwJPh
H+ZDidCq77jkjAMNGIPgQcsNIWJsFYGJkzp32QRjAsdZVc8JvWgabe4NMZuaZEovyzJxYvbnczQx
eZ/avKCH7LPUT621QRsMv546AW2cR6oxwVANRt1Vm34h2GuDfxWfmTWCiSwRMAqjYZvik7+Qvk8i
b/dUgvVVMrXK4XOlFHSHsWQMv9r0Lfe0baFXOn7/GgQ2JoDlKaZH+seTF6vq1GupO08h795uACdw
csbD6FKf+GwcceSHUctiFIQziGOZ1RERicUhm1eJhPeRNW7pFAhU0XScIZysNv5FQrQfKp/zG4mk
DeER9CYJBVqmTsPT7p53p/1SxQ1UkLPc367Ei83lHpAQnQ8hX0uFPmkdvO9frtk5H0pprIHF2JUG
LCNY3oX0cUpXuev7/q07d8gmPjC5/yOeN0WovlbTxReFsfUywjPVXxAyME0LLAQ13KwyK0JHECtT
9fnDXbtMNjQ+pVW/YxpPrWYKsp985XVYuMIsjHkN5rA8kP9JFk8z2Ch8z06cAVCpBiCbd3unMClW
fIa1pxcdgtpGyoKIB21apg4KLhX33Bv4jSfNo5XbJGvAEaLH7W4TkF53TCOlhFf9WP6/s+5Ray4+
vwuxvuZHGk7UC6RqpHKD1ny6VQ6eMmT4NM/zCt743uoj6JHlm1FFzt6V/VfOkk+k7aGUpcZTHuec
YuVFdGXpWtHoFmvjo8GQdav6XAzk6TG5qKXsFvquKwkMH4zJ/OPVRysHrKG77Tsy+Kz1b0EYrw1a
z7qDvJGG549J9Xts9MzQtxWhhnj2NXZdNX5PEqVl/cGDJsOruGSdyCzxlOdWmnN0u0NQ1CORM6gb
7+DLszYmVfvCsAZ8q+btQE5E843pESkKo4BMFWdZeL1bY2I481tm7iJGFw+A2Ahxv15h2ihXPg0R
GLzTyYW2Pk4mF5fzp8dcXGF5Td01RQ7EDljUOAEDowtySHHPEMqJ8DdSLwrEAfBQxfCF7bO2VN/p
9rHdtFzgS0epDZIXrSxMv07wiRwPQFKRu9P3tpv6pOfzFJmrv5gItmzrVp6ol8F+glpGdXflAQFD
4np79LyhXaw0WUJL19ISK1WRbnygfdvQSIp3kkt9iMVVg8Mg7XZ4YpEQHw75SnuiTi0fOZ5ZgasC
o4B1EeIuurmHZd6Uy/IkUfJzTUqk7SYVahj6onS7I5Is0JsO57fU8tINYpV4LqCsVhHfw7RfIdEF
oEt+v0QSUwS6W7uIy4vvtqBrAn0KZ9BdeA13ybQoNuA+960Ay6DMuRc7OzeeoInpPnKeplNLWHwG
T0yv3MCri3fhg6KH62cy7NW3U7DsA2KTqLSRMno2MthFhMuqAxhxrNUCur2k0fEs/cadbTxZgUSW
jfcglqjsFf6ooA5dtvUd3nhZs8JoaFna1KM2iEQd/A1XBRx2Fh71xEWjlJSiuA1waChCJ06F7XQO
E5NmRT7jSlj9g9fmwrrIOb210pomq3rrCZ7cM0EXcFGyF1AZJOGu2Jm/oGrXiP7+3+24jMFz8Hb8
t2LPiNhQcnPtmLapze4HdvixMctu8l+fr+WZDSP2rxBwTghB1P4BOffPITzyHXyCu3ruN8Gm8p1R
Q1HTBfgB8HIXUk7t7N4MTX0m99QIoAWVkg4e4kERqcrAU4dPh0Q50mBA9rH8E5EwO42NvLokasET
ceqq3No7daynUS7RziUjKOlj4dtlDhI2zfnxA8XSkgRjTPeHcjCmxyK1cH4nr7swZGOWkFNVw6kb
caYqiCnwOqxlY2clS86u+f2SojoYNWDLKKMek5xMMSAsTcqgeJ8OyV2sNIVNmt2gj4VpWGrWqyhV
lEmkU0bd+JenVHKxQya/2Sq/dvDd9mD2yykV+3NcJ3t5cb9b8O/Pz8zYro3dG1ePX+/FXZZTO8/t
mO4KSBaAEB069peQ0dVwDbz2B/h0Kj1UNGvC3V14eWhbKjIHmmGdZMEfT1oDlrFYeBiQOuqO1aWY
K6cGcJC4Wxk/B9g8pZl9VoO+eu5KEgE8tmMAkECJEKEdkw+1Pkb3w9HK5TrGegEUZbKUDZPqlfoi
xZdv2YxZ376UwzIgSln1y9igXmvFCVd+l6YPkNtUf6iJvcjX6M7w+srokVRYq2yasiWROVsmV+fB
majaCRM5tuNueT/xP4vmeL6y/yHcPCNHOZp6tyYbMJnVu88JZr0Sv0DXeb3VTeHKafqUrloRFxQT
WRbrV+5Prl+7A1/xcwzzHT4Yp7WXotY/uH/OX7jgpTdK3vzG4J833OiEcgf1xJZ6z/BDFSBtg7rR
1Muau6/v0kMtWuHdWmBSzm7TXWxRynd1tXEv/rX07doCBXWZWz1PuHX4yfWHGYCf7A243M4byveU
kC7iFWtMRh03Rz5bPAfli4IjL53S2cS7vIrcfVTzOADb+RUJvNYSq17u6XuJzkZj9j8odIFMOT7Y
VMo7Ik6jOt9NElL2/RyE221dHflMxZK2EOsTEY8HG6mnecDit2yt75aDzfmgMG3r5Zry43OSwic+
ViSKOoXh9CY079qm8dpJ3MnDyEGOaWp82smXWi8HAFIiya9pvlc+kU1oAHgDxcSA2pmY5W42zpUv
nUU3MUfSa534TWf00pcv44QsY6sWl0gn1S1Q59xqSJw/EtWuYFAmteC3w5X4JoU8NgD5xt9QG5lS
zBxhJALBZY/odkfn2Ewo5+1kDWIHqkXqGXHAVA8OYktS8GCDxYxpFSA23y31SFGm4M21dtLKvokh
VxasScYY1i2464ZXRQGF7iNdGiE1vPwILnC0Trek7FTWglAuO+rss5vNIptfitoaeBAS14tHnfLI
IttogaqMfkW/70Q1LJ0hvG1ZjdcdPf+qNpkjfbmKbSC2O4tN/+OEEWconi9FqqJRNan2wZtkQccU
wFy9umG9r28MNqKz8lO/6jC7iCp6qEm5xGY3cZM6f0M8rXgL1NJBfR+PKnCxspEr4sTNOkQ4Ffn+
4I7lI1x2FQ7rQVcOqnZFfC+e9vYwEizcCltS4z/LNq39DOwNAnEZ98Fm/dn2CYB1dgF9G9xNXHjW
0WRvACbHGZ7XxYu9HWbTvaVow8UPuOQ0bvvxN8gWHaa+N2Rmj09fhO4L5mB/d953rgTIiJYw/Dct
FWliK6MZOGyVDC7CWCGm8mH5o9MQTiqEPNW6RJJMxDQq3hiFdhdpq1+BpRzvRC36xN15nmoxkeG7
6YaOXPjJHwgpQeeIZK4EIVapYmvjO+sR/IyUsJN6nprGSYFMU8QuwtODp6GctnrZfNdqeV4U2taI
O/+xYSuyIl8fsusiwMghk+TFR0FEuM6OoOndkhedOG5E9lvCl2AdHXdwFUgV08FBN8KdUWej9feT
/cunA6f2/jK0BFn9y/zyK04JE76lHnGw/v5elr6Mh+xWjtOdpmMqHSKeoO58naooR90ieEaJ+SA8
KPHNKB/p3lcrfJNyn45y2wVq9L8iB/1NpEZUtc+8MDp06vwKnaTHEvEB5qXXcvJp0+lsSS16Vkry
9NRkI3HWc6MfHwv52bv9Hw4pFvaeFxZ26CVYqmTDN1P98/CmxdWQdnc6xcftW+GBGYitrHSGR5ms
kXaNV23C8eCa7oNEtXYNJOcbN8R4HVpD8sn1qYMsTO2BVH2ys4LKJWfrwpfdrDn1l/41xBDbxKp8
37PhWET1NMgbJKAlflVT8mcEySxXK/hLCKN6ndCCE+lIKXnxy+AC41N7moCSmpcyKFC9s+Ci8/Ao
K0OtLGpwsRQfwcn5LdW3/2iAUmxpkl+TA4++Tt3Z1qbYsW4IBDYU0ItZPJWkin/lMwKNa0H1iFPp
T6U08+tYS0qHfugbMKh2bt8UYUxfQzgCHFHrjq2RNIvpBZ3T/RSyfGHTxhtnL6MzqqKMIDiRiDIW
rtUxhDsCoz/D87fmbC+v9OqLydiUJY0NfbVwrUH7+Sb6QgyVUDN3LuZEYW+xmTfXLdwS00n7J+JL
CTmIwi9v7oNIoWyYoNGezz6KoQAmqIqap0uNfSGnkLvOZs1ceCHW1G4XIGKtjRcouNtszWOUQthi
VVwmwccRePbZ4yJBiPN7Eq7bHyd+TH8uRMUbYJ4E+usLhlqeznvJDTQve/NV8DZweUC71ENRXZWQ
sK/Q9JIuRzuS0qUPL2IvtAuk1fVhOYcbWO8duRGidAEUPoio08GMEgKKK7ErVmS4Nww9oz2TGvru
+G5JtLP8UUyxZesEGcURvxbYRYEhVCtLiSurQjbIXxuox0dUWKupgbcZPVzqP5EOSQeHLQcmW7Cc
vjv09O5F9kwm1VcYhCZP4I28V9bDtrk/7nD23wLfJhmo7mOi9WgTn0yQrUyppNOFItnUU9yV61io
OP9RMwXrB1hv8Oaith7FcExZTQSeFJKwdLje/mOcogEdX7+ZpHwKrP34DYWxeX4O9CR1Orq3bAB2
b9g5o0qYXnC1fTMzVOurwi6cPw0Ib+yJAteMvesn8kr/H0GWvrZeYR3kfszmUXVMD8DQmMTs1Oal
wSvZdE2WG3/sG6YI4rYqSsObASCPBrtxFgtKust07eRTG+tibZrTLDAwoWJkfpzClQIJ/5lMHgna
5S5HOtvol5DP76kB0c/7JmDRj/4Bi89pkzwly3mEdxYf58/0dkSuKH5Jhp4h2oWjgGEMAYY1Fyyb
vrMvjdA9s2V14+rFWspMAUiJJcnKsUCde2+2pbxkqMfviCLfBMDfGDIaN2rM/Voy14wJwPwcM29t
rNR4FU5Kwq1WpAqB1ohv6RhlTlrJ+B8YZVJG8AV7RhBDqHP5EvL6K+Lv4RA8rpzByGT58Pjka68+
YjziCvy/5orei+G36B3nsSFAwuoTkDVLhJ54uzbaBDB/NggeZnnGIUg195bjbe9Afuwqj8p8Cvds
ESiipn80kWA93y6bmeFjBCUY2S75EdHMU9lES1vMb/lNYF2ek+50palKo3B1jypOk9/13zjSCbwQ
vfWJCZNVYMBx+huIWrYZInFx1GoLs/MA44JdLjtHLO2Sow2ZfNpWy0Qg5Qj1VRTrUyHFBXhKI7Bw
OR48hO24miR5PkO49BfF7UYXP3t1gM4qoyUxBJM3enAhD4X9sQpFR+88jSuNcgWEvpCyvfSdiOoD
XhEb0kj0xw2y5pqVKtJLF3enSUM/p9wOa3CYSxDYwWXeJa4KT1w3SjqfQn8/IeUw/RxEj5R6Go2V
Mxgw2/qY3Tko0+HVhGLdyj/ViOCEuwMmEorRL8Ii5IwnM++CMB4Qwb54NPJT2USxiOZHU1NUpGcE
FtfIfSpEqbj5KJs/msOfddollZmFO/Ch156WpUaKCER/hx0hBTlUnxxA3iZY5FzYI26AhX0LZUI/
mB2y1VxYYBIpSC5h2uS/K3WI4ZuSUzquuPdNzj0mimwYQU62TaFPLpf+sI0g9m3zrHnaOt8CCQbl
EIjgLhcm+wigE94PiLK10fkN0lq4iH1L8OcGHYkE6w8tL/b4CeObbiqW+6wqjvWBUKUyAtOx9wTO
YxAq+KFBt7uhe+6TR041u0xTniOeD2iIpvvTcfWpEmgQ3DhfcyXBYIVT12snMye0jMzbtt5eZucn
v3e0URvSJVTq/zwGMKJy9qRmNd2SpbjEpFP+zkshxTcXUzTHP1UJgoU3aPpEVySSZiUBAmFYNXHl
2Wag9iAm3SdlARwWt7d/tZoyc3CTfkJGWNfXDnYGIfaonrgUUV+uqPmV0l5RShH9icX2Pgs3JNbo
mxgI689dsHQtgDwPc4nkT4ZwI/eHdv1XqI95s4BpyZpij4M+DrQd7z3NrHHReeLvOvepgqx6pgs6
f0x5ORgo74h4Glb0EJmpT0gJaOt16+czOv9wx3QAxWMDyZ5KLcte68IfROXe8xWDUIx1m09+aRo/
rv0MEHrhjplZA9CpCq/G5bagHhbUiIqN9M99+G7J7vTkgM79LOIpbH5xKF00mPGWva9ScLtcp4rw
GClCMmYhtpm2/ynIoo6tLog3M7f03pHu+9q+zg/9dpburrylmxS2pj6m3DZvwIWSYIlR4/zefC+Z
hHSPcFzHSM3EElMWh04q/c3PImA+tM0jXEpPuQREhAIEnJ3RzHKQsp69smVfquB5WXRvz2mL1A91
2UT1+3Lf4bmq4ydZ/TfyANS3o6sL6N9DHma0UmIABQeJuysiWTqJpJokm8I8pH12GlrASuXdMOxU
KE9k3RLWU1rtiEG244Hwl36D/CEdlmZidIgvWEhhkQnd4vjC1e7JQRM/X+Y+YU//oVDaliFXhKdv
APGgTul0F8FxfPtYWn9uJM5Zrb+z803w/K911IY+9dK7Zk7rqdS3sV1Ypjp3q7tN+QmvMV9jpsOu
s5Lbv9CL9VNjZgmhtkqhwA98fpKBMwgcNJl/4IYJVLAR9Zk2EWn/VhNA8diW3wpfn/0GbrTXZPFX
9meng1pTgJYdBifskOT0K4k7OWO4AFqsG1GS7VMea5L26nB8a9/MbgtDdzg1iPd6URr+XWz5ocS2
XHBKQswv+HsRY4RCHdgVhLCI8gQobzN86lYzSE27Lac+pU5E7Ctdfqkk+jKjt/dZTT+Vb0W/emqq
9CYJWin0dWF3kbPH+Ken0eSnUyBBVVPpUi9oNEiqomXzu9cGLQF5aeuYVomzjJNaNbCmlRRZdct6
qZb6NR6jMoXiqcHIcWj3yik33HzN+xevCc2wF7jBhQjPCU1+J4kOydh6tO3ceyVm3+F8TkWtreoF
6zIuwyc43GZboDkQsOTYsDge/D2lLipeoUjTUzonEUJ28pPK7JDHKAy40hvOWFhpdG0hhx/2yf31
8B1b2X6Fe3shoo8whrHNwY4WSwK/nLX3AlfxspPsygsWOKY20j2nLLq/hzQGsyggPGYEfUiYczpY
o73ZVzRC+JjKzpBiXUG7U//xgyXurXclyRUgUhcS/IJ3+y0uOUSbEnZPx2QsYGxC0FSZ/+f1WLaD
EMLUWy/BaxbiPXDH5OU+p6RylP2hXoxph9d5+JfzVifPfeKA/giB7RBQoPDEmvy0wmWHx2AzGF3F
TdZ7msvTIPbrqMw9kVkw3KAmoqrqdrEAQJJKjkFyMxiaXsgK8+gSjhVfM3TbN/uco/xfKqWZ677Z
xGYflwEzZ2vAAvATZ+1uKeI/oaraGHEbqtSkqPXExiV3Y01Otg+XJPuX0akKqRblho5gIM22NwEF
ON92GZ+7UJ6FONTX5lYXh6sQTJZ1rpAyZ12sddyhTbg615M8bfEmHr7cxHhDe0cnqar4WVXXJZrM
TqPM0Zqqqgp5R0eksTnfwCOcWEjvvHs/37oMESeyJMFLq08tuSlfOepjR+37HU4+Y1Ioz8aAhLUD
w4WvsQYRHFFAKNU3noNgbeWKS48fFFHw9SX4TzHlnnXFLOe0VBjgH8ODyqqjFdAANlh4LwDwJluu
y32cBGqMfeWOTmUOdeonFr4A4Hg64wCWL8bg22+8N04lyf76U9y7WOwN1SwikrWh6LIPWur/m/V4
fuiOgme1sa6wr9sSdTrK2R4E3s1lIOYYcYd5ZdtXCuffGTdntVhB9kxguVyuofs1VONVQwoUp202
m3SfJhlXo+PI6DZ2YDg8WE6NkUSnQdtbCq2LxLeucotb4mnGEA8Pi/MI6/XPtwUnIsj7ohycePs9
5SeulsLWY2dpTh3LSx/dSI1ftjZ9HjqTRni/o4hgvU8i8auCb/Z0GGDij05IV30SA9/ZGyidjB6p
ZcNYqeNp0HUAjOS82rYf76C8XGO3/0CMyI4ITPtZUGLGFjy59s9H5fy31XLjbWK4wD9bLuuITMZC
DbLxV58hLVWdvoOcdVqMj2JxAHuiJohDcZbaFsow1QLtzbPUAIXPSUjnD1RLwEJZXA84UApZHwm1
cZi8G6V+invvdwrlnp2TkmIdpm9O4w8JMgfuN+szlPUmqvKYQnVmMPIU3Hl4FecxPwrnoEBwZdAi
YvRrlLDcmXUDMF0ZIfcyLbDnreZSA4xsfj5ARd5Jl+x5iiKQz67QOVczJGtcjB5breUm7afagJKy
Sc4kWhc7B9YXwL/imb0meI1z6ugWUPrHcbOcUeQnlBu6QUpOOnr1mLQXIZ3KNvSIqn6gQQlTHMup
cfnRXOLQ6HmJTknLdraXOuPUcTw+sSmSJwcUCrpQK1ruSiaOdpAc3mPhhVTPINBLmj/MjqOBcJjC
XP8bUSmThXSzO8NpAn77RaLVBl9jfdcYzaG+472q2t60lrt8G/etsx+0jzr0xgIsNK8vHJGvMGce
WRkL5HYFs3V2o0PARx3epYDl/T/IUb9gS72LXcfoT3MGmN+GA2Tz5fAvgzrnApTnIFUwhi5XzAbS
xVro1WoZ8R35Ke2XPLtnlIslCCAflTM0dF/BcujcxGkT+88+qbNFxN8GFLViijyrszMgIAnzbcqF
x551d1dtXOP51Mj8AiD6JlPBdH8hh7wYerO04Q+LKU/elN8G+we67zHHTCxiqy7LBQFTtybLjI2K
wCuC/2yyw8IcCevohIKBc6j7v5HxAkqt7UweIRqJvoC/2hGFaINT6S2T8MoltTm+6szWbNLVy1wl
hK385414rrKwEUFTf5GEiehwwNC24zQGRBIjoLMhEZS0hJJ+XemwBKPrg2giLAzw2E8DLAknZSy/
nG5owrkk4iKFL+G3HfZOqCRsUpl04mjjoFHT/3hUP8pakGv6uxij6wdebkwIfMWUlqGEflnGE6I6
suRJf2yhZyehMKV9/9D0R5oCDQv1E6JozFY8WF6wDs4QZURT8Gk25iW761YkL1To47JADKcs1V9v
fTYrBNzOwnTP5u88FRhwpH8ZK74zx6cKQE4DwbvhbwTWjAVYV3PuHnp5eRxvOR5OgR80cbZrws23
mF/ncfZ40EPzL54jkinajLFB5y+Ieo0hIM+8fLPC06TC89opKatFPUTm1SBdY1pFcC2drWeiKmdu
dhPpRIouicLvJTt2CQirv5+E/lAh6Mon91d0F1/cW2WhXleeVMQwuHtmCX/pXVv8mJ8IuJvHsAvl
b7W2nitSHE0if2bNVNGN9o6UolYJMWJAee4D5+HP5JoJttWYaRKsAfUq53xMOF6FrMitg9mErolB
X3wibNynBpZKqhD5ohk+SJaCAnyn/qCA08oNSpZwNxlPCJRJlkoU/KQMANtfVvvZBP0PI2y87u9d
bNuEadhIW3qkDKW0OpIKHXL3O5zELgFJCjIwX+tncfvcWYRbbLVE3NNxG2n6serolpiYRVkJup2F
aTDjF3FZyoCLbBGHwp3QQPPjc/zQUlsLd3xKHenzt/c8q4DOY2W2u4b4ipZxc/0CmUPq6p1Ccc6T
D5HG+PuuqOPrMuvrkVVDn36jLtkBb9Cv0eDB+C4U6znyjLg4GRrtSc4aUFOEw1eqYlXaZSEr41WY
hMljSaDvZ73H4CyLVQPRn/rk8KxWx8Y4OBZZNIE68Z+lA3i49sDYgShRM/Ld02NPld6d931+bxDY
jJFAzKDW0XkvrL8OodAmwQ4McPuAQlU1wVKrYprdx8mx8HVYyj9SnEf28q5Kz2o2WlkwQk/MJYTu
d0i+DqOxZhqzY45K3yz+gezKROvbgZgwMoz88bjsgUlRsF/8a3IuczFByDrirVrOjNMy1xRyXnfP
2BxqJ33cfEJB7/MEzZggPd5+RPRUufKajQXmECtFTwBM3r+w7HTGjXkY66T/zRGcJg+U9PKZhCWd
3l1DPIHGJBSw0MctcRtIHiA/hrRWfKSm1Tashm1Hrw2novvBwLhiws1X8LJ+vwvQNHLVySoNtTyd
Df9lp49dRhYSMFh/+bdCTY+Zs6kqQSEvZ9JkF5ZcB+4lm5p3G+PNCD/ul0e8j8nhx+Bki0SG/Q4Z
HPVstjU6Jv24B4W2647jEmGKaj3mGbgUvwHgZHwQWJAfUclZuQELyB5dgaFRF/Hes3zHyEh/CZcF
M9pzficO/WsSfBh2I3v4A0nBr77qlNQ2L3MHoPmujKTHTwOnie12WAVD7Uf3pvL2vKSTEdkS9A/t
RA5+qVmm4VKfjMG6Yl4sB0/+n620Bq7FUQQiYtil2TKCxsvki0SlfKjFGIqOUij5Ml4+tjx6CktU
LEAW5BuWJUJFlLT/AW77/H20vlSVb7uf5/NkjD9kAQGClSdKYw7WlKuL3Gi9502QmMKeb0CrrkoO
pHRE2W1BWMBjAVb4TS0Qltxc4JGU2L9/k1zcqWmrt7mX7yIBs/Oq35IAYeJK7+Gp6UggQoxewPQr
qtAebb5Zs3qb/Ps4cioeBgphRcHA76DZjqOSdlTrrYrMKWZrymAeMFE16ImtMUHS/8ibmjikpT07
YdDv5gh4DWD1wa6i18yxCTBBYdHVtCAUIV8AdOMVcoiYOUY/1Il7ySicVGSNOrkh5kQ7h9DbTkqO
z6AYbxv5AthQw/s1O1PdNNJ3lm0P2svMClml2WiurSQ2sA/JTwidEsO6iSDFxslF64mRSibmkgDo
+qr4o/EwjzvbHMcLxdwTAPigA7BzZ4oOND84DcdmI9v1GHVyy2psfHVdLQDQPU8bPSnMZ1BwhgRV
FDqzKIf0pUHAUh8MBfK8th+ijreRsz9HM5dIYQU0cxSrVvaidnBQa5BXjV2sKYRtLfdjZ2TslB3A
klSr42GM4JczNZNTTKHvH2WSmVUSEeozHSSSVC8HVecNv+pdKkTGosWdMXTEBQ72OsJyse7T4nNp
Crl0SJ4YtHkno4VTGHU1st/x7pts3cpfRW9GosLJeDcgPDr+tzvb9XXZJL6e1Az1q/dZLCngsAmq
xa81W04bK3qDZyi8JpX46LJpGSbqDk5pcHjsrT8IGEbuy1hVjCNIw+t7iAjkwWNpz7a0HfKkGLP1
m7ilhQI63hgQMhzd4k0tYYuYksHHGEflZvc/+CBLOA+ghd1MKt5Ngh2lmwJpyU92hbPe4VQQ1Hzq
0SKKBZL2GTigiOZkTzRXu3nE+Nbg17iQNrqAC1AkVGwFXD2g4mmnHkh9iSyWgwfPhIxguX1Gd8eR
yH15ajJIlHWdGZv6ofZgjk9HdwsSSdHQ20Z8i4dxYLkDyNLtKvLF7iN24YOZhg0KYQh2Pu7DEF/y
8yIjh/Xf3PdOtWdq3cf8nVL80KxIA6/wRo2b1Z74UF8OHo51HEXkcPFJzdi5h8RkdBpo6pgCKYvC
ESWoJR+48pkR8dP+VFuRj2WPuzoXMxAJ08qcmlgUXwZpDZBKPVUbuW+aqxWpWT13sgeXntV37Fja
/vk5EV+Ee/MpVqb4QJPjk2GyIj7LHZClKvvg8RuPGW8oSSzqmmTZXVREXJ7YDwNzINBuklmaTvlT
VNiuEMMTPLU0OX+nlbGLARNvgpBAa/c17EgncIxayT96HnZy76KCOO8EjeCNL1WMWUfDlNwDW2gh
AiNhikBkAv5BpBdIg4A58Qyx+rAX6aP6IP+vnVjA0BeAag0gP8+5X6HvE7aKUx0RMmIUupxRhuD8
D4nD6FbjspJ0YKEHZevpZcwxHD6U/YbyGgC0LwWSBY1Dk1QbG/3B9NK7AZBfGWVXUUb3QHcBCOdJ
SGm3Qj2HNs2AwzujwOFdSKgpy7o0RDQuBVmj4tzarl/zKwN9GEeSaDh3moOzjj7V+WHrFJearQfS
iq/Krt48CJusXCCYMAAN/n9kL5jduJyqlr+UdK3EA9hivLcShcDBXdHUjPyYx12uaYabaCC8DEGn
8VXlHzEWk3nVZg8F1G+ZvG6ZEt0XaIv08koxT+r8dOnNipSoexxIIIzdeNfar6vNiw5JwnDGSXlu
BhSFTPmEnk2h7fGXv5NQaI+leD0Rsxxx/dA7O4hYCylgg1Wg7O+zrALuOSCxXvd/hxJSz0kmzWjM
NLieZBbAp6oexPfzVPKvJdxsBlhfRs0DZKjpP2lfL1ur6p53Hix24WTG/9sjU7tAK7yFNXJamcl5
KculsBTbuubIZX+K052J64ZrXQhbIPaD1Z4x7tSZeDkVOrF17kC5lQjlgASjve+YG2a3eTltfxk/
ujKlZRmsJviE1vpfOROIsR4Bn9TTPBFg0bcYppEbOpjQAmEPF6wrnPKh7D5DbPZa+IZqPl2Amre5
w2Ws+4B9hjK7AYkIOW5a5jJDauENPMHot5bDlEgf0kYygoDgmrMQ4iCsWnTzep/DfN5JCSVxfYdP
WfVcJRYUJc5mY9OcIYfGkiQ4rFn1BFgRDjVYgm2ofMyQ6ntx8Bne1VmJc3Ap+zw4bBtMxKKo2XFl
FR2Bcq4IxQHEENP9kzZ08UFbl8p51mPJ8gyeh1T0uOBRHOFkl5j/O0LSdi+3bocsjJt6srzrL5sH
CGUdZ2tl+Fx1OsoM3IaE9OdbovKyqVn/QYDJuyBU/AZywD5Ya4vq5suW6MzAHK5999yLon+YOR7g
zrSR6MnGZX25/2IUrwnRe/i0xk1TgEoXqFtFb+MvHN/GkvOl3/kiicKhV5hQU0d1XtSXez2rSlT5
Yo5LH9VXaitWIBnEngO++8Ts/EB4/iTnbtYvhoASL7Y4Xnv92ABImASqIjk6t0BK+CIcnZHBt4iP
hMQ7So/KwaLRhVYQsgMnb8Es03yXaJhwqdnkILTRL+h9OPcKTG0JNpf9TLB+HAbJZfjGYUz+2xd+
Lyero+ueBKpJOVboNFVF3+0LkAA0x5OnbxWj3wFn6+J4XM7bZbAyIuK6WnOPLzRmm2IHZozRzbcD
pA5mGul3jkfexx4MuH6v9/fan3NKknoZzUxRlT5Hb1XxQVq/Mf9GkVWeesP1KloJsWIa/bUZYwuB
Zb9aMskAdV88h7r2XB/+SVo/6IqBe16mtF5mGzP9OGUpw7IZLLBc/xsiQcBdRSsXFG1sRDVRRi7C
bF5yWgczhQxGBc8sfQ7zATnpoRQa+oXHswOnXrpeY97YM6ai3Bz9pg2POwI6LbYkE0Wb0rkmnWcg
4MHPHIqpEnQKdVS5r3rxUwLgj3slTzxPIZ5PDEKT9l8Hx4I65sINJrQV0kFtpfKZVou4seCstOAt
bC7KBbxc8qoIZsTe/u6+yInYDappljnKn8xZK1b4x5wZPqjLEoXi0CjBJV77OS7B/R7PblRMGkOq
QfjbCaFA7ncq4TDHaQbcRgjQFNmAMQ8IJuFoXX9JgUc18jlSxtUJrz8b1CoPLahQYI/ppKn/fSTE
HPIeEwlfCLpyEfrM13lgWxkDm8pAStwXmbeg2hF6oxuidcViw5PpbHR35QTldlQN2mJutMgRwLcj
6wqTvNoIDwfSak51cHPa1xoIK4g7vVrKN5D0lYrbEWrd5vWR7haKU1sRd/6j3aDGjVTmW8Fz6SgX
Jvs8x/tk5DBXXNZzS0vmBYIJcOWNTSjEDKIkUnGp5rfQ3NsRZps5au9AnxJNdfVzTQGRntYk51zF
HQsdD48zjeYzIxihVgk3yzYkNsKQ1DCPrbX2IRBISy8yWbTQUyD7xtYsa2jlHY5/0NdF0xRY4GqJ
HRI0UXb5HkbdSZ798/O0db8poDc4ZVogIvo47my+1SzoiRw2CtC5x0tkmkCxmNnJRJqncakQhfJM
66EkuBF1TcYPw4FIkHJ6kPLTnxtmyrQYPBPczaM330Fxvs7GTszVgS5RpDpdgc2cemJ/lxHfgiJU
h9N8t4zv5qRzIbwVmYWh78f/nQJjUPtpHT/jt626I99QOirDeuOcg2qfA3ux0QKjxedki7ifJYLB
ZasgZGhHlBoxJ/KCzuuhZ3N+U/fIvAv1l2EhYR9YMXCwW0rTE/U2x82E67WgFtMQsdvEoUkoTpqy
5Nckdaqf1hjlcJiOwvs/XhFj1/QaQoSnZrKTH421NmHkpgOWkZzC1IfABC+xgOOOB7xBDUTzXeg6
IRjOwaa258mVQR55fkgy7O/mpa72DdVHfcjV5RSuO7AaO4srEeqVA9eUkqRGCG9NQLbJ/MxiS5Os
YvgXxRaxVUsT3c3/NBPJboAxH2j5MX0B0imJGCqj1SxgOlbBJsbOJHrlZQ3SsigdhjlMaqZiK6c2
6g4XEGZQQLmQHfO3sHqQhtigKxw+lgjU2kCNVQI21kNA5EXrk9BenuWRu5OMWBs5JFy0gutvm+dR
HWMvA7tqSiL0asMMgK8wsELW/4ojCjzzwEeonSdvJnXIIh+madtNfOtbHnJv5o0Iw7jpzojj86yU
Mj4kvA+9YMbKRNNRIQFzurrAas0hyFwbQRF7KtONR+kQWk3Rjtt/zuIeAc00qOTH0i0ZH81g9XzQ
JiWfRJi7uPtECr1jJKWjWjqLXG1l4DrUBPus4SFoDcLed8P4H0I/ngnDqDVIIFMY/4zm0oRKDpo6
FoKjlzeaUOb9sAx3uVEEL8xAEyE0o9rp8XWYXkK254Uq9NwFobNIZq9NDyN98ww1Yr0kGSmeM/th
JaSC+btIYgVfelXHwovdIaZs0FqQmt9mGwQtDwSz6RKwJWgVgZ7dNwjUtSRf6SR0MvaLUQzD00qs
XFnc1plhb5tCzdTVV01ataOeNd3pIAeA2zNtHLDGo73kmZA/OtNuoxl1fI6cVXg1KXWPZAwbd3dk
ZtBRW3jMNZ4kjXd51PKog5pRQBDo0nmp/2OHMeamOP1V/4Z3MAV564Chj8a3csK4dkB/Tc+JBgkV
BqdqC4ikb1sxwX18WcrfAaFRzRAnTM3eqatVTp4Wab3ZTSj2G5591/rYBDdCO4usTxzfo1UZeIOC
oG6yqC10ky2gQKEHELGSvhfcKcLtOgVQ1hnQwunWN86gTNSpZ6z991XaEBQHuM2TAmLOrtg364rc
40A1Qe+YUeT4O8rHUTEQpL6qHam0RwF3XfuukZHJj9+BSQnE2+lmrXqZvl3JB5UlEQrZ/bFDBfBP
t18jeKq8dsnuxr9BAatS1e3L+Pp+iYIHVIA0m3K70jE8sNIqmsFmKRxewexzJEAiuTK8dBLIAmGi
UHyUHAddKORD2C29prYqDCGD3V42ChbIL08abZfyeoDx0oP4jYZVfdh1IY/z748HA7e6EzBQXEUr
GTHqSUC1CdVPjOV4A9DQFErOMWGCCgKBXoH7L9iZz60Ed9yAkBZerNVBBXTb+zcitvOaBbbcMC1k
K1/nu/rn32xuwcRqifxXsOaY0raKmksWZPugfqHN9dnRbSabJo+fj679v8EHoz0QneERatgzFhd8
3acJNEPSgqxtmxiHOX+ycOKkkfdtZNHW63UmBvRiLVySgHwvQdPRLrUIvXv1xM0YpBGgfekHJpn/
uFetaKEavK4Z1xT8bOHUVRQrWlQHjFv2ORf8MrlalyuMy8aYbOGQ6D1qm8mB8jQGEtOJY2ThpAvH
0huDUzWrujfKMJx7RZU7T3SP/aCYXiZH4ss/pvq2SPQEX/CQRH/yDBg5AXbHi2H21i5qjt8z8hge
T/uAmZqgwpx8DO3jPMUdPooskI2vTUto8nrucdiw7qx8dLmWOwyYOEDRRKpd77EYUbGVPhsXbaRX
3cMDw5dC7CAuIUELHTHAkKzH5lGpsMUfKFz1PYlx3iMl9Kz0aDqyFjFHgQo4u4+VSiRp0YCKsKAY
PGG7KIb3z9WSLFbBk0wIyMog19zd/sZAGd2uvCVxAUXQUqdVlfiw4ygydKOiRmr0V3UU/Ll3GUcx
rsD8L7cfToZuHz2gBUaCGwcUWXvrHbs7Fq5BnGyeORw0/mxRpJid6WjOhhTZjX2iOhoDAlOtqaKn
m6Jqrki5I2pKeaNVhHo8BcJXd8F8KOiiAjrnZ7/XlOZWSILGgfB1RjL2Bfw9NZ6JPvbb7Ab4gu4u
6oEe7pOebB3P3LZU+ZT63+H/5L8IebA7BqAN2wn14YK/ded8XtiRHLVp76fwepaW50xswWDFW9rZ
2vdA0SKNyPZGw2KmOn3rd6fDvDvkKrHGTuuk0hYwmzq6wclOvFnJHw91DsnVojqhdLW0z/Z1X+xi
vm1WC7iKtpTroUOlzLVuRLt9Jj2xncQsub6dbIbMvPDLo7BEiteCLpicDFte/3c4YePWax4TvfON
/H2c1vXlqTa4SdcircHgOeBjwf1Lhg8YygPky70cAQDEkOa1crNqweE1UNt09pOi+dRbO+fcy5jZ
hvsrvO4eIoUTR+jY+H8niagKj3cfNDiyTvs9xTCEzKVMG6TCMU+ZkuSz9bYJFoty3akVIxqQxxqp
w0Wh3dRX6blDvNvarkxdESokK8OyI9OPQ1r/KGBQjr1QcAZ6o4rfGbrynQmig39mzOD0IMhgsuaK
NbZ4Fz4VLgeQshxrh3/DWKeVmhaDPs/1QzsrASvbQLmRau2rdQPjmf7htd6s2JOP4uzYGaIWxERE
Y0KiRZf3AGlM2fQmCHPT0kHDQHbUpFNWM31GXGDluw2OEL77dwR9tJOrDT3eBk7XaWv62ZMr5mRb
mS7B4/VDZtWx8sf+F9ZfN3cioCUSRohrx6wSryGrEEfSqJLONaucYgVf9gcjZTa6oLfzhg9+qvbD
inWiGYHduMAeuXIil3LLhMtHCAaxtps5Yfgy+qWzaHUb5BYGQoGRIgEE97hC+TIGbaFYfAxuaYul
vVfKrtafeyQluh/RaxlgfeM2z9ZMZsxneAw8jc+77P/x2lPuKh4iDy5K5y8aKsoAXd0DlB8/OXlF
bJgGaG3Oqcru+aYTLqkoHP3jB1CH25D6LDX1oaYd/hXzKJqYRAefJJQhj+2aS6onmI14n8bUatDR
IM2DL5KPYrqr+qBM//iPmFyrNCnr43KO65UNNcO/XJsUgBp6k4eR+yJUTlVmdh8XL3LRhb7qz3HD
69HmuabG4LQ9iP8XqCUcXPiEBJG0o3WxEoPcGrL/0czhTCh47MTz6aBh8I8Hy1XG2ODCX9RIOqMP
S/uS+STZpcQbOBKznJBvTr3UTVwpi+ym3Ex0jtEGASv5Fx8L06RhC0ZTuiLfL4bP/u9NLHzN03rk
5T5kc3nIVRXIgHRPiD5HjV3oNIZZ7Qahur1/jYnG4LAVqgX/98tRJFtMB7YH8aV58ZXlB0xPXOFq
+X96T/Y3uLv+SXW/3mpoauMR/0sCl3MRxqJoZAB6V8AG32FUwFQKeuAxv8PBr8NZsWUOhepOZWmU
36DVb8Dua65KtBP2td93hKQGiiNpMd3V7clhDOhbMM+IOuVz41JEhYxFL7UhcOW9qML2wQ/TQBVy
XjUgP5y4zw/bra5NC11oNLRLHMaLhlz2udM9iM8o8qLgXouCryYE6N/QhcqBUCHyHIcB77IwkWdZ
6258oXd5YPUPUZUAXO3tB6mfxj3yKNHC2pYcbwv2rLrPHwKeNor20rFmffB4IelTt974GTMdfwIh
oEfG/Cp+QGIso0vt4dWJKjPhwuZmEgIatSTw8i9VEyQryapXNO3XtBo3VSE/y8zql2bnvTMYgwJR
cvpATnG86sP7tP8jylWMcEHXQeh46SKXzyVIgDubxMNwLTF+rsCqKqVqqNrrnMgDkSh3zbkbG7u6
zmrPU/y+s7DukU2aqsfn1hhvAyVaKZGdKCKx1fdN8cGm0O+crWriWN1J9iD+MEegZx9TjDxeo3DY
8w3Z6T0ynR9hlGYH1TN5TJfwimWwWmnZKBpXMhXftYV4tYcWIAdhpiyTm7NNvtLSl/z8HC5kNWtv
INdES544zeB6oFNQBysD7KZzSBa4TPZkh9mPBymOrodoHI7D9bFbkdRQN16jc8MDnT2HrZZYbKKH
tzT225yNC72P61SOs0t8n3xRgi7O1lQgjXU1Wjlx6c7xxJTFCLuvgcQi7SSNnJ2shvJ8N99/EvLV
xZdX++KYmqFXugnlswSKDXvqqHoKmGJzZWLj3zXldRrVxkkHtD6itpEuxIFXdAufkVlI6XRsxKlU
kWFaWHM4ZR5C/n4d98pHXuiLZXGnwAFhBX7c5lue/B908paF6GnUN96wshZVcXuvHrDrzbflrzt5
tXkFlB7gJ+c9tR4nkXjAQxBSpEp/zPhbfsnZ0R8h/er5IEmV3cB9Oi2DJFkDFZfM3MDVTkDxNQOB
IhY+5RP3OTaU1yMezC1/tEhav1h5YhYslZERU8OrhAHis5/EpXCyDTLdwpN/7BUu/ByihoutoOCe
pebn+ghZEHBTX66sWUWt7L3rFvBNVqY5i3Y7rNeugbSTrd2vAX+SB4FHG9uGc9i/ZR0AZW64RR3t
cRb+s7JcLfiUrII8TALNp9ly886Fa6NYgcrwbrtWua3Pb7dftjEe8qOXWa2eiMbjr12Z2rg/00bo
3BdVX6b7dazdr53PUrgKgGxzfrbxK4FBLERNugIvAwavI1AUu98wcJ50V5bADCTd2/4hCWSmE7oq
sUqVZj439mYuunoFrzMtr+h6GNaUnuhqG1TxdKanR7vMLn6RS5iXoWJcu6v6SQwTu/mHraxpoAOC
B31KRZuMhlCWMSWf74OJo1Fh8n8hJ5TSDRqKP6eB0pyqFYWbQpySLqeWli7wkvzkhg81qTkVbjp6
jUqAKSL0ntBYzZPcdUC0E+iKzsTTR4DxDFqUd3LgwqOxzRz0kEIAX2DarS/4Kbsv9SzD3sCucTgi
uAqAQiCM/hGgwPxw2J5JQxnvseHjxd57XwFV6U96rgZLPhEKkWpDpuD4mIEH1MAdAwpiZK6Moovj
xLl33cPLpcGWbUJGCJCii4XyvD9ub0HcBdKk8q6KN9nA2OCVlKiZxOdqRdB1YxwZ6K6h6cO4xHWB
+p1QNrwmxjeEMgbkJy4zYHnifJAmL6OaQzKO0cbnGYKQRCr3zAImr2Wdet/sYGCBFf1GbX7AjIVQ
mEOSENT5XYPFw6pFvaOSO2ovnusAVhoa30dUR6OuVg+q7j2tGNvGozgRBMnTIkOUD6BF06FiHGlF
eIV7P8N+hJoflnJqOy5WwzouWLSapTTArX5P2Be8mw9sAi/J2dWbkyyV95OrPJioFGJ1oQqu5jQh
Ri1f1AGqijm8v0roiWgyessiWAh9hBA/uiL16ocIh55aksRfXB7svZ4N3y69XyFIPxl9g/2ZxNuw
YzblmO57Gk8usOuLP4Up6oVqH7ocibXorJm1GkS3YyeVH9ehHzeY5cgXgzd0dZzg2xThQDLyWxYL
Q1a29z42BgNkDDbhhKtVWmATx1zYBo9/9FDtjibvdux3E9L/A2zuZZvBWnc5ggJSwwFXDhGUzwYk
fMOjd+i9YKICglm4r4KrYNS1ZD0bjsUsXp6z90MCLUpPTKGcUFWFscySvVcPr1nSesYz5GCdVJ/X
Onl5zGPHX7cvH8W5w4+nQyZHN1gz8u+jCUELy5GZEwY2+s2EjTihvSNq/PjzgMSocEub0uzIOlRm
X2GC9EwdFG4Z7/M+RFrvGnKJtK1LNrT2NYFN4SsuU5wvyiO9njV7OyyuLsaH6djhoXqB7Q18ImT+
P8fani3ptKK22NgHuFHh1YnUbb5FEYvHICmpeC6uaH4lvDZjDrvYZUzrtgEBDB0+TjrSk0dEf0sa
GH0OULhwWXCh16QOWkJ93tN8DHW/zNS6ej6z4Mkrh4BVsnJg9y+W3RWyvO1zk+8WC2aJvTmvUl0K
CB5YOZShRiVxXrz5VvaCL6vcLPXMptuNUbfzbHVosbw1Sn31JQyPr1SvapQoklIROaYDZvm4zTl1
iv1UohfwmlwmMLACDt3J0kCboDjrkOkTIN8zVejitgMhTCVaxtugKj9IvC4BhvmszDBVWFnM+293
jYPZs3yMw5zItfjPh18TaIPZXnNpKXbBgUu95t6t+tJz7ZXgTXixH5efKuUvO1jSxBaTHsgQxFPs
BnYtJG8figJnOpQiymvKZjyvjoAZsDLELFu0Xcw+cxZQSrP8Pgf3WVt/29mVFfxh4B/8Yi3sK5+K
xL/OEMAP5a5X/S37zRXqgQJFh/a31/59qrggSMkfifjC2Wz+a4981hlsxo5A6UdXNEJ4Au8BMyur
7paeVr5E/dRo0JP5FZmnCARp+Xwjt+ThStjTr82bg4pM6PR4AOi0CsYZdbxrI1NPaUDw40qb4SUF
oOY8pf+eBpDx2wZgOHhwUxKNiPAOTzy2zmygIRIv3iMkUDHpdbkw00YhlgiCgTVG9DZsiK164DQi
dCvGkgU1jNyV/O4spnzDmgMoAymIQ0aD6ATk2/UdUNKEcVM1hm6xGE4EiW5Kc3C6frKamXXgL+EK
NqHg0ZkCQpo847sz5xoLp1CYqpSyDalWhu/3B8rfLo4ftosAnbH14AY9Z8MZwJiy1wfmXKYvviFJ
kn4TdDEntliSjWH8hLi7IXAarBv7c8mAhGmbtlMQL5EcRBwzJ4sdimSZUuYmicpR5HREJRubPY2z
6OKZfDce29hbsv/GoMMKetnGA3yjaDLZNunseE6daM7C6TPw4biJqsOCRjFq6kSrVa8Gc9rKEzw2
t6kjuSQ+mWTQGmCs+OEvFw3ti578dCzHNDhaU1Pco42QfUWNNXZOJxsFgTKLpQpYMCEaEknX2f0h
iWSTy3SgrlNHmI0il/JL16bSDtZlLrkOUPSk6pbjXN5SG0PG/daqme7rFpV/8BCGrAl5OmhdDF0S
RsVt0zZwxdbVmGm7KhlZzRMf0fA3YLLb21P2KZJpBGxduqWQw7BfwGdjc8tH5p5CxVhW/Z6cQ471
jHIKyinLOkE86GY2NMy/pscoNly/SfLPEaVF1+xbzTTCEuGuTf4Y3z4ORekF+nspNn1Kvk0XnR4V
3OG25MCo8ELLLBMkvtbZ+uJZhytTIHvLF23f4DpjjGSN2HodQR46pYJJbvd0jXtXEm7lypJFS6cH
h/W9x54abOfp3AmuMpgAwUQamhjAM56AuLWfeU1XYsNsib3G3FutjWwrkl8qAEsl+eoXIq6Lf4yM
DKH26KanlFr1gjeAQws7Acm8CdAsS2gvB10RZzhMrhdDLWeyaq7KHtLA7P4FE9pMaYuqqBXbGGfB
5n1/27yzf+fP1zryA366F/Mv9a7YgBaq+PKZ9qhbsLRVVzXQAgdboevzPmsTsceo1otu5FBvBeb4
YR0naFstvdYs25+03qEddOeEY53efUWxPglycXG31ncMtVbmeYykwv46Yuf4w1mtgv+57A+KeVp9
r+4+7/IJY/+XH7LX/PDsqiU3gwIdrAxvAnzYyuJc3R/lAWBEcszIyQA7++NfrmDeKJySQBxx+33T
cLcdXbTtuMNGsVdI7Y7pgd/FyzhWS9buAdCP1sgb5oMOBSiyRvUv6cdVOEpFQyV6I4IZbHkN5pUS
wDKCIX1RUzYy7eSZpmoiHVVDdHJSpQp7rTflnEulA5NYxbLbJdXobV0i4HP0r8xRtscjFtBemDc1
fVNiazPsauExLRFWz+ezN1GtoV4eBojMGVcXDRNo7UuSeo7jWfOKtlRsZVZxAZPh2MRjlDzKRM/f
w85H1pd1cVtFn+iHGM4U9r2oegz8qotr+1HMbqcGdYCYdi272RyQOsZ48/V+OssLpE5qi/tqrUrw
j2BTmttL09AuX5ImwArKkEClmcH9dUnaF+JCYvyrWaGoYXmCQR2tltWahYBjRKQeAWpf/xbc0ndB
L/2vITiMnq0Tsv2k41/3Vr7us0YtumyWlW+CjjyfFkbZOpKpWk8ijdVWqhwRldl+1DTm+JicP2HQ
OZQHgRSVDGIy/q9hHTE2K+OBUq39hVQ+W0dDR3qHpC08qd8d9DnFOJl9ihuKFjY2sNKOo4LFdxr6
w8UYmu5elRLQx/31F6ZGSygKXf564bZiKs4vB+LAM+rQ75E37Xb4LYsfK1quyOP6z9PTKlVtp+Q8
A4zmckJS8jiqRwvGS3nNWsP6HFQqQ4VZjw+sZj3gI+vlN/FChSq8cf3AI5+gVktLxlo1Md68BeHx
VaVr8kp5bre005j9bMykcBXFY4ZY2cof/wfY0RKHsyhHl7P+AjxdByt4amlWnIuZfKii4CoGADNa
NC0Pk0dgTOJY6eJTrxvmEkYHU2/gF+pvzi9WfN4eG9bMWQwlXlYK8kMIJwtvwbTxmaL09YuTCbio
fZ4BxDHZFDVCQbSCiC88WKWEkMhIEjPOAl2Hdewusn5dJijGClKADb0Ro2kHUTrLwczz1nBiK53F
QEJi4pfC8dlFDUgnTUeDRxWiimKPg2ATQOZ5Wu27NbTcbLoKs0b8Cxm2M3irVHQxTmvsQoyit28m
wAl9bmchhotlvP/IUoznYEOx9Jt1lofvPXgZqQ77wtH+WpPCEKq01Am3hTUUxi2JVh6gBaHR5t5V
yjoHMr/8iAiGqBlncME/gi9PRz4CZrcvUBkJJ+K8MtjL6Mig0a+8x5WAeM2HAjHinthkuDQqctHc
dHWkKwcpAxT6SMT0q8r4m+5WB05ML3ffzrzPXEAv4x+d5CDsWDzp1VAZz4VaFsExCToOE/GjftUc
Om9r8WwRaMENvzmIjKU9dZ6U0n3auPpLExSjPDsPqHAnJ5H1b4McOIXc9PYATrC49tDKo74hTD9t
6hnBh7pNaKItPM17Wo8Y6QzOnAtJvlOSSA9gr6PF2SUlKgW+BNzFWNYFTliUw9e3Y+93YGxYLDMo
y3AzspZ2auPDsqAbxWtzFXFZsivk8l6A+ZdfPm2SDJux2C3d1OGahBE1/hwFppv60aNtCT0PaQPy
MgGoyBUR00ULdY26GAp/e15GhA8FKMT77wHsARNSqCyGYGaRMYoK9CNrJUAxkAnwGMhLt7eh3UhQ
Y6f/tpuFsSpDvHMC+S6MS1DOH+j0S9RcaM1O9LIY3IszgUkPSehZ9dibs/VKo+cx7l2HRos0UVSO
V2FrGlAUl6yQ6ampX3TnU5TsiwGAEK9SQGTwpZ/B9MKX4QQnHMq4/8hJLKgA7yOBsq9TuNBNiQIQ
AjbvZ/t4bAkKWTImPwkBtRC9bEQi4mE6scw4pLMQgXOBk7gL8Q5LTwyaiWf56wI9PDFYBSWpS8bM
gixMgZd05Uz2nWF6FqX01hGyMcThrrpU/bH72WSR1cR3VepHbAtYn747WmKVvIJZq9ulCGHbIKSt
FE4pfaf6J2x2OJHeP39QYgOs5pvFrJZf5mF90ZxP1uxhjvO5TQYV74WeO/zY+GFbfVy5D7yG8ryX
5TjYR3CNh9ePkhR4E0juGE0zE/VX8lA2u3Zr6kduCmQrFB8ykBcSpL6Qyc384tm65SzX+gLfhuo4
zITYNpGddIcEDavCFK+cfGBkU5X3ldgGgDLkdvIQj9iy/6U8xZO3TZH0hT/3DK0XRVRNclsk18eD
UmrSIU5M5478DsPd4wn7w8PDVu3Vj5v4mHPtBSWqaaVpuyhsIyweMKMFUHG4yB3rz+k3y3yzGPvk
xPrGhP5ibtRntl0S/IlE4qfSsPQ7h7TUOWU6xD40InQxak3GfUKiMbmjaZeAsvhmMwbSyBdXh/Ga
fF7ewj2973JJshtZkI/Y3pdWe/VodSRKXLVY70ko5MduLEfoSwMX/2fwVk+dqw/X/SwZtCzuvg/9
7RHc55LvH9jsg7ej3O0tMdqPfdJ3EhYHYgJQKT2T+Wl3qeVc/RtzL6q2qo102PYoDEUO9qnFdVHJ
MIFu3i7RMLxHHCrdhjkixSqbnwK6Wn4AhVaicDI8bpmRVQ2stgXgf1OoGxEzy/KtIslr/NiAdBdg
JXJfk357HlWAYokn91NoOuk+LxYdGSUwNRjuES5xhUphpc9Z/9CBFIAehnj0tvYUmpNZPbo8p1bn
qU6QPQntua4yuEHuQ5APXYKKl2b3epqnipODf6yZjO8c0Do+cJEjWdlH3+whV5Xmg23IUh3hYI3y
m/82C+Wli5RGTgo6DaBrA+Z38p1DqWCxTKwFSpLcWOvkhjzUR/hFLo8W6OLW6qAKw/oZ9Qgf5IC+
qzN763OOtG56QC7NSnQysADsmzhkEeSJ7AvBPsvrJrZU0Jc24wHzT3jJTfc+4M3Dz74Ybirjs5y/
rIBzIVWw8w1jVMzEKW9FGOHCKMv1a7GwJSMrXGAjf3VK3FtBbjHlbixsgDcaOH4CBwqkvL8V1zLk
leA1CZZbiHc8DGAR8BP2H89lIgbKLc7557ZSy0xjRgFMq8jji3fK8EFQg7ZAjMeX2fdQZJ6IW+PH
+3bBGzw0NVkgHmzrhcYMODS6KXlXE0LjgncXR9aTltI2qm8sqFhPsFssfb/FxkTZltmTwoKpoGX2
Zp7T8vxcRqT6cKpRcYPNKB1xOqfRp01Q9uRv1+KX8dY5mw8qdtMO1j/I4ChVNRt68yFNbAGY6bNl
zg7w5yUJLQjXfEPT7eUDDQvoXU54LpFO6Mg2mNnazwXnlevmilcN9fk5EBCRBFOXRWNeS0ruNtda
LBvQHVI+xYAdhUIUsSfStu+TVe940+pdKV4pxN1WrTf8488RQXxtmx3xziTcvW5avquhkmTdWiLg
v1+KQH9ltfq6B4Y/1pmZtI/gYEdy62/uShGJt8lmQ9UwQvKyEirxd25DrSG3hBDVDT2yjUXHCddY
mq8zXK+s0zky/nsAyQ9u+4uJzpIPYjswIw4WHe/DGajAu9/yI70Ahix6FTDNOqBONuRe9CDtwPVA
ygpIH3zwriuTmEP8eQCqQZbs8oNrGqpf6eML3JGMh8TMmTwxBKP8sh8UrH4dXRWXFGliHzk6mveD
/l8QXunmvloL0PbM/UjqNe8UJCDT3j9XdSDwHr7Z/T6PAAkNTAUH0wodbZ6/Ft8lEaB7Oge7Rk3R
y5/xnTIrJNTK7lZie8KpraUeK1jky6aQxs8fcx7UP87c2AE/Z3x0Y704DJ0xyJoL5nuSHU1DzVdG
9L+tiCHeqKflrzEIi2664EQ4k63sC1WSVr78gffeATMncsdzQPralXSbgbtKFyMU46zOQnMKXYpf
nkya+Qq3l8XZj7V+SFdioU+JbBeytqR4jvkCcqowb/pzbM+PWbNCRtUz03GuUwJ/JZe1EDjun57O
UAG9NHPgG0aTwNLB+tXAHyU1//8ACQoQ/rNpTEbD3yIKryhkFLWtjYzmlXTM0BUxOarmgv6TPsUs
SCV20EUNfqFACIO+GMJ/MMg1FkEa0sGSD82XEhi7igu4uG2A0r1IqnZNm/653PLZS4zdfyGHLdMG
Ux45krh8DXqNM5cL9fkIDK09+xZ0kPkTik3Yy5lSalED+FRB/83xSv7IdQPUObL7Ivzh8nTkHZ52
RtCUkdDTnWKfYwnWR1O332/5GIykjRdngFkF9bN9XfUxwlTlvK4I21HUBCujOIMDfiX0Yza+0DaS
U8/qBfRSitgPQaVRk9Ej4/rlui0LSa+g9HIObXzHhEY/BQqmm4kP5SLcP9zKwCJf6aKe/s6MVVes
y7whEwbmdX+q83xACqIEG7HoWJmn/whaf5GHZFq9RikY7WMsQCHYYis2f+ZweeUTsc2eAwmRDuRC
clahqJ+RH90CNZ2a9ZJNFu685Kz1+RceCegdvVthSfwseSsxKMW4986l5DWS6TDlM7KuSblU21E3
ofjbV21h5VlAhVz5esMjNxQoEIfrJH1Iun60hKW1kCejad4RNaytfPCfNOxh2X2JndBI1yzPBP0c
zWYoFZ3ub7EMwS2taLGhhEI9KiFT2o/SLiLSzT0zfksEsPBaw6bk0gI4FnB8QcteTErvkpSgnwOi
UutIbKNbdAU1kuVjojD5ukeZdOa40ZtYeIhKs4CHDJzlnfw3idu43u6Yb47TFjkbacjTj7TeNbPi
SOxvY1tlznZK/2Sd2PaQGGuEfGN0BKUW/Zho2hNO6kCaUfKSMz2u0Deq804ufWHdUEq9dB4xWR50
YS/wmHyK9p4CxtUyKk/g+qYqTLEbcXbQlXvjYkZCyg6LrlZ4hPNEG6lYURQI/B1Oxb4fWpgGFGm3
puM8Sn6I3owt9k5wF2ohs/WLTqB9etPQWzedJfk/UNALl7z1AxgldTYI7Oam2uEFm2tvXLjbzBjy
4lyRh5xW/zwzOAAC665kqbRok+7PQbxMoyeT8Irg/bfV8sO4IS5rAsbOSuB1uunlrn+/aXoxVKNB
SE/nBE3b9CbbHa5gPvFBbvQD4iiaqsTl0dYW7Tr/k+9QiWMzntBaJNFZq8bgKukJe+87rwlzQhgI
IU5I1U2+YV3B3srNV7bObR+cF4Clmr8bifzddRQdHquAOvwNuhkrV2BsfFYTRyPvYzoNL0sBkyzx
MCrLfQR5I9wBbGTRcaJK10cow+hGgGWItGZoRiZx6a8z13RtMW1kbGm0KlQaFprjurLXVUcAro8A
w8CukaWTxq+lYOHQtrOcojV8qtDCNbEtAonJV6vjSx32R14NibLXANki1RD+vSRkH3kaBGtzDAKq
anumU73d4SpoXjyYvr0f6yglieeEnux9xkPrBK+Yf0uh4MGHggA6oxWWKM7tDbKaYDr8R4IVZiWH
lQ2/U3s5ZeOQejTWH6MdA39jTWyibKkCEMwDy9RdDLNPlYheeA6bUOHnpuU+i/As+MhSJPfO5/gD
c9NVxeqg0JG9yw9AS368wwbjm/8OLePFu2u+0j5mNjUriCT49HGVZQH7ChYzKXDFCzpE4e/+Agyq
1k/SVK9uTeBGthLKrdHI4SKUFxSHUkS68i3anZbSsdbXtaQLvhgSeAnxPMbw0Kb3abGcT0/+0jgJ
FSeD4LsOZfzOg0eOu0h92MVmaayUy1uO+4uuz0novvXKs71NrWkUTFSZTMO361imWv5Nq3T60NmZ
fnH5u56xMXwaujMztEUrALX059PZd7qWMxfV7LWvmFV6tcqvuPDDybjRpHNH0Xgmg1HokMDCd2zM
po6mqmA7/PQL3me4nrdKo/JFdAHEiamPsTQnXd3pShdR0fuBFuP+7WV01BOGwarIrvRMOGTtLEhA
MmHQ+cupswGCE6cuQktWkOL5zO7npADjTW9q3qPFiSxjnFoRmZDkP/krAYv9QhKDmxtsKA35O2U4
Jo1FuBU2PaXW+OMjPrBJu0M7OIo8KBh6n3WVg+uUDPLBPFGEo7CjV/hFJXsFLgP/BbG5AKl+K+67
xXUf6hcKyoliUNz3WlUNrwfAZrC9yEjTKURP+xwTm4AIKYd7X4ChKG6p5mA3/WufVJhwjEsTghE3
vdMcUKBrQxfFx/mlPOMbAcXLHeWWZIC4YSG2Qz92JxeSPaqQj5dIeyl+LYtWu2xFQ5RfmEmB2mvQ
BkjG9g2e3UFKok3e9CWG6Ed/kvW6SaPpZDt1Vs3FCYXZEveu7mTtZhOTVjw9mfY0mgWwcRaUMDr6
Yo1d973GcvPDS+XLfQyDqYaZSdMotRRZIMiozqoIP/k1tJMxxVrwQYyNQkwttEUyd38L4NX490C+
QeRZ2ltt9tcfz8XZnyRmqMejWcVP9SaxSv3xBg3lnamsc6eSkLFxlnsHeCPg10FlcixzvxQuRAne
RtifollvrBc95ggzn6TjYjTry0VAlX10l6OWcbR/rvESdzCmfIJSrlYCzJLQgbYLxM4gebp1IZP0
lDFRL9syX5h4SClNooegbAYOyqb+98gl0eqq0fadi/zizGVXUgGnXz+EbuVzKepV9smMDaQ1U24u
bAp05UUG0mL4HD68hvfJxOnBztfZkgn7yTyMm7yF2xTtOd3Fv+2l++WMolI7Ftj4eNdiTg7geHHp
6Ji4HR5IDoEn1s8jcEo0mTrfuD7YY8MLM+TTMtn+lbkpkUvDNFsnRrG1YvpN0vMngUP3l06wRtT3
fj6CyNKHUqtLFD+GsEWttLo2wUgBLHFCJD6RdJhi8f35Plg0sD1tg+W0mFqBt7fozRAlJwjfKvgo
8HkISsnpLjQRyEBhevAWQSIGGKbqimAVZmo08g5TAykwbylZRlxf9w6JMLXlw6038EmnwpFPT2u4
IUbbcEW5wIobqe8MNypCrJRSe5JcE9Jhcj//eKAIXzkZMogpWXbebuGuZ21cWO/OsJ08/Q647ePp
FcUWhx1kkUG4v8WKmZWjwraHAPXdTBcnqtt5AU0UtEcQfFoiO/v5rWFbpn0DfOOWfQe7pvycCgn4
pV3WdfS8pjAoqEjIJE7psc0Kmp2wrtzD/T8YcHUkX545htYrWkwNABbT8b5xetoaqe2F29Ne6OI2
mxG1gDqEJQnnsYLUqJIYq9ZCEzPc09ygTAr1rhS1He1UKN9apHo4gmERHaqa+x4pSWxwiGJxp3nj
emg9YGSMEKvgatnqJlR3CVLebJF58k7z2PphJ4OGdvG0qTWJvkuJHNgOoXqf7zsQlxbYfrvZuO3S
s5NI1UfnpOE4VoaQPf/gt10jFSMQDL72HcT+lR6v1MasEX9rgbVcn/h7THHMiW95ephbMOesqVAV
8qQnF58LQG4LIs0HYBnZoVlSUt+R62zKZPkQ+Tw8seWUv7JW10tJmz+znK22ShIqEnqUkxSNpvxD
521oOTpGg11QmN5iJ34ffao/Ki7ZzkHDi4N6hukJAggwS+POAQRstsRoHJZfMjriBvlOC/XpU54H
xu5arHObRFe0KG+Aa0QR+dAciUNI20k9KrILuG1t8cv3N6XjsNKo3M0zUMxXzU9QtN2dHSflemKK
NfognW2r39tlVdv7h2JqfbR47amOc25Hh1ZQdZbICe43atEeudcD2/hhnNOCgn+StFTk6P5o/2t5
PBPN3ievytA7rAjYoieBDiIfzR4q0l0KEnBRqhfjjWxzl+1t/wQMp+hWNK25gNdLRf8DE1GN6rQk
9I9P3uUYN22HfjFxAzqUzyZnmtczGzKxKpx/NSzVzqNDgbMjgX3NT0eD9c3QhuF3hIH/VCaMYdfy
EIJzEJ8ZMy4lswu99d2xJRzCeKY5y+4yBhyGaF7d7Xq+nXTt4U1MY7j9PqTAzWFqzmOTCE27TNE/
umHtZyiYwOialKO/HNs6ZyLcjJwFx+XN5dLKpwm+szxt8jlR1FzHFQ9Unqv4Imqj7O2bzCoxzG0z
uqwKFMsfJPY5GeyLmGouAYUca9pWRKthPJZf9CJPVTwNRau+ucRePN7mmyS3CEN+jDLGrnS5fYMh
+hi/FXPR5wr+vddYACEl1p6IiU3CHg0N7Yewi9M27AeQW+5DEVeN5nT/xCIslRxASI9XVQS1vLAG
HqYaGZBJsukFode7vvH4L2hoYRrO8hUGXzfvGrx1ZQvd8H37xuwD/sgpgmHufhJBKMUQeDjmPF4v
4ED4932HnKtid0d2s4oT3e/BAi39o1nI1nPE+DHAKtqpPXSqsgmDL+1o3a7W43i0wNoM5BpQd4+n
pJd+N5m/hKtXP6zYYlMrrrloFpMgtk6mzgjNIGJPoV91kI3qnBASu4JlV96m9QMWydXZ8AxOWY1J
EeegUhETOKHVh5HKFcZZRjWliSTPXeWDmRSWtInajAt5Fossr8resjh1Yew4nFqFsL1gkozns4YD
Dn/VKDNDCTry/adrA/rGdG2CUcapyr9SMv5lO1hcrDydePrb3tk6Iu3W9lzaCarrOvo8aLxod9HJ
GKsxX2PWE4nuh7at2XqbULcx/TJSou+J2qmSFFJAZogYyp9JRtzb4FICNrFqOBpjnpcpnRvLciky
5bliQfNmdJjLIVTZA2VdL9RFliYwdKTENQRRboZOepDzBpl7KccSG1EETFvfrHkSdCFVDw1ObNYv
bIzEgAWc2r1yDVer3hfYuBtAwncNn6qNK0xdSw0yxj8FfY3D2tKkfLrSfP27o7Eo2ZG8ML3jQlOU
R3ffZ5twyP+QL6pt4n/Q3RJSyr9qqP5v2StJ2ZrIds3G+jpiSavQnuyCP1vI7LN5TO9KppV/Tr4b
035YmgjutS9mEP0J05dtng/+6sQrsgnHuZ8Kl5jDwQy4j7wk5/uQZBz6hRIbBuU4wBe5tUsYzPdH
F9YKTLiosIwyF2WjOOSLS7mXlDZCMo75kLUj2n6GD1mKeGmSCYuKTLYgst098A+ckBmZhWJ1RL5N
sfG0WaV5KPkeAnjUVQB1Mz5omlzZvmid7Epm3AzyCJvl8DezAMHMc8k7UVmqKN1EqJ5oWwgp4QOn
gJR8q12Nxcl15zefP78/7EwO39siROxITTKrs6dXjfXSHSo7Z6F0cHxhu/Tt913asM4jrw7mcY2V
3mNavTtj5hYpyIDfW+LPVjz6ezgCBiS6ihHbO3mogCLa2HxfTKGcyW6s7VxtuDKN9L0cVSohif37
MaJNdG56dL2DzUcVR6tKOtHxvQD3ssisADZcn3YLTXfFU7d/rRaKZWOQ7LIwftZs7ymWnxrwZqtL
eHLTdzmLGeX1OHFRrP3KRhCcgyv8tTVikYprKlkiBUkdu35tzT+LuuQkegS7UXrkGj7DmAPI0GA1
EHSZP4fRf3HqsFxa98+EUjYKIUjb+kZ1OaqvlX8s0XZj5/AJViCFWIgfCEPtRNYPWI9if6QnVaeR
LuXeMZND9W2N/NALXHvT15dQS2xsKUcZKMK3bTR8ffZPcVJE/Tqex71x0t63u+sH3Y6K1WWIWmy6
AHi3SSBlTh92D2+Bhvv4kn2kmkkfmAADOyJOjFqtFDlg1SzgYyIHtWDSTC8ikpExgrurF8fadbji
6c1Khe36NzLp7MPs4eiqg+4/f6PMM24KUrKqcZIQiEbM9WaQREP977K6zcoEeQNu46IISD+C3wii
kuv3DtJWYxBmvaOWZVlt/YtcJv2adBvk8cl+OXMsPAAjR+PkJwmEsuvO6GYdZDHJoUF4GG4JoyFO
3ZXDf/gQ4uJ4bNML9p/4o7RilOtjfeV8cxkBqGtyT5hCslyDJqwNnuo/smwSnudBr0LuEMU4N3Ss
XyDdeGnk6mxW+NnsN1AWcpAPwQV9x21lY85M9yTnbfROTHP0prM/nIZHrYHWi8a3Fi6EgrFj3Dk1
S65xkGmypCZj42zeslVxXsYFcDQQ9f+Hz5/6FtSc5P9X4U2jk7Sq6ZQJEcAQ0MnI+PYwV3yIdfLb
v24hIPNIVXc259AG3GeTdbAhR/kiKUKpMij46Zf6mVUAI4aPXQC4aYWSdwzTr8qt7aIyinpBXFhy
t+WzsC0jyZ8OYvzPhsKHY89deNSVaoMPtElzpTmTmUi+SUwmVVnP3K0u55pGQc7CWXmVNrpkmAT2
g+0MGmveydpYxbZWk2dZPVeGaQY3ka8e1dO8mrITFSABfn6Lcrsu5a2Tn8zd9xqHnHybgHOgA4X9
fNI38LVzweNp3v+lQuTWChgscNc5O/qNohhVYjfUo9vxwti4fIWpCUZmn/XXYhIlsOc0EInlCdy4
qN26fOpg3J6igl9rdVs5lvVoywGAxVfDSs38XzOhuh6DdDMceW4tEx04bUHRVocWdVK1f1uOmqrh
X3X6yqe5UKfqIxhv0+Zu1Ve6Nu+0/W2iTx60+Qlj2wg+hZMmDeU5/McDK1KpIhHe64JEccBQR4S0
KvCmhjU1Px9aMAUlFNjIIUQ4Og5RqjIufFlfdWgpAVjsweckpTtc0NhjUNhyd4y7Dh6t3EUGgBYs
2D2sFlu3/rBX8SIdxPpnUmJmVhJ7ZvSa0hSsV07cnFjMTrf8/Ja6yLUKX+mZRxbYTrGjW5UuRe6r
ozIgPpoSsPvQl42OuS+oaShKo9b5CY739BgI0f2bKHd0mrByj0XzOuEQSTJk15S2IAthTHCNjQ8M
/IFeTQv82oL6aFAmknsypRiibGjwPdib6vN3xXDx4dLi+cw+b0o5hSERcw/n5zTZXstLILahWgat
J9wx3OhoRLdLOgWlJaNSNTOoSZzRvGyytAmlYim+HAqORaN2JkrcygOyXAGlR9TUzJzCsqeCvszQ
pTmfurL3E5SFJsWmG0v0YY9nYksgxQWoOUvNW4oB3wGPSp7CchXNsIUpzpqss5gFPIRsYoHIGdrc
a+mg0n0J0bbRvgh1otdhwrZr8adqmYg+PAbvCsydegB0Wz5gPJh+FIwfk+XdnJUX59dMKn2Fmevy
Xo+YSHoy62OBkMcoT2LiQTDCTFxHldk6H39E3ju7BW7thUfuY2tZcz9UTaR4ZvuZllJjkmwIs6Rn
+kYc60Rqi/qXoJCAu90iITMWiFevhNk3Il19yie3Wj6BBkE+SJh7GkzoRQjsBisney/4Jc/sn+cN
f1O1KEjFqjV4X72GBcNucPxx9b0ivEYCQo46YjMm8P2GjTQBhIHaatWKjrf16GKwCMAicSrqnNEW
F1ASJGLylA086ifk8mkL90EMQbahen5PMmP1QJG4KC90uuQQw4vHW/t31nNxvd4ZMIIsboCKSuDY
5VOz2QLP0Phocr+gkJHOv6hoNyxx7FGyhAdoDksNVKbIAklC7CXRS/ls4OiYgKRxXc5K8yMkS7ZW
UQOeM/CT6TKxSRRnnEYUUwUjk8yxdfS164+GMY59Wr+DVZ4paqeyaDW7p7EWNyGIvrrifuOIIlWa
AdyTOVHsrW2XX12ibLr7fGa6Wf2JfoF8y6Ay0TAO/OGDwygwjWyBUs2oeJ+WPyxr3xGBBae7aoXp
mBEIjK66Ej1+/LkuQ5FAsLWxsF+AUbjhpdbecMieJchja23JoVpGP5nNt5PCzvEBmBuSTuAze8vr
kdHgxjHfYAwhsG5ZWA7RgzIEuijNy6gohCZdpO3axHYdZpRiOVgJYXXwwxnHc7F2Cfmec7PoM5xB
FXydByIP1lH+afQOaKdIkcj56VhZwahzndSK0p0XEZs7o6Y7Eb9Up4Or6KMo+HLrya0fkhyDC1hf
E/X0yDeb4qNe4ZGXZmssb0iTF2M8p0+gIcrRfj7FbeVe71JugmtrX7q/NvBJ01zhtTibZOjpGuej
t3soHv60/rhDAAYPSJRX/KBcrpaKq0tlatZ+AiH4nej0JvfGFw+mwJpE3xQn9Xy3fNLgMipAVvON
YKDAkQRmO5+qfhl2QYIOs51YMTMgl3foN2vfJP1feZHhI1BmJpfCiEqy/qwYTc+OTUn7GCw8Nr2H
3lK3PhIT+arVCKQDwqm0O0O3+MSBe/a4udUSeGeL0LAVtkhoQCHeLddWIisSXVUzQuz/TZnAXcIY
g+NnSM4t5w0QEdZ3JPoXvnG6DO529TDduGYq3TL4OERd6FCMtrGMjy9wrMMcggCIBu8z5ZA4TmX9
av7uer9TgQUrq2ZI8pmYYnPvBJenuXnSQ8yTsVf1K2P+kDv02raAA9zYBYcA1Rab96Pn0Cumerp8
qdSIze/TMxg4R6TZP7TILdJF4NyiHbBeeSva68z6fQgnNkmNTCLWf6SFx/WrHvsGcN/pPf+b+Gcm
mbAi1hfPN6TavxfhBd675u9Nv6q4r02pA/icXww5EO3050W2F9BFmYcSbtKcgj3yWPolJRerMQp4
889D13aUwPRNPgvjvLSTS1NE/HmU6lMCEVh4LGU7tjLC6/ACQg8ufxwVd6zLCDEZDgSo6jzWfoQI
umybsXmwlgpRmjezRqVsEaQmk8HX0eyIpqZBnaIcga2GuXq40dcmOPLWDWIss7ImMwi9pMYWWFCN
ShiL4XHQCuPWfGGAwr8tuNAVHnnxWmi14OoOpRQ6LCN6fkl8VjjDu9TOuLqfdMPNLk7p285zokD/
zrMKxjL8Cy4T0BIBlB15QBNU7w43K7X0IMRreA7BDvxEqNkc3iFH7JCyJDDdzzMZ0IAnvps8f1hM
1ntR5WAUVUM2SzYlPK230cKIAVk0puR7nn18QVHPlkzKzHy89gETIzc6Tcbvd1rcjugh19+w8Q4w
K8m/Eu5sh4ooXFE5kEEpBGiWLbDNTW7nensfQYuPl5sRski9grGzbPoFczGUExs8NlddDhzbM9y0
VIo77zyZr1l38We9XA7iy+F6PQhnvwdIpfv6dLa45X94OLndbeR5mHpNl/7QZK9GIvZlqnuQHmCw
HoU511p0WP9aqVzwsJQK/5okmb0npVUhIrQ8xo2ulm5+/Zh0ualV1nNmkg/CWLyzIwbvWfiPAWo+
/iujv530W/aTg7WYck28EjaPHnljmZrWKvK45Tb6TiBjyFBvrAr/UzzmwJisHq30cqdoYap1KvjZ
bKCI/zXJYaozwVmDRpzItxorZGIxOpmHvMsza64sn6DSWkXYqsCh93YnvuZDWAIIiKWdxY7kia8A
uc8PG8/enXpFqLdQUkeZPjWIZdBeaIWK+yRKSZ4A56skid7EO8pIHgd3T3nwXeL7/qhB1jx2Zarx
2hE2xtnEKK9QJah+sqrD9QmwNCLm2pmP6qeWj2TVrHR75hTnqRglGN0XQzGpVLxuWl32TRE9dfEv
QrLQTYD8saJ9ziof29eNj9QWrenprAMdxj55+EP/XUaMleLxw0jhlO6RK51SYJop2q3+IMlF0fop
HuA/DcVRjv+Uc7jn9CEny7GJvVLaBJVmyd6D1XjPhMkbDVMxXe1f2p8hy+afx4fdDPCHFqr6JF7y
cy/6oZbTxLrx9dUzdyH/sc+e8cmxWmaSM4FjP+AlP0eg19x8ASPvdSm2yDmSdNPDdIlIVHtf5cln
0xsR5le8u5oS7yjCReQXK6AyF+c+sVEWL3AlscxEr9PlihDvKvu2PNerLtG0fBo2onpQpjytdTcZ
B970EcrDjZNXf/7uqfuoDrQ5qQHCAQ6XrrVkLIngzTZU6R2KgZzRR8h7NpEKE+CP7TEFMQ7V7cV2
iASMmwEVW6ekjsNqN/FS5lEqEgkbP0UzbxJcdbOj/2gnwfNsryBxS2wRDwyyIIXDoWJW4YjFGzq/
GkeUKKmlT/sDLn3mHt0demNvsQj066BWAXClJuihpkgJgNuMinCZPqeRaNVaYlrFyLw6IZ6UUihz
DwMxbecd1T/ArlIuEOso06QbqXSDIM7beNImq0UWP0Cyj0YTHrWI6cbB/QfaLwN9YengArV89urB
DUQTeDpWWMoCP7rHaSRrqyFLnlVGvv20wT+868j1ff5kp/5gPn3hLeOAhCxJDecO1ojjfBq1UP4m
bo3BJVNnxLMS+/NXqOZG5s9E2OAg7eKwFty3Qqtifo31Im1TuWPVkrWMIjQ8Hum/Rf6r9iaox6tG
YoAJVi+lmO5G35sk7TPEdUZSiMCGync4YG4ZsEcsgXNwZQR/ih7GRKYv568vfDqm/mHyqm9sdOLP
QIJZaNGRueOA+5rXP6Fvth1s1zodi/aq893JlyZjCFv4ClI/6w1XzTOEHKBySZhECOX7SXBCqTOY
En3c6/hjjCepKWQEHEaPCRpmTOXqi6AOK0v9W5MCgGD/+f4Tgc2fRA4L6gTCg7vI+oL8ECKnV/M1
F/sjK21OG0tTwafNoIV+Rvj0jFGIgNfO9cOJLhTOp33FkZN19C6Je2xGEMqTQdZa+IjbS4laUFDt
e1i0Zbi7uxdFvz4OA/kA02DsFM2CLzBggikUJdIjpv8X+/FihUliv2Di7tj7H8Y2xNu3fu4bryKe
UHI0eC5NAacyHBquGnpXt2DLEpq3H+wghCQq6LYVG6+kFPFIRUrjn2NuCa/aGYs9VoFX0Q8llZif
tzpcTVvyvpAXOA1muKKXfTuirQDyGtdajUo5VTLJg21CPg5VWcILZmAFSLdywfHJKCM5vLM1U1DO
rJYOyUBeSV0kBf5+wS4ECc4II4yznk90LgMO88/k5E0wSI64K/Kf8EIIFjct23S2Hk8CQx0oknsy
gKSoRgnEn0PPepBbVC6kdutnt1sG/1xOmuXQkwuv3GJ3KEXRZaQWw14IM3mbmLTT2pKA12CB6ZLb
kDbLhwmYgXPU+Jrt5cbff0xTZYdnJMA9PvlQTQlv4yZuD1QgRBdOP79dOzQ7WakeUr7aQvgkb1Jc
XSRtCMAnPuD1tAz+vLFVljcEcxxulNUQ22st42I4mEjQesi/OJBdNeeaGWVBbrfV06hQ5jnAGC25
6cGfMd7K0K4Rjm3LNRMn8ewANoGRG3p8NiEmHcn9A70tXvPhu+7GBVIARRVHbf4BDiAQ68ndGxnB
y4PdQjF4gpw0eIi3KTcKB8lWHRbjkMu7pWM5qEjyyGZDfKx9u3i8ASb7iKpeX8lor0R63wL9Mtf2
nrQdV15tWPQKvTm8h7aCkvwTvivPcY5rD/PCtP/eQPRvgZAf88wu+ajC4ANIvCD+PlCBgA7YTfyk
sTGo2aGZSxvazKp6GQ121bC3GuSOF8j2qcSzVoNvLEMkJvE2muT9zaeFbNOFO3gz7i03g2Y9p2YL
fw3+ljJL8aGrNMoeUDF17D/M6ZqGjQY5/zYfsOhXO1WYLVLE+e7Z6wUjEN37YhR0V4rAwAmu7BLq
DArrs4nkFmrPDROiWgPa6RK/T4zBX5On8b5vmyAahvbht5gSLJdSsAQ7wWuw3a2pgrJlT1d46gWv
ObBsWSBM7DYZ/0JFFALA7dRt6/ovSLIiSzddtFuEoytjzhNZv+aV0ol5E6ZIJO+/mbD2UGRJ+xgJ
SsTg19TIiH2pTACmd4uuRUKhL4bK6Y/bmzMAW6B9Yeh0l8IAb/7h+8DCFaEzToF5rS7d3tVQgyhA
E3lHEPEch3rLIXUw5mYGYUmBVLIL8XSzXMe+SXp/gFJc/Iwf0PK8EwHsuFgYrvJ7xxgGlSlx5oev
xxNWl2AZH1oibV3VfdHv8zkMOkDQDz6TbyYQV7dVwNO86waZT2oQQtgOBZUK/87hVq9QPmBdI/Fb
+IGBMDAQ6iJHLswjuSmN/GzYIJ1EWyIJH12Dom69Z2Ozb3yxqih83H/l1vzPu5f0D93NTFyYZHza
quorQHHn9sLF1ZbW1I2UUOfoRTKpMRT0Wiyox0yHxfTZspZ2DhlHXohUog1xfsaYbfD9UnQrIktO
sHaacSpKqgxuVMhd9R6VHaNnjKdyg+DwTFEH41P0cF+V6YDZSdJIU5TleWUPoEIE2rnXhgMHU8J7
NwejZZlkt9tQM1BKEWLkLtS5kG6kRtclcYw04xLWMTo5ioeKISoHuQgPnKtoDDLr0E0+7Y25iK8l
Qq6e0nhaYauT8Qh/18viUQu7YM5LXT3eUAVBz/pSI6z7tca5VAxe+sU6iWpKfhg7PfqbAR8vD9zB
e+XFiqxDaaSprkHbuuyv1t5PV+XzIsH9pjE5x6M98HYY71Uwrkgc12HdQK4hkpK9MAXEVDF3mGM0
TyysjSjiuE6OPhSy5001EtawA1qy7je7uLh4Yoe0MlPwBiYzAmfvt924jTMK5ZDqzwXuhvuN/Ia4
aqZCaNu384ypCv+KGSEv8Rya5feNivu1phG/Gy7EUVZvCDudWiRYyq1YqpsRqCXWFXzbvsqAca2K
PVbppzRMU+c60MAAuIm3CGdB7US4SVraQic5brJb1i6FdzuWdgkscsD1SU56iSXgIoOW++CxbfZC
GJktsWx5oKUfwIyZar1xwaEKnB7qOsrO7zXzWo6/7i9ExFAm2j4NEmgSqM6kzW+HTkd+0rq5Ijwf
qGGPBPzFbQRd+ETC33IJdBgXcXZucQQUK2eV4dvIYNUBsH8UQMcYqI5aWPMMvMgbmja1P1bGbxPD
E2b3KTZDPrYpass9U1E9l36zshUiWFXv1HTwGkNt0ducsTfVCNFAQjl2Plp0Rqetm6TmLr+VuAzn
/km6tAyHu4e0G+6NadfiriOi0Y1hWwFjaB6wO1fFjQKPaXmbPTYFNghvTtZwoNMiW9xdpa/bNX5S
FYUGesGkcZ1wrKE+iC9MLQWmovzwc1aG7GXJZj2J7XL3M2laoN065NzM3wJUcFbb3ZJYu7AjgJ5g
JK8NYp0VE109Pzvk/5LeYA1qSPTOz41yJii4n/iLiEwG1qef3/IgAc4VFar6BTHQzD0C8XZ/6/cS
wt+tl4ff7CuOgD2AoqIeRVFmlUROkp9B0tdcDTLLEcXgwpwT/8PCEUQsmS0XrzSdU0J/Hn60RGH4
w7tjxjvgSHb6ld0Vu947rnFqNANEDrjDc0qnzEi4eYCZFvDpw8Nc0FX0RI6YOuRKicYJAX9mBbk/
8rArias6XsPfnT9zV1alz+xr1+fNgKlYSti9/yYIbI99WjEcT3fndJbkpXFzP7yReSWgzjxoO98a
szuyatNGxpyFZw68A4CrKBKan6c8YQwN5oIsxk8SohEveYglNCQwDzy1VtIwurYL5nWZuCQ4/06a
RMBZIABoVgHAIfuazqtVfZMYSW7poyqjSBG8ggGuEvsmW4kP/fn1HaBXf4PaN/qIzpyQAwaCStXx
z9IDdOxxKP3g5hc004lATHK6O9YZTAleske0K2kRM+MKckYZ9SS0KBITu80lBjB5W9GtcYohSDz6
ssHGQmA4AZ1Wr+bF0c0NLgsXJYCvU+Dl+Mqhc0sY/hmuJhInpuZ83Qfg3plIgvfm0k5/wbPHYpWO
lyNmeb6RUk9mxhU5sC504BScIpi2pxz3IpuQy2YANcRcwABNfVtDVvQHmI7lHaujFGAC4rK8wc73
KfyfQGqVgejPO9KQ9kB6Utf4Jj2GQni9KXrzEzbyxdfkHma/fmnISB4hIOklzfIiEl9YiLva6JO4
tJCW/xSC6F5mIAIWRpPXcJQnxYrIOiitrS01ALuIHBjHSCdpwiQGXy9DtIRGGIAwf7v9i1anDLi+
8I4DlTbiolRaC8zVdhxBqgbMMzbMjIdsm3q98poBH3AVBX51HMCBSk03KPvEOsZUYZzo6ZPEPC24
3ELeS8VdK2039B1PGJjehoVlvc7vkGrlLnZE3BmIcAQ0srx+pVZi//WReoRGWGeGkYaCacsl3Fcl
pIGo0GiVWdfbh5lbahixD7SrmwYXmdtF3vLvMxg9vYW6I/wENOTxUsgFI0sSStYLMZ7OtllK4N+f
fPwudUqRoKI55t6RtflpK2yoJzVHy0ZkzlRcDHlPsmrTEJE60Tfgx9/d4YZhavu7CnLZqi5GT7D9
3UEeHkS82XfKi+6lQia0w0Cy8DeCkaGxCBmQ6xYR2JxhSBPoFKMEeA8wAr9Ed/olbqNrUbbGOFOh
R91ss3HXIYU0SPPAY2DPk92+39Dqsbjkj38T2mOlw9vrp72YTa8wCRj+ByheUj1TG+9JLx1F3JGk
KLd75MGbVuEMJYHPyJ+kT/LF0lLGBXWnfIrXS5yDMgz2IuQT3gEz1cSL6BvazHVGO5xS0xZ6GmWK
fi6JOHKQT2pTjOtiA8rjGvjt+tEYVOxcXBD31QfRkrsgiTAX5ej4YNcfdC9a+/FZXr/IaJiCHzMQ
kG8SzjaMikuX7/rUOsSmRzRLbpfg/NFizPm8L7+DXk4V/wI0+4Q3wi8c3mjA3DWMWwKM6O2Qx8HS
2kNkgHxEzBrh+YOicAcDi2Qbp0CVxqpf+50VT9oOwz9Pm7wm4BEosDJJUiFQckdyLIbpROEEdYes
4JVh+3aVF4LY7O9uKLdsKU2/LhUNyF2JO/xJGTfbMGeSudWUpBjDGWdYkLhaPwP6cPe8Rp5ZgE7J
NpdpCTRicqISCe/ZQEoNfnGOWPjPxecl49e1o2/gMadRR+zbPRkcGcixck3dXoHO7y5u2gOLg4Va
eJmfWgg6lpkrMa2nixokYYe3MdeDGAwUdEi8GR0c7z7Il2LqmnOWzZoDoa65ESH9mm2FwGGpV/ck
ToH8Be+a4CfFJLSqVtRp59N0KnIPhPEXZCTeIl7B2tSUxjxdAWFKxbaljTTIuwmQT9HiZ8VpptvS
ED3HphIE5CDDn+SNoCRGbxLmKU3P5qnr1sMZyGqJSb7go5Qk1fkk/txDDY1fQ7YsZVGG3qTitxVY
VYoU3qDG1nbmBN4YI2H6tKx0k1n6WDVUyXMIaWnrAmuX+MZ0+0c1QxEKwuhMbpf05mGxcz/9m10o
2Fpwx0SyXa8G/uY1Ok3yOrWuAAR0sw9Io6vQ+SMAQvpKUdY/IIQBVvrRLH4IUAKucIdGqKv8unhm
KrOry8UIAyFfYV38TEh/mCH1Qdhvd4nN+lIX5ikvOyz48/sTJB7/0fGgFktQBPBGtU5XrJP/NPzj
+/98378buNF4A/JZ69VchFXJNBJ+QRNWmWXMp+5bEB6/TuVgN4APyP4BGFMCuDB9KWEPAhJRXtMt
jh94yvmFzwDp6cUhC/df5UmrXe0HtrliXjv3Ue/vPmEsmUeIcMyZu8wRs93fX2qxs5V0t4MmbBm3
/hTDh2oiFPC7kkdnavNjTisZIfew66cAlnVVgD8b/jFxE0IT+tsblDzVnbPGNMyNdJ7ZKkBnq2Oo
ZoWmwokIqhbHBN+1sqS2uPYq5OjXZUL2EfMILhYNA3jUgaX/4ynxh37QXarSGI19EzK31wjHDlHk
bhWvZnfoZ+A/7frImKGt9qreRxKpBYa3QsL+N2qtL9gLZFstfU4MlavSbGka/bDxaCsCxkKm+DH3
BuIJqtB7f14UxsEiLl1IBRzzwrJaEYU8T9FncUhAc51GNn6MHD5UfEETSAIx1pi1RdrFawxGtm62
td/vLn4BLMhrrNZ+jDZuPJUxR5PYmtoz41Hnh6dKhXsorpOF1jJ/KFzcbi+E8Bk0a0ABgM/XG8eq
rN6QtzLkxWxfyO3KjA1ZfYTjC5aN0fKolQvEgpb8WvyllmrCuq5L0+s+6tXt6fXNR8kyv+qCIb6e
eQgX/Iw3eYgLqcDiGwqRJjPcV2bOU6HcvBzP7D2f8yQr1KmsI8hokTakNeO3MNTmCn3g22rkNgVY
70kvsGDENe/Q62b/xlvF4o+S2Ux2l4tsPpAO5zYJR2yqo/NhuuQrwLqWqO6PUxb0DzsLpBOP9V7O
ztFiAdQsiBfzb9L0uW1anKYZYIjJA03V0Lwlkyx8TsZGcD2nUS3mvIwogbNE0MDcNxYL8jW011NO
cSt8bUrp94/vnMjuAMefQMyfdGtwxSXMAMXN+GZCm9VqSXP4hASy7NtHT4tyxhaU2fzRG6YbeT+2
pljaIhbKtJ6B6k49SsMGWK1u6YsqDHtpAYchwF01qo5arQr+hEeVFgflDh3i1fqwKGOkV1S7UnfF
SrZwIHZVjANaLiVPr0NyZeRPH6vKnLfioQOU4q5aCLotJQG2iBDvPNrmO7cogy7xVxier2Wxu+Tg
XBcG9pBYwPxtnauweWn2/hjZC8lBbJlkZ6qvZ9oT968JB5zN8w7Fw+VnPIPkxN8Xn01WA0EtfD4S
JvGCqXtmgLP8BjTDgiRSHvc0qcq8Nno4ZjUJcEAn28n0HxEF6S/nKnjz0cw25rZoWXgZiS45wyOv
Dw5uu5WT5LFLxR27JzWle4x+ieKb/vbAgdHxn2pugni22q7VyY/P0ed101zWU9O8HEk2fEIEHuX5
4NMUuIWa7PMBscyQm4Fio4TmgN0/2jslF5QbJ1GJXBPXN2AbLix4y2zEiUoQJBxePL/CS5O1icbH
qfpEe+hwjP38+4wOzx2yNpHMG8cuDA+V7c3+8PIr2n490Gsk4EJmQsinfsHt6IoaZ8DafkV+Q8u1
jaw+CqcGc+YlFNBQSIwaeYlGQySKv4ZjmUHKOoTPNgxW3dJnX4RJqoJ4DTeqM2ItF6LjQnpJusta
wy9yzM3yYceZYLZbqX0sKazxs3sN7OsDWyNb5W1oZQEm5tdyx7pko19RvDqAgn8cTT5mOVgRnAIp
BvUyNQwGPQLkoEUWABy+2KyFqNZpdcQbZfskf49g37usdTz11O47fAsP/Ul/WwjwDjjD4e0Xu3eQ
VDhIXX3iPjiJE5D1R7AaObzJ19i2DCs/wmYZ7Vd+qzz4aFmAg4oZc0gCsJ3lyItyKogmJazXMtNm
4UPybMsimoMC/TeXVXufmqlDqh4bYwifR+O84ReX2h3Ed6InjmfxcUwsqpYupAjm3olaXIcj0xdG
pr6NkqoRpQ54VudvYpTZS+EgYjIpFxq9O4GUbbD7P91srP0DakhwroboRvl+aeU+Eoj+gy28Ww31
MQxdnnEhPnT1GqSu1lbsaGjAclIn07lQdkc6yCLJh5SMuX7boA+NuGeQY3fLlfBbevhIqA8Tc8Db
9MF0Yv0GhivT96SebsPGy6nSPYvsntrfNNloU5Pm/qmd+OkJNImy1D2eseO+QEr/k9FM/Fq3znyG
/9pW74s2XN2yZIC/YjUhenKCUk9/45gTKBHNTauqR0qwwgUQqedIkx+sVOsSdv7518ZrTNBJf3n+
idSR30GUj7BKsUTO4Jvubn093jCPYCuk2lX9UBC720QKsxgrGfJbpL38wuQD/+fsbE3yVIhKeO+9
pK+ElO3rVYboPJLlPoOxxG+8lgiV6zHUkjK72wi5ELtqZKgZt3XQO39v2DqFKCb7zqSFryA7yBco
fMxbb4LJFf9/4LD4QLA2T+Kol/6SDEiwB6oZME24Xpsg4XZMm83Up70/vO+xMVpiMlCcKs/tizm6
bUnVXxwlrdWkdyzO7ej+QIbBxGfOHuPT/2zc+xXbbiZ4pr6WCqJBpk7ldAjEBjDeYNOe1cDw/hIp
uHt1KIqZ3YnCZTRDcB1zQySrcKp/hIZ0W02LNqYaNcs14Q1ex5vGv9JE8hUvY1F7I57VJzXQpHtC
j+LjTouSCnNepN+lilOe/eHN0gRrUvXlVmjJtKUmGujBoePnSFWehdkJwlizVs/IkcnJ2YoWcEv1
LtUjG1BYKa7YJPaE1rlxtH8bbVjd6ua3qUoMI2UA/H7zN7Apa4fkK7kbodOlC085zOv7S59qWY+d
dJ+b31P/dnLzsgca8c779ior6ultok6WxPhyRQx/LSqO2u0xvRyoAZHuJcAfwk4+Cgt1fvobLj1h
QORdOomOV1mJs3i8/ytK95h/iF4POoWEzUnrKe2OhrSO8+hWLHkNe4y1RGfJxbL8qKnkqLq/T5Qb
o4rncba6U+nTusxht25zgIS6jmJmBcIVjhdNWtGGD8MQvAP0r6aEq79EyZ6LBqFIwo0HVbTHXbwE
kOr3e+nKW+JHlc/wONJsTlnH3TcHdk/E8NqdlOPJsZk/EC4cc2o7Lqjl0zJMOlTld/lFn76yRzjp
HtNBB+wBX4B8/qYbQKzw1qjJFp5AHRn1djPBSYJ3LdY3pKdCaB1H5vS8Yf05/BHGLxEE7K/Ph4Ms
MVaYjH77+rPtjcNwSoztwTuLCbKODrhiOBeM3bMHEwOvJDbXo19sr4QTIOaNFoMxTRuYbXjv6/pH
rbrW9ka5dKFDKq+At9CwQuUHh+tjNtk/DHnaABOBH9GTQ0JcajmSQkwWcmKvXIfgaep+POCUk4qL
54PSc3AD3NGjoBfY16V75bpY9YC4h07TUbgHjaccxJmXkD0+EQKbhKG8GnZplFHZq76zIwedoL7Z
mJSAor+5A5Dehw+/Bt37NysMx4AeU+DdJUnv11gJ99TOimeUZQv01h10m2+uzX0iWHyf/6F+reET
i9C1HkhgkpjCpsFI+QiV1MOF3q0Bv9Wzx04aaVUsGKbS5ne5j9rDZ5uib/W4WepT+BOdzRM0Wp62
XVERnVG5fDj6meVAZptg5mP9YFf6XPZsXqyBRNQcrpWIN6yfGEGfOupQ5QKiMcGiQSYypJVSVC6C
t0A9zgKHslu0W55CqlmVi81ZvKe1Jex/+eHTqHLpbBU+d/m+drKyFZszXDggj2XxlBVnHiGmxg0P
uedscOQZ43r1z402edeR+wlxX0s8mAAIt3Q1GKFw9vhrqhOlaOLFUf+cqEm8/59yT0vqp5+cfP1K
tLOo36k4+xbYYBVFmgtkt8a4HL3cABqK8urIb28rhqwxQQ+t8kChmAHMN+5lYouZi42BRZyP3qZE
ADnIJtqr4DUL2ZkDUchlUSJTisKSreFJFLs23UmfWLtf2mYsN/nLSIaIAQz6jAgWNWdN39e6einU
cDEHtPO4r4D0Cuy/niIeDS+LFlEhiMDjXI1YMuVhhRtXbT0zLduIxdOFfGgUCfJHWG0s5XxSlCjg
/kHYnU5Q4XzQ3OcFaNrP2JpMV9oc57anmP186z+bq4AV+hOnmcYC2V7XkFZ1WcbllSClyJgwI56v
yIvSk4pmmbKh9OJPei4pJ74XDd3EQWEXImzEvxScXdltFRd/8eocJrTeatKYtD7veF/2wSzI+0wO
Tx5fXH3kRhl7oOWDAsulZ4OpGWYb0Bxnf6VbMENQqtQgFV8sq/IqIDIBHmZuyCl6Ew4A5XeysT4W
pc4Gpm9/y2aj/wT4K6BO1hulqiNzpx3l3crqRJN2nlVbEYVih6EXRBVViZgDyf7XTSqFL2a50Anm
5geB/27rbYUyX+f7dk2Sf5HdVlmeaQ7+autOaBBZqoebm3HF4ZpJ+eKXoe8f8wfVSxXx/TXzwQND
i+yeMFtYUvRcX50gHBfHbB3KshZoS9JIdYRg88vpijMeXhVdAjgROcYC24XxY4Ja8U5l6U2ddWRn
+vL5E5tUkHN7TCD9VX6aQRE3CcZV5fQ2z70Oj9L55EPq5qHyO+5INGhKpmrHJcOlBue/zV+13Fp2
MzlmMoteCwO37HRXusIbEM+1FyNijnuhJKQEkGDJN76odtS1dM3VAkGXMMtr/gYGOLGS9iyYaTz9
Z5XDjyc9zC7J5921Ji7Zv9mOICFjwUMBJQxrHufsyAnuIYTMJ/mGSd+0mNyCMpZcFBrDDA1bvJJm
72HhR7292tpzgRXi5r77RH73cg8HLDHZTB47mcqkIUpzQD+vqnVZfZXQhyi0Hq/0pLBfL6P3/S/V
GoptEe95QPVPEikEzg6EPHuzcmbhXohtnD4QXsN6pj87/QtEjLTQqPasWXOOI7HZHWYVHel2+BRG
DxVhHkDFlMn/ROgrGGeIjl3OjX4yaFyB/Ba/57Cc1HqpFtdM+0GbJTcwJGmk0B1o1WQXjFstrZ6j
72Y6He9TfLN2uy8BTQYCGKMgu2DipwEa1JUK5mpQfT8K+ao2iWDC9fIOahm6IeUeJNlgD3KRGLyn
Ze/VmCbREnjcKCMynAqK6foUc5RwTZOB+HrSFRb43EpJuzoKczb1xzRtIhLIhAGQUeBKp3r2xn/x
T4PHlc1rYwbvODZYOSwDp+xHFgM5pglEdVgQvmQuyKQC4JhiUA7VzSvi3+mE9NOHuQ27IlDNGBpm
f8v+XYHPNP6TycfhadjV6luZaMpAEcguWjcRknYi8+/aNssR7O6S3qRmZfMAB3yI94GZZQ4GkRAU
8VRAUUAumGf2SXGPoPk+C+VKUnrghG82V5xz5s4SS6RSw6TYGyRFEYz1Q8jMnPNE35qZVgzxtTsd
YuSKrm1HDm8P0CoNVxUCO/KhT7Qi9e6dcfj3hQ9Xdd9bMHjIYAEyskHcwe6wVc7gUmmyNzv5OwBB
PiuCKf8lab2O1RmLUYkGD+6190yLlBEw4TtqK8ea03hDCXnqHJ3KQX0xC9KIkgZCyQMXnG2e4XY5
YSfhe9HLpywc7nAImPIc3gg1uLpszDdGRdu36QuuWHnzmawhFHArx235Meo8Rcux07WbreF279F8
LnkbKVTbqHyxquoW3w5qJA8+rQ1b9p6Gye2aeApwqg3tbSKgWL9HF1cqhrOKmblrmMOQ2n3z7Vrx
yPUPB8tgm2nFjCP1CDI6Xa79DJBKQcolfoUI10p4KRmlv11D18bS0VMW+ZWD2IsifwR92KZpGE3u
4vYqifxriNWEF3tobNub1jnGpiLJ9cx4jLlTEVKbIgTamu8ju0u/GP0LIc7PnXRizOzaUS4SmmFs
as913JC/LxTZ4anblyqcqb0rXXr+IadC6elG63jA7n3D8jal4tFv99/HcxYoxtbAd7xQGg9Jx/QM
nq/YrR/ojsJJkexmYUC25mB9JMrZCxbAZkoI/FD07pBXpbK6TcOILPQq6SewCgsdG2hS1hr1bM2h
P6/DTG70qCyHsgcB+AtYBV6cmu62lsWf635xdOKA4C+79+kiExiei3jJCA6E7g/N+wX+t+SwciWZ
CgEAkM33IYLGH+2UJdxN7Q2M1WmlwUZ2TyUmbYuXdboyV7DfVq6QlRKVnXvMGLDGur/vtRJyShju
Jca532RRQnLPyWqyg9xp6/ZHgRRpIz3k08HVO8eNNogOOwPz8WhaJgTx9ycM2+wL+bWro3rPcEdb
a+hs6IvBffMIe05dkReHARS9tLK1sjUCDwC8osqCD9s2PP0y3ZCkvqm/B+l5IKIf2yasK+YXfp0L
P6D5kd1ZP5dw+T04eEjnzjsa6q3YpeDL3pfA9uhmLrL+gW68glqR5WrWlU9hECdOTC2cg69tmQ8s
ZPABPM8N8ZKA+gihnlYtpkBAC1w/yOtsmQhAJ4Y8zKFxB/VvFOcbmLyUoABS6xAuXykN6CJq1iMj
77CkJbtrdlR8dsesb2YHEnH3nfuIwBC3eZZnNjKlye+WM7FBoCz0KsNwGThd7qVcirH79Y46AQYz
yIe5EiCxhJh4y9AV3voOYReWRzttSYDTfz6+5Y1SZEhnP8lCX0OAjasa9he5r8No5hSYWhEmTp9z
C/n17iLieB75sxXQx2rhkMbysE24IEXymF9h0O3sAe8O5Ae15p5ARQfCorWCxEN1ReFyv81DHoJR
6F8VxJiT/WM+xXHRNM8N4gTyFA8LbbhFF73Ja02fSFo7dJaewTq5h6B3MCiHfMz/QY1ZQHFh+L4d
eAuf6mUOODHXhzTEPu7ThAjYfalzL6lF3Nz1OPxFa4eubqeyxFx5+C692J/XwIJTxRhT580gg2if
11BtUCNOmBfqflHAmzMMgbTKaHnaiQW4EUSYvg0jDDiYNCdvCVSrZGoWFiOksDZTYUuA2sZ68FRt
s1BHR5h32Q1IZi4SYTDABoeVnO/EH8mSkzuCkjHQeZMhHhHb0uGIh6x7fJu/wqHKrwg4GoLKVycP
BO250kScukyzDWZU/M19NVKY77vzhywB+Dim6U0QmP5ZhZCXy3W1VKi6mAC0YP5I65PR5E/7XFnl
ZBFo0743GypoYA6xmu8EPCMOLHvIeXakUlC7Q0TfTH3hyQODTraHDL0ZeC/lvpw97SI9IPy9IEcv
MvTOrAJFbkT5IEI57YXR7ExFVu25ybfEuq9eL9H/0b8HDfYMVXJCJ7veXGPbm71BoCfq+/iglJ66
AuuKZY3YM2k9e6Z975jOuYsH1NJrbxx/PfUchmJ54gR+4iyvzK2F2p+RYtHA6UWvsvT9+2kZdVPb
0ySxildKTHygN1o/9Nk81CjOl7cFrarlo7mPOUeyEEnSpAqvb94/iqXbllWllU4m3PrYSPvirIvz
F531yx+a7/23Q3l8vykfqdY3o8Gb/0V4ybOCVqiwUKVXOP8j4fvzTv2buMPFT6kUeNvx0ovVMDpm
IEMK9uc86MOcEnjCMF+80m+bZO18EL7im2xq5qMDWqM4jMbapRDvLY1nYOkgARh4SYdjiHgOykS7
TRXNWl8z7Qe50tH2ueAKdQCQheAfi+hOHRHe8uqO1PvXGKNxL7ZXC/c0I1wS2lNrKMTKMYTvH5VJ
+APSSkjCDAxoL6JHpcrHDrU2kITBCD573NXvqvSaPL+hjb/Rwap9uZcVc7f4+RDFVYGgRGOfVPql
NL77wr87v21e6cs+MFP4cMx1GEUfd4XJ3KkmKOWiQe6+UhqS+ZNoFnJOMQ/T7qGfHUgt+3HeVcXn
Zb4q8p22vwsQs4d4EQ7jCNq5RB5lcYA3nMlzcfX//DjRtcDR5CSbr9jCH2hVrBAPMTkh5sycNTBa
ys3WbEg99Wgew+wNIf/lbVCCOzgY618bt6yiZg5xda9chV+Ua2N0DWZm5xtwBnwlrL3bkIgqco3p
G7KJ/jRcjyQMTpLTC9Hi2rzOJqAXC6ob9OpAjvsQ0VgiZd9qsJQWbeT+p/sINNbzidwRUxK38i//
d7GhKOgUtciGXxyWVdhvVGjGSUYNhJ5kcs1PJihg4+hv/VElh4MSlDNgQ3RIfSd88FKRe9u7eEMF
PSV8eyC6NVQ5h+ATphNzx9ZPGA/BBB2zIX7Vo66K675nMxHuurzjSm7rws4v6FWXzF/VMq+mIBy1
kHLOTHF3c9lP5GqyrQCzMVj8xVBcGqYf9j7rYkOpQ4FW3FX9+2Pp+Pjle+0s1rk5ZRsKpqDug9BI
//B4iZMne4Iy6f/TD2+1UC5QBFtgZPS4NtoUOCP2XqVYTWu35PEP49PsESky9kOk7qDiWAqNtVuE
JvKthSocpxaaqXYet/SnIOpSDEqBxiSiBRPrqttjh1/e9/WgWznQ5ICDieeV9SuTWUqjpNI5RcAs
R25/R1iRh/V19lOG19StX6VcZIfJJ7qNtPXdKHaasjc1MjzTTHcBEa1Lbz3b4eifmfY9mIOJjLuR
3lzvoFJJ6YirRlgAmN8t22MVdZ/Vzc0Sj0U+9ouPOhDd0kLf3NzLM1bW96AkP+QTe3zpgdsMTsJG
LiMRwSofuJWvsO9/Uos1T8hHvuYfOWvBg8SDRQleGvbEppnuyakUEdjq3I7iwxYMeUFSDCNKgzqN
UlW5MS9y1Y9jKLfWCabI6XogSC7N+h+HlccXqsklFokmcn8+tU5Ywy9QnmOzzy7K8TmKpxL38EsP
MsV1uazli1I/rh5iPvco3qfuXOA5yasI6RKb6tb3R0ymW+rjeNgne6BDl5jkaVFhNMsruFgBRN7w
w8E5f+y/giHPMNCeZ4TCrZe30V/XSKEenO/Icjicgh4fk1kd2q4hfvW3TKT4b1Yv/Mk62YTSEIhS
r/sAht93Zv2QBSliMkESh7IKpXTKK4o76J5oYIKQ4eFDHXXJofEMGxMZHiyqCg/1dsoy3OVLuEFu
y2MnzxYgBIAhS13wnByVPD6BBE2augl0/VsRIKDWsZJKKty8Qz7QzANPWAeyhuJk8OjgJFqhfIki
Bz4PK/IQpzfNH4MHJUJ4mXfSLhh5KM4xI+I/nTcXUbyAjc+CFaLC4gYzfVIJleebv6yIyQSSqR4k
iSAS8nKlrd1lqGJN8RFsgPwOp8Wlw5lsbwh80XFx/Gx9Cj5JooFPYIu6w4rxtD0MYMV/2wSQB5Y2
RLBbxCQaKactvya5WFwgUg7ub3gGiJFhWJGC1Q/38b9NOxGA3YslIafPsCQhpE+5Xv7hhDCs8NmB
MgDxOjps5pfecKQ3eptB9E8+IAa2Amyiw8u0of73pQv2XFFMR31+i2zZ5GfPnqS0ZlQUOU2Mom9p
M3SneFwipRpyZkNqOS3MzyUiXoZ7zeqpl4oDBqh8qGNAySLmawKAi4NLMRdez6XLhkXQd5ZY2cgt
Y4lViJ4TZfPbDV+lPBWSbbJwDiMDGwHh5B8dXGn1BhWNmEfZ/HG/0McmQNIbI62phuXitj73L1Sc
jn9de5yvu3JUFLH5STJWIz/uc6YigiSrZCVB6XFbW9ZPY24H0bWY/4wOjd4EvsqITpfAteB9IATn
q/PklUb9EpZTmwmwZ4w6gILfyIDtRTQ/6EfPtTRt4XAxgEYLQctxCg1j2OhR8j1SVDfHb3AgOpi1
zUdR5DU3Hmw9TBrZDNC7fpikC0AjBYWdD4Oe3DWVhKGagCP8WDxdhwj/EBqdmZrlog294DUFP+bk
Rj/Lb7XgUYydBz+Ofese7zpWYcqcbIyPe/Php5f/TO1/l0YmTqfTnjnxc3o4nq2E5GkI3DT1cJle
1jZmMimKgEPsLDj99Zs38Kn7XuKkx9coxbvcgEaEldcKBSr5gDhfv/Wcl4TPA/ZWujjDDxWgS9l9
hu3G9L6CyYCj7ulKvWlmad1z1FcGKZqxxLie6irw9pQ2nfopVEE9nTn+/+mxazEzd5y+FrfmXGYk
HClCtfr/rguz7frN06HvgXetHy1FROCt5L4ykj1QNmfNA24A1L4P9r1oaizljq4RqulDqVIld0sk
Wm0tYf1nL5xZ1jYAXJuKWMxTqsIX7H4xXrdjtzaC7oc3UwY6GMXm0sgPBndDAjLqb80a2fwbMvxZ
y+lj9+77ocnLcFOCxnk1naiYrebTd57+2Hdx8Q97yn3usMgVx5SChFZ/J68Sn7TJRSV1FzyVEyBb
hZ8wCBdtL5JB9ddT4P/zKnW4YfgoOzBp0VqYnKB6/hRMaFHdduj+/syZnPltYO8IvYDHYetLvIP4
b/XrMFQb0zCuyT5WzZNgpyKOQP+xx4TboIJuAdznkvhFVdZ414M688iM9+OKuYW3LN5gPbkAswY8
ftMKlBQkZbuocwEqUPKFEKAoV4fwWy+iVoUjpd7h7Yc+AfGsfkn5JX2VpdBo04GJ2SwEFr4XzqJ3
076/ECAOdNd58dmu5w1PdC5Y2SfGS1+icgfrn4+Q+OhemQZDyl0hDvHVg9jplTK3Rli8RiICbzBF
evVBxdGEbk1iCAkiGLyePQB1c3DEz+zXu0+lzFOzq5afMN+bnU7XB4hiWC18iQIYBsuHeXobJ4HA
dvQEID2Y/Od7IslzY2m7VrIistB9ra8/gxEH8vy+XMkd/wsvPsFlRLisUFrK1CyuDJ7hSi20fRPd
Ahti3vhkPJxDgwRxxc4pKGAq0UgfINL3/ralHArKmLrMFLT9pUwoMzUnleyjfhV8/Ui2ujtgVdST
54sPCekJa2rNPiICfbfbleySz0nbd7rhIVI37J3n3dAgwe1kD3hx8OPMHvamqQQg3oSzCWk1748t
U6/W7VF6371ndG27yTxc3y4NNkN5gr2/H6fDxrgu5dxUaRiV0xcxAV+xb87BODKrMkkZrOxpY8ig
Tfs/7/QHOkpGyFopkl7GEe370CtW7I3NKm1A1HThqqkwLAMKTSKhlAwRvGVPQp9gC7KVDP9Wv7FT
irCAETXsSZNcr083qWd7ExySF+Fp/qdfHm11W13L4OIU/3QCsWfL52Nwx/05IFWK1vjC5gasjD8L
mMiUULQOi3bG2NCwq7r88E9zwDO2HDpZjwBL9Hp/SX2ObqyoNn9TuIjjQzvdIxA+MaIjk5e9Xt7w
O8Jo9dkswNu+0m/RX4YAMaIyxBEBPvitG1fczFhrlYpC7flDEj8Ns/tK0Y2p/Ioyd8zk8D/cFDZf
U7yrzFo0KwNZI1iFZftNUpnNP+fzDHxY2zqgiZZvPuAhSrEuyhp3p6olTD+buDagl3xG8lIbrbYG
xZkx82sZFc4a7xOypOx83+QhXerYgWagSc7aXlt9ZU/MOlWxrn67CuX8yND2hh0Yqk7EbTUq9WgQ
RTy2PYMzoPPfJS5MODfGe1XDo5aRHoxgoi7XprR2ebjrQ3fwwCu5qLRKcAh8UWA453CQ6mMH8QqA
qrC8toOeuuIsD9EQZYd9gZlwtIgwvzY/PnKYpK05HyXBXrJHhT4ZoYcVuQvJaLlfKXeiuqv5guo3
lHNdtVC1V3/j73aboFOPe4h0FVrHJbeWfxjak+7pyD06JznPHyOx/sP6gzzczBNFlnfpnDi37R36
UFHW1L6CdZBUMrl5tVblzdblu3dioBYmj4fUZRdsDrTLIjOfHYLN6Sjj09Bp3/3D9fvPracVjT5K
zkrFogfcaVq4LJ4233A2vBdOpImArNefnjcUU3hhNN5Bh0fbETGyyioBADc9xdgX6PfDbyNkDJhq
6oaxjX2P8lWRG/d2bxIKe/YV/GKjvi1KfgL6VbVV1fItqd7FuhI3DfxRdd2m0r1DNrgRe4KgPW3+
8qZ/9zkTf7vZtTE61uNPSQb0FSncNnhbbugdjhMAylfEy4/hbwPQmvGHhNapBBj4NwnBeQUc7Lfs
1qVvVH2GiDq6QBQrsdbD8XhpICu8ErGID9eYdT905pVMZdyjlfyHN1G/DXVgWIucH0BIAyJbLuE3
d2HpH9w/1/a7tyvHC8aMTerZ4fwQJOm0AybrceFYFJ0kgKhE72NBgZPEynA3o74HkCAkPEv1B0rt
Sl8GD5OQnCZXxUabQ/tHedrE/Ux9hGedDAjiGh3pZfOqY3MkNmFkoT5JUxYZpxruheH/P1M08097
TLMZloU19KUXoHclfFrVzW0gWTakSg6+X9Scwpq5TJcdYoPfJG0p9xwI4vsDWeX4vMxe2ZDuVzBi
b0QYFI4X7do5yu9U35BSDqOG13lxoTXuYNhu9RZPGLVYkQfbImwg7Q+LNoKioT0JsWotM8XsL7C9
xiK62yH5a5/SD/c8fhlFXW626LIIWwiHQFRyO9Yy0V1Pmzk9hEiLd8mmvFKice+79cbeF+TcIhpO
7arbjcgUXfaWWjmH/KBZUTjt5EMVfjXxT3F5HbtNgsVdKdBJi/vr5w5AAz0VMqLE22luPgxDknPU
O46OHb9534aD0EJ1zpV4Rj04C9jCIOU/b7Nk4hnLH+F5G75oG3f/RLcq2ecY4WTZaJpQCtRxyLCl
nOlbdA1dQvf26B6WSMXPAdDnLzztL822SL/iZcJfEMFUnWh6uXXRwQNilvoDto9t5pJO1ekD/BfK
fzJCq++fo7jsN4nq/09K0/HASURChF7V17jX5FL80OMPIe7OGSltw9lcP+HxdJIKn2oOuvxg//Um
xETkkP73vjjamJuSFcyQZSRZgJGJYwH8Veyxac8sW+nGOyVButux4mdhfDqswGaFIjnIUmkZA2cv
IR56FZZS3WRPuu4rM93lDyzxBsmrNXzRobcPrPeKifbskJAVbRKgV6i1KMGgCgMWjyQjcAUaBsWm
FiacNx15xpPM348VHyhXMbgr1Ky4fubzIyajB0Ffa6L2/QtBf+ctCVHx2MRoXFoLypMXdB9A9wRo
+iCvmAmHPPN8ccCOd1lcWnlTnrfORm4xYlZmDiSTO+ZffDKvR35nbqmFc9Ka7o54RcRLic7kVPax
8V7+2ruTqNQbD1Maqg4BaeAhQl0i/XBQlpc93cfe8dRirVYERbPogUVIAIQOTwTzsQASjWt+2IEJ
but03oplAmrmP2GIoRYjx3t80YqGdgg0NnC4gNJXyhH/HWzJcLAlF8cyFN74Q3AMYTv7GapqALqi
HDSlYbmTogmQpffjKPOvam9pKPkHHotv3Z/mP5xf4ChwTJ0MXUE++I6TDxDgZurpAPZpzALwIvsF
orUFrygYd7rQYD9BVu4qr7nQTAXg0uJnNGPvvIs6+jJUMaTyCOF5ipSp9/F1K12/F75O7zxxFyzF
PffUKe+PkYxmL3kfoVabMLbwlis3cuqLcPAhWMlZx2TsGOSFrnD0kvBnNFkk8hBq1dOViCI7UyqB
RzbQjmsL7fdUo1rSPkIYxZtBCAXly6YMAbpg1dAe7W9IfIwX+5XWkw3VAJCKQR7nY1biVdk/hnSk
LfXwR2WLhZLRRx1PL7ruCFfkrB47npwGLMxl82aW21jhmUjhcz2VJ2Omskx8AMdH5p0iRQprUgxy
y6E5I/hRgGSBwB53aYJ/FdzsA18ZlCynCH+P5lLMt5fnmYqGaH+XChuHd0UGBczEV6y5dmvV84+5
+zBzJjKaet/CdNXZLz5Oudzg+dAGyiE7FEOryFRxqhNs/v3bq4z/tV62jpxVH9ekfZrT1B966lHa
dfhNsVjKRli8AZzwROptQN97c8O7TAzUhLzQaANcB8dj4vSY7w6zIzGPUjsJ9QLa2muP8gxxncGk
T0AD1um723ylpX9n4Nd7eALxAk57WKRl3akuqk9H4wxzXQqQKPjFztx1nRw6q0rJPZpSQSujQOja
5H74s5wOnseX4l8ET/+ht+Smpx61wyd9TZ89Z9nk3filHO1JsA6HAc9eqUNcOC1qnjd60PWosEgG
7LCSJeCisQ58X614IWjAz+oAqFt1dF+30vy++Vyk1zAjlCZy9el9IN23F4xefRun5AVjtn9dNGyB
i3cKH/BWOwsJDp1MQqcFWGE2JTMmtXRmXwmOi9nJWsrpdMlrC7zhxHB/OdjKiJIgUdAmMiT33n0W
qUUD1aiosJENm9IuQa249IVeNVUkqjMvf/XkqEzOyxqwnSbUBN66+3GQ858LGb3kPP3zZhL+NoYY
0YMMRPaAjDyeS2G8AyhfgTiDtaKwO8PBd+kAywtvSe5FHsL//YORiBj6QI2G0yRqdI1FAaw2uVh3
uI2qG3I3lpxArdxHaMIPpyqlXLJ/skacW9S0ugSS4PCmipQUtoPJCxZvCK3xraJjktyVgpt0Rwin
vRLL11rSz/RsM/k2SxYTIrDYT/YHTB29W5w9iMrLALP5fdPhNe5voVrYdH1U6FrCk/p+8wr7AWrQ
LRRGRVG/wLJdDC8J7qWZLOsFMcLfBuQ/AhYtcOOkb20RKde1iB5uPvWl+8WVFKVPxoMaPrqCdC0S
lTdGgNGpkOpZaVZJR6p4+aI91sGMnuR4fMf97+/xJClVF4Hs7WBP+GLoz3XjDL7gyvhv6kvRt7v7
jcDsp5VqgGd7wT/RYfMKJMiSo+ldmJ558ecLzZbr/torzobdfKis9eTENCQfiVw/U6u0KoqUIl0Q
BrAueIdru39ABvPTiPF6vNMWLgrjTBKTscVvceWyPnm39a5NIL8HyAi/746ccHRW1PzE9m0poBcu
mkvCJ/LvMN+9udFq5ft65UPh1LFzeZfjwtV5rDpdqmyqF2bZXnIWEFqEtbOTlWDxXm2NWYTozK9h
HSJL6MLPuAcxDgGFoM0GAz7q8dYXPe7BFhbpunqkaF81s2sjl8cFkVUTe3pMkbGp2to5NAJUDk/E
DZDBaZFefWfxLBZrXYu43b4jMo0E/isoyN/DKvkTbk4T61r6Ea0P2d2ESbK7UMWG+O8prYWmbY5c
iedYEYx1iRnehFYwftbp//e5gbLr0iY5mwT6frTQRczodLakrnxYqJ+J7G28LZUMR5ULxyRdDkUd
cMTvTw6XG+tppozEERmku3PFk3YkwlzsvBbmjgr5CMawc2c75a7o7LsgNLc2f5nN7c3CI45ZTm38
H9SUIWIEC92/LI8N+tDiDVuQhO237Yw7XKP5DioEU96PBKnNbq0g1jIRqm75Qt/WNOYso0Lq5+XD
Uu4qQYpod2cUO3ZR6G1OPB5r+oVkipLPig6Nb75F4LLGjOQUqUDficouKbKgo0+4crEpIkbbzuBo
HDcyKAFrHh6i6XawpR6/uG9U3jBOVYgy1OPsW/oPdodrEuG9HwebIDUYLp3lOgtzde0+bHXmGvJe
FSl19zc3bBTxgUs3Uy842ows9jEzIQyyq6TvaiY2YOPVtSQiTM+eWnLTercuy2pCDOgmq4S/9NnT
0uSY+FEs4u2oadSmWJGvqF2An2yJYKGXWqXZVfvX9MlShPCGhrRs3MIUdOmlzJOosLDQKpzSXJN0
7DCYHN8fQmadnGk6LZtBhqNutTRFAlXWDB/X1pW+Akvw/3BrXRK5XRFGUgHf9pGYNixe9ZX2Iu/B
/Tin1tr4ihw6OXrlrKn4CbOv/rtnp+/Bd2AkHPg+RiVfxtPxR6NHKNDrY62Mh+aGqzdIKjkr2sUQ
K3U3ORHcrtLJEa/I5tFhzAU6vhZq1xSQB7VPqrQ1gSg6b83FNjk5rMPlYyquWhsHvWYYjyKoVYds
BOGvnUtHsezyxZ9tmzvPz5ej7J1Nr4iu0qbUH53/DyZ/wFdOTFR3Kf5PXFbAmYXIrPaNJPoTOxz6
wdUvq4o2Iik6AXB+H8HF3gJtE5xzw4+U5Thz7mdryxr5ZrOOu82ZXA53K1K/dc7ZsYAQiGXDJ9Ku
AxNlAD/GOA3atjB2bCYqG4cjTs2NXFlH2/8o8eaFjjU5bQ5r4QqiORwiQBujOAh56LU0NG1yHgIn
HkfHw2nBZYLMV5pMDmkm7v7DuX/jdXpV/yr/+61N0s2AsN4HWL1PEc4xrSC8wg+yUQZ6ugdMpzQz
fv7h8TEWzPASrcovcJnb6HH2YIFSdK9hi+Y6P+RAMzAgIzKHagSoqyrfdeNm/4laEK6tCvE+4UQo
isZu+nTaAOqTRU5xzi0FE+mnVx9+cHxD9kRDQGeYeQIlbFkp2kh6e6dCzopLSQVVjRoff8YJ6AL8
Ggnv1vIuNjGlAPQtiSvy2ApQr4nRnEszhGrGzROb3bzEJ8kBIjcCHuRBLUmjHl0gyBMVqFTKwQLI
CBGHU24MDu96gaEe/+dUrM09726pya+F9mE96Ie7a4/LA0ADvqXsRvrqm8UTI3TRsGZu6EaDXQFg
JFsrN7dAVhnMHL0UWvtzlGYIw5M0BIrzO9mxRR57gK9W4HWcYLFuy6oAFJfYAVJ404mr/hwObyg7
1T3i9pPSUZRLljXzNfeDOFM9Or1yBMXSFD53fpmH6kJQFVjuovymQtzn4cSQrf/Ch/CGcpB4dcij
vvu1iWtfhc7WsEmJR0cdI2dC9pdjAFRG1NDRWIImGC333tHTByd41QW6LpVKcGafjAFb8D1mqw62
z5QUr6J88eFLAV3wixwCWO2/ahddH+x5GeZGo2tkzN5cfNsGyDukg8M3QI9flnzwnMVFlSSndBSI
wWoWcdCZsJQ3ql6xRsWH6+RtX6qypL/be/QJLkZYnKniA319tBSaggqlkFtKSxkr4JglK/qrtylj
dBnxg2mgad7krQtONsXrUBTqv72f9j2/EiyXlTSZBMc3rqQF6fhMF8PGN4Iug6bs4/mUNQH25gvm
/fDpX1/k139SKqjNglyerhdnk7gJ0tB9yx2c8XetR0c8kTzmfUtjkhE+dQ2NX7S3AYA2Qg+tN9Fk
UN4piLGM9WuN+zpN3YBkFjWKnRYT8ixZgF+l2AheEIAGxbqKIkkJHiCUjEnPmRilosoRPbc07NU5
0cKo5AulHN4+6hAKQC4Jt1XyNKzc4ie4//5/PGN1aCgrd81V3mPnPn7svgshgZYLVGraB9kqvd5J
oO7NSqbgLsC+xK/6XbzS3MJ8m15jUPmvlog00ruxzZZPwpf5ZuyFv9hSEnJ1qVI9Rnv49xngiL9F
tRE9o3ysduhNdyZWWOtfQgW2ifwyguKkU8U8jX5U4CKG7o6sET7VoSTovvuEuD6vV8/NaDe8DdF6
tHJ8Dx/JPF0IbtJeqs37bMz9uNiIJPjV3Ag87WJqXGBPDbI3LQrvBkigThss2VJmqm9LqmVBNXth
PVxrFcBlnLn6ker8VKBeiZuMEoGntILl8pgRHkWxTzIPIR/N+7mY2/fb+FmC7Qk/PWsnPzdrfICT
fZfshYhQffI5g70z2oZOluKfz8oSVJdwo7Xlzreby3B5nvYHPeaD4sGxiKKZRp9xmrf7Usl4522c
+XhgXBSwjUUD5Qu5sU7UeFt2JBE/zwGnm3+6mI2PRXqVr4Rf/dYZ/5Y3DLDUWpgU3VSpRZAgBTfI
MYQTUWaNl8W99OvJzu8uvAyGNaqE4Puy4qJ/EZo4DAgh85cnVM5c/ykoFTX/AaE69PZPejc63mOj
V2MWHDSIA9vVzTYzEjZoKRqxoucQ9Kp4LLTmlG4jAoMlIawz6uLKtz5YX/4fwhavZhuVT3yT2s8y
8sRSxVHqA2KiS4U1clBEMvPzETb/A9cXLtB/9Tjhs+AkqPifgnA3iYCAtuyuESAQmXdYhAZGP+Rm
4eZ3ceE/chFPo4sX0KzVsZv+SJq0qPbzZ1i+w+EnIDTnqBB+lLkKJwS1gBb654c+agcz3Z8mkrK/
mvM6v14z4w/DgEWyhpdEeBDE6FhSVrm3ioj91KESyTAXiKlstKNAFEI4FwXE46EIsDcYpdfoLPlo
qQ1a612BtZtsS0QXEILYuaEbljmvDp6C0L6tYuvfIZAYvjXWGs0pd6lYN7qvlzvSHWfFyxE32mj8
3wNsRnw9a8HPqJtog1ixAtBl3FCmbweubq8hfbcXGTAb0W+DE/39KkjW3jHj/BioYGJLOqEU7moU
sESz58bYzZC42DrnN225xGQ9X/0D2Gia5BUnMWM4f69RCd3+HLtxekzN+W3A3pEY6zo0UoBFy+pQ
F7Re0XvDyEt7h1x3fJ25/YOuObZgk7fsd9Ue1W0EGMGKOpmRZ3LxY8VCwqZALnlV9aOYHycIFvyz
Idw10+L0CFfqh4TtjYCX58Ef+/X3E9jRake6b1t1GEysL3YCM7rj1EMsiOxuX5qNu4uAjwa6lAmm
Llbw1sutn/zxWqkZS48ybYGxjGmBS+9EZCws4XzNH+/GEmAOkN+fXPDXMHInwvVk1Kjz7XYD2rid
Mses1Ds7/kauGMQoVp6TdDm8EyNIZwanl1q/LMLnoU7ASngtX6seEBJfvXsrpaMj+KTWh8v1JztC
Vn/3eSkrXjBqKReOMcU1RT800keYHBPeJJQZQYfIc/PFZZwK7ritk+H0h/679jLXpeVWt9ZbM++I
fqVVuh/2W6mR44g7DcOHJZn9lXUFn3bOksYxu9flSs27yvXun6QNKjaZiNOEDPDf44sJ+PCM2qa3
dJQe0HREYoyksxfP7v8yRgKgPzM6f4mUvF6h+C+WZ4PuA12GgwLTKZ5lVYT8a1/zSa9uR86fBLYO
eiigD3JHJ05Klt8heMwRT489n0tCUJIOJSj7QSVxZBWZag9q1iZrN82Bma+crMWhU9jPlz6YN8+F
0jPPMMqVGkggrimsMVga+mqYVp/Eb/PF/LWDZPpb2j5WBlnoa63YH1CzCK7xRv/1HjTl7MszcXxR
iien7dMY8SMXQRn101BrYBxH0YQyw/LwAkKmucsGomFk0OQIPcGBYyI40PKqPz9n44lw0Achz4Au
u26VHClEN+bhIdYEGTgUW66uxlZSSiueTJPih7JMjK7JHBBrVEI8NBtk32N16WnzvdgGwMgIsZHQ
HlrLNGFN6NFq/fMSik4/Bv3zASWB5k9jbW+1lBuonF77WZel4WNad3/ALdaGYRiEbHlagB4d4uvq
syQP71mdn9lN6+3SA7cd8oHIyVQoTlWRCrnR2GdwH1eHVgRszqgzydbVFnQZrXclv6iQOtcvhmS0
HAs43txGyVnMlm5DFFf487ou8B6QvQ1DYFDy5OTI3zwpwNiE+ltnxDiZXMS6S39ucb+uQm7wJUwB
j/NYB0Be5OomYK0jzeNZ4i+7Q8gZWV6TBGrlzgQxjCbEqQ3IlsuoHdlvPQMevSNHCyjN0P1OMp3J
jbGnrQmXhtbzGGNM9qSTpeDPTRt5lGe8fk/CB+RxP2dPFOr5MxsUH7H5720iHUsdpday1aBPcqFJ
DaH8ddipf2HyCLYNsswN1wQIYQ4u44jmhclp42T9MVphe8Em7hTelftkVxuNPNiAX3zYtWJGirqn
FE/OBTsnfFH3sdmpUXR40raOPO/rDcdWP46bUUMZzs7NDvlbS2zPS7QChISzewBVnQ25aKCAUf/Z
nV6QDg+Ze07w+I8/LhZqfhRcqHyGEi8JLFiJ8IB+unI3vGZ7de0HzBTtvsmo9hE/SZYA3Yzrl1Fi
GB/g5iES8XNNF1FcwyIo/PJ1azCewiIPPeNi6R+HP2vNHzz4FabnJ5r0LRMOcCu2LELMzqNqI/bU
8gy4RaHVida5JT6NOtVYgC4s1WlWyR/5TdM++u8WQsiimyaX27AciduPpu5o9JltFCOmW1ylj8CK
JRHH7rNx+EtLh9KTXgivpcptFLbU8MNLunQzUkdTduiciNfNjmuYuOBLOhjerps6NMSO+Wh6J2Y0
LjJAtyCEg/PUDwEKCdQb+XgusOGvB0UcZadXoX0wRm2y5dxwMKtIumVdCDSzEOBcbcbfjuc+RNXK
YQz6DRSKwPwLQsXDO4yHi6IBzCiEJ7D9mF2Uzq1wEmFAaz/pPrqAaRpDDKw6JF+7KGX6w+5lSsZT
bj/EG/24kM91gDPHg+WFraZaf2/ramvwrKJk983vuqR0eQFzeoEWDVK+MQpLU7gWvuBsFnfrrTz2
iKemQi4DFjIqUdpUpdof2vyH1F6J0GOeKyW2Vf0YycxBO1WzVFbLxSJKfioHijQhba3pDuDdXCCa
DqJl4Nbuj1dDsHXoTWdcL0SnjfXttvpYXLO7uu5UvBHEUJTaAYh20YtrHrMYuOvr+yw2HrZ/5iUA
W5dxVnJKpnWaynUrCrEFYRF3SA8tVDKBJ5FsSqziwLdvvI4yRADeYVdvGhflAU9zesRJ/DquNuar
zlHfIHMPpzn29fRBXNzS0DKlkxhKPSGr55FUvlNx2D7Q/+b0TPl8fr3B3fX9QzPh0SV+mpDVyoLw
eQp7Tc27sdo0a43ULWpmQR2Y5jhugE2buE3gX4BdEWE0+5mENBkZzqZSZoCJRRJa8ba9DW+49VE9
em3GP9+cv678kJOmU7RCiXjSboS4+Gw8ATxkcS2NE8BcVEv1HInxr8Hom0R3ETdzvGs2M05aIU8t
g/6SzDzJ4L5h8wrK72iC1geNvKf0myn8Ca9Ua0mQIn/O/ylDdbv6GQsGb1sPKp+2AgGllKqQ9MMG
fk3QCDqxDqi8nt5aERrVIBZQS7VNzFxb6CEdyLj/24RfZyhQ66JGUQ+EWZD75og97wFr+Zkcz3cT
FN219DIiAmbFvGWICgQElAomIrMvVu51sNtsCHIki4bqlKmLPlgdViY4/H2TbdmYeSnEsxbHYYvi
dNOYKUuTgIBICOEpNh0heeHy5prZEKSfKRHE1s4QXvlUs9BqBgIhWpxet33OrbL678ADDCpsJ23m
B1nGBCoc5CAHf/B6I+2qYyzJK8mbMRe414UMV8RPdzyQBFWszLWty2cFERmG9X9paPqA2XFwnoq5
RrjHoRAqficcPBPlSMEoue2bgyBHQT7yrTKQFRBo/yt6PH9tPpzx3CIH/FLwIAXnwo00UHUcLEjt
b0DOrOgb2btTnBbPNdJ2b0LpXCg3V75+q2Wz2JzSCxBRZB2Uw9oU9iXixu/KPF2AtnCcv8nhTzO8
ne9YbTIQRvtxdgJLa1Wgpn1Sw9W89nrWygWcSiS4l5Hh3hCjRJ/RK5B009V/JLdZe81lBv9MSFPQ
4q4eYO1b+HhZWgNDUHpU3JYAv8Uvmsxgj0jPGgEAdXJJT42DbIFh4qY674v4dRjE/yX0AyGXA/pS
+JKViq7Stb7X8X6Uf+D8JjT4IBMYVkPM/pVgHkNABJrDpOxcFwIBQDN1Cn1IPzdQnLvgCuvcCllh
08Wy310xcM1bDRK0t6awcjfc9d5HuHXe5uleid9HU5gl8ZCiygxtXePjf/6MYRjOIm99PB3/Ac8W
NjedUtBRsCF5/58qfq9/gFETeLfPBSUbNgle2BbzhiocL/xaJjKTIKD4Y3DWFmkF8jkM4MIjvJ4e
DZEHJhCRkl1OGtGaVlpVJD5l/XxRkXZt0LHfIMwglweMscYia6rfRU7v8EQU7FpMEVp5WjpLjvvN
uwfq+P/G4ecRBoMlOSS4V0vj7qxsVKyuKE58d8xTHTN5EDORPibZJsoGE44rVRz2ZAh1Ee7S4zvT
I5nzDU4jke+kIKDDZ1SFA1uhVUnhu/xRojCjP8I+CPABmciXncp7uhF8z1PIzvx+IROK3POMBcZn
WuzuTA/P7+dINzVtPl30LrJgpQa5Fc9PUUPSzctj6zNydqcOZnwTDl7H3irzvN0JCcgtghsCO07L
zOYfutAppXF3qyDnBqvwOA85bdjYNfveEZAT6BJLrmTUuTo+EaRVNgsH6LPv7wfUaPMoFVapjxlj
9jNCgmJrm0Jq+v5Cu5pQVpIHK8FgNef8jDmZH2QJP8Qk7waLYS4AmmEnb063fPmJZo8wo3AOoQqb
5l2vemLhUDI8HZA/0kQKj08dObKjlieexcyXuguR4UALiYXRs6hVLVKLxLK9MaZPguj9IKBduOj/
wIMkU7ho9e9I5eyvJfWaRoPKenlq8stp2X2jtAAvAs4tIYmlVOS2uIRLBDkJUueM2CwE57UB4aR5
EHyjH+GCDZpwwwgUlUL+jgKohloO8XvbbBxzeHqME1cWrRca3utWd2y/r22zAxt37vdUQgRVwbbT
RSwgSxM5/NmoaUZnqhMjQBUe7WMuEIuC7F2rSy794SQJspdH7nGjPeehkONUqedBPNE1h1bjwzee
sgC3Inys0mYvA2Dg7gvPKtiNen9F0GxsIgEjG7w6IMKBu6cxGEQw+e8bw1Fk4xatcrHErg+CxNC/
tzbBK1tdPg3+Y0isePEC+RBE9G42VszZvEystfC30wmrvW/M+F7AR5S1XjNdHrGhAIrDcRNnVCUC
EkKW7NITSQ9AdwVSsvpj+NE4/NZWLO8cw0PJDen91s1HH0wT9OKfKd9hrXk26JNgoX6xjLLK40XZ
5QGe0lpsv1yKt41MmOywcmobVlyDL5ceS6Lls+cpmVdED7rPDXcwlbiRu8xmpTQiFcB3838RFgjt
731NnaO0KDNgD/5/R+iSIzIAahEvnScC3OMWpwlua6AuMIQtzhAQW8hs2ATtGKFlfFp287z0R068
JuAJI8sX8FbbTIr5Kx9QhBuM1RkIFwejB09GbOTTwiRxPbXcz8l0T/PIsgXuUd4eVJsxjP5J3ESe
ocXrPTnti/am1ew4lTfeQPGjvZhw/RF0Vdk4FtgPrT/D/j9W4bNtG1CV0VXrVYBEVVpNgNVvkBEI
hgsxsNcko3X1+S8185aVxDl0Q7148TFZumfR6aU3FX79zuxZdbb4J29ArgJbNs1+VY76C/if1mVn
yr7TmqLMVkCpUWbzRMNz4oxVB1OccvA0hoYNUil1zSdx/z0gd/dm81lXhT2yt/FIqpAMzof5Q16B
EKzxOHwIuXWsysfFbUL1DwXHck043cX/fSEzzsiIn2kpGBnq6kKmX5KoAnKX7WPYeXuUetXMVnFp
V71a0YitYuKRmKkVpd+C4lKtIaAgWDi2kH+L0lichsFCCOekvismrX6qcCA0qtD59cwEzn6/JLj8
aVqibr/hY7KdDhqLffnUuEZyN/jN/HwcvPAr9w9i2zLfLBp1zCPNNrNmxEU6zVEe8Fu0UyPwg0HZ
oaZuzVlp6Xy4u63OTHoxoQLWtDtre8cy4KCzh5C5+Gw3/JVN6dbF8T6nNnVGT/Alo5OxCh6YwjPb
EIaFn50nZMQ5470OKFFqjqys+73PiMMvDuQL2u+dzpG6fpWHd/nkvThM+k4ER1yvyHFB4CPlKlbK
a7SnankGRhxkFXjVopG+OtGc1FrJv8QrzcsjPpPGA/wMY2y1q2QqMkqDc8PDnobFNrhfIs1tM37r
cMMMpxp2RCGyoJijyHlUtQHLUwO5v4G6+P86wJSSsn/3PK20Oy9rn8IvuKwPuVYdB6CbDmFD/Bml
A01/nLNBEABrBqEsPBYBARQqSj308fJmrxz0RI+dCc2EaoVII4GYAKmxjayhCVyJi4YVCW/G0Sij
XcCzF2VW1EZ270VGGhSSkTuzRfPfOYITlKo5g+sreRwSojdtFJe2K44Jx86XOpiY+UeaxAgO2XWl
fs8fF6RrvVsivmSA/YihMiHDAcYQpFDbkpxBDd9Xlsk8Saw/LaIefGLkuekDuC73jBOoA7YXjtPC
Liax4UmEejjC1ZmcuE1PunAlfLIrENdrOv9Tc7HINdBzugyf6In1+MzniSvlJ4RGnhWh6DP6jU1Z
gTc/q4ZGHQl8uzAU+Toi+Ula0N4s/rqrLDv9dDMjFuLbon2etE3UDg4n6w+STfvq3Xwqw66lgjxU
mgg3Koxe77BDU0qUwAmGpJFVQDwcR/40F1P2ae1eFVFsO7W1z8gzvjeliU5Mal5CFIcsJGEoWRHZ
9/KOdbT/dZSd9TsuGqCpCSPnTDWNsbY4PNykM7n+HnNlrwk2XfBc5EDYLtvgIPl4dqIZBRru4Y20
OX+05ywuqMA4el7e/qSlHB981FCuNgQ2SB5Wl+ALlShhWWnMQSzWwMi8ttiOGpmqZ1gtTED6T7v2
9+hs+53kCFge4HeF4uTJh7v+cWfMBBV9bDdACwiLcloNw3MVN46PYzQiYMLmPHxos9cBoSs0fV7R
oUmQrC4i1o269RVHVpu57eI4nf525HunJb7GYPv+mFwEJ6LZky3QQGcvViwoamY2PW7djH5laynn
IS0dll5267f+GVqB1eL66HWO3uEOJ4yLoFIF0bUyQy1MhgIW3noEoPAm4OJM1QYFs/NPzQVUPq/c
/mrt/MsvW9B92Y55To1YrCVUBe4uOJWhQYbvAT5fiqxa/IsDBaVckTQl8v/8y5RrnZtuzmJai/2X
3Qm8jinR0vHPu9/m/1r9pDEnab4/NNqIhaClkcqcZQHzyPWfo+9A/dUJqJHMw50zT1PSmTA6JPss
/xl3z6XL2kS/dMNBCPXSrXRKW6fbbpGRNiI2v8c9XUrfUtDWwkkaOW5hCmeUu6VgakvxECRrG4A0
r8qQGCmh3GAcmztLVbPN7uz/H9kQcpLj+dWqOpeV+AKMIKsXP/DLI3p4cxGskqIeHqUu67RYvjq9
SkwipCHA1MuSkSl3O66+hm15wXe9o7bUc0/7S54Gaib99HyWjchjLFPMqyBUM1MGYbDneiwbuqVD
w9JJzVesfTC4FXG79tSNoLJF7tlP3m1rE/R/1Xb5GHErPpMyFq5fV1NzEBVFlRi111Jpv1D2+sGM
YR/WEcVkO0HRlDMf+9I6XLm6rdhpMjjAISGp9P2llFgJRgBgxKKVx/LtLfKxVtpuGF7C4i9lAEU3
4kVYmQ3QKN8+I/jJwLZsHxSGLISsG5BkmdBiTqwzcyCFjsO8HmFHchfjcxekJUOG5SyhvyhBEfKn
QkjZHzlhozk1/c1yuay/4nkDiCBMMRNyOTFGowbIgxrnZvBQTwbdFEobsLJ8JVUBd+DkFonLYJBK
Xh73w5FyYZiBSOHxz4NTy/sydXy4aaUz+nX8N96MCOzzpL0vqknRBQ3Xtu39356whpUR1YYzw72u
TIof8oThpGoRNmGAy+F4Pdo7BmHTlc4N5f3B2vMF27zKY2KrRJorrFxTmhz+9jhNnwmZRlCphhyK
hvd78qLoYXWncPi3mYL9bVclpwOhouY9wdaYycoYApCkh0D3Kh1bC6U+Q2xx4sC455VdsTU9mP7O
n+7SPGsQY/4Zb0fKbGWAQj+FOXLN8jpwDqlgg/6Xj4Cemr3mllHDgJNV1qkufWFt3gO1XSC7ogiu
6HjtH0+ob7UwQp2utzt+Pncti38QwAjUdVf1daIxhxg1u3mBrtwvxS64+Vhe28tMpnvmDNU4NEZP
rcoFtHpeOCjHh7yitRwXEZNwC2LDohZO3ehiLbDRJws99fyNLHdPYCm1/Nk+BpWlV8HvVj4ZmYKX
3otBMWaLn4l9p0iwYOpK8GATBHDyFyeowQJ67Qijiby0G5wpqkBWOaMCpMxQbBibpruC/R6JV999
ClznVAsvqjKkN+PwVMdE6+bKvE3rRnrLGcr8ILUN5xjZ/IH2cXZR+TKaDPWZvNcZOgiIoK0CbCxq
kHBCkwZaCPTAlZkLReLdi9EOQN8rQDjAb8WjTe+8l3hnAwyTqy6pfobDe8tG4/I2NaPycc9Wgu4b
c+wdu24rywEqLDFUgnT0/p6VryuWk8e63WLGVPBLQngHOqNU/4QyCkVh32v9TxLhA2OWHXom468W
8TiilaKQjh66Rm/BkSxwRG8Z5rbZ7rz6esKbrdvvwgNpBhZluijqYPJ3z6eCofCftF2fjAnSSNeD
x5cVgZUzTTecfHsUzOg+UGQ6eUgxJu6gOT9xzlnS/EEFDkcQI+jiuDCXE3KY3LfIZs8bnwrrHuFx
f8mL1r36Y0k3yxB72nrR7jIPtSqpFQSEKsJO88rIN53cH898t7+d4sqb4RrxpCkNFh5IpiYY1pi6
ZIBBolDz8WD/AN+fhfvKq9hNzK/dZ7ie5sQ9C7h4ZiEv95Y9HWeVG8VF81ktERXSP1vUuVJWLaik
ueAt9CJ0dWN3embS9nSBLo88z08zC72AwepTph36j1tDBA4Jzf9s9mfOwlz640squzDposb3IKVW
trgufPFCaSRs9WZf7IGW4xh3BQ+9YDo+6rB+KAAWBWLAA74BZWVP4TBiod/TV4LRg1AjWQMjl26G
tB9dDcHwDP9Gbykg9+9K119vfoK+wLr3E73QJO/s1eEdcHzwbWJZYAUPAo+sZr5Qc3fs8Y3ICMWK
2CNLcFNgEQx/yEUBgbbQlJSZtBAaUVFZhQdUpWjdduycJMa5fnefoy6H/kjPc3ATwLXMEBmpAnPs
BFJy9dBUGBi3X5Nqjt7/kdeRG2mvFKGt5BuWQ4IVH4Hi66bZnikp4UGu4EISLtzXOiiJCHvlde1x
5TWHWeJAhnyjdklz+xlrTfRtqm90qd8j0GVVPKDYRbqE0TTbUxRebajK+4MPs1ilBww2D3dr1GrK
rTOHot3eFL+/i8MYJbTQOegWnNhRPqMoWHsS0mnJR7H36O6zSJ5qkXzz9nMyG26besh2/HDIJt5C
VOWvhlbF4Ar04MUHZUdEEpBoPOcgfekYuKX6Z0Jecn1cNzdX30eI9oJO2q5kqz9SnEnA9rfc9+wx
QyOJ1ArRBf8JzIt1TADXJfNDWEnbiITRwMXHakFPPezjRLIjHuT5iuL5voQ98xpXSBfXroiabNkX
7dIRFZrHL7VZsBEI8tsxV9aFXzGFhagBVQ+tOMBaZbL7tptzZiD/M34sNETUUF+f3DJQ7rOQm5Lr
7j4xqJlYs2mJ+dVniSsNazLsDBnrmNV+D752XrwdRDycHUmJsSXF2/J275nUrVmFXRNn+Tv2PTI+
BY+P9LrUKBxtE+vzwwmBr3isQiWM9Ai35LcATIH1MZFRjZGw6gJBo5wgOsMqkniuWV9O3UJS5b+1
ZVmp+qSXhrjcvQQMZrGQ69sD58OcYD/+nUOcp5bwtkIYS5QLXq7AlmTAc6P5v5PNDewEGmIHRMjI
QNaKLn73qJVcqhNVE+zKW9akTINayA2SJIxec2d7Xn3sRhx0qHE3FB6ah0KvJrDON48kOIUB756j
8Om9/d2p1ISzAg18ol4rfWnNamYHXqZrXyd4ve2f0crq4OpOFHwx81x3mF+KGpz7HHE9Aq+jlXGk
xJRruNGTcOBbqnRkOzDZd8ocDTzqLntZ4FDA6BELnixTwG4pExEZrT4WUFQdGdMdBbxp1BoU8rt+
Eau0Hnao/sLF39m6I6pu0Kp2i/HCnjcr79cXLfROzjjs/ddm90//woGmAcQOHcBl7zwbhDo7BEvZ
ug5LZZPcfJ83H9DMOCvgUbF1zIMGwYUov2H8XvF/kMLZVpwsac5utkM14COPT3Bm//bhVW8SmK8Z
e/8Y1rB7lOtKV35K02LXFLt9u5NupLVrHtRXP+pmvubJ+rxini+d2tHffui/Hxpsa40PKvwKNZhu
Zd0HqtkwIuZX53fpI+aLmuuheP4PhkTy6G/Q5jm7Sm3xnI5j1WtTFgScSykyhk+j4RQYyoqiwxg5
TTeNzWdkGUe9jjgGmVEJUPZdGM81bK54uqW3g5W01axF2Zw6vecdbtpuWd/gXjXErSSY2qyGk8lA
DhuvVgGotZpOgQhiVMk1ici8OtXuQADCysuQhhVfhlSJPSpzGiy05KitzYynmE42c4oO8mB48xu/
NCcOjG0iyvYMkH+Yf8KZrAJzVCFiId0xwis7T4BuN3ESkVBlsfxhgFSE+6JFYDWKZy+eiXGlLxqR
nibQ5uBeHgAQR/k8EvjQo5lKjVTh/3y+dHbVBYME/LXxIC+8ffIfsVhyzSIT9bdAsmM9rcBeEH7g
QgFj82ZyI56rD/wSXnfc+9xn4EZuM5ZCaefJtEE6hUTsgqfANxqGRK4KpjZMixN8pRVbFLxW6U7+
8WSG4yTDiIg3Af21x42ivi3j41cRET4FfCXttcEpiI2xDB1nW08iq6ZvAWBBdUWhUgrdxPYKTTso
we7eyK3MdosBI0BlsmGNIYw6B+6NhEJAZEiJTmb8raESRyR8tsh84C3PvJL9VebDAmtSd3tQj2wI
gtpIxE0thyYVs4ZABsU2sKSPhoHCil9FBOk+t9xIKY1hQEIIjfPuhBPrHWdEf4BCXXD+VSUYjYPn
8O8VCWSGb8fnEatvi6n7C1Z54bxEe2HCAQEhfmiYmm4b8FSjmgkG4pCffOjuynjpXCPUweQcQOed
DGKGEeOen5WWRZwyx/Omj/kkpr0znlMRREbJWw6nM4fUEBJbqXa5AmxGd9myJrMj483nYaQZNaxd
xwyvhj5lW8pY+cSPgCG6rFCOxi9O7CeJiIs7HlQShCROSeGyqRzD2lnw/Gqh29HG9DId+SfCvxHn
qDkPe6ISfsNw9J+zuwul1Hn2K+y5tpomcH8yWo8DF8HKaKX1mDynpFoEiCvmWyfM8QpLRI4JU2NB
Us/Oriq2lnhfgh+9UtytCmUOs0kvDphEFd2lyMRQYQC7u2igZEShyvC0V9tjaHYtCDcuHCTAY+bO
FK5hgSgFU54mH4yitWQKbiGIFKTeZ5h1e1LvF0VJTDJ6ppQxaVX+/lpZrRveArtQcyjNfUAqZYNJ
x6jFKP1uEas03yK4M8s1k6qpeXs2upg/CufpnKEDwFgJGqLu5+Cz6nl98EvLG6CIv0B9yIwGwlOh
oGWTIPL0rR7s2RYbUTe0ZglRyiELFRBj5htezeNlqNSC9W3KynXbY9OPN8Mo2v+L433jM92KQrHQ
0j/yfnEPy8BZIEvR+6FqK9PBnhMD71uNR82eyWgpVpFQ8TuBxaeV2FsNcrg36+mH3dZ5hLq3ASu3
fqlVws1y9Hnu2q/n/DIXZdGcIsNre8I947HkiedEAf5o8XvdCa8cHH7//a7iFCl2SVVGc5ca30m2
6ly6Pk3S86DOSkHyUUbGM4loamVC8TzQqL8SKEtTJvvSZhvTPtr4qA3CnnFEwHlTNermVTCnMwso
r3ErKyJHheRnBxzAOGW+kyHTiwX48hY1l/IJvsF2XB/IB8otdQJtW3wYNaWfd1urMuRCgr+8VxDy
107zKVPnzflB5C02V1OVj19EWGwr3XLfgVX0ofp/v/8FYsQR09X+wAMMkLaspQ3Xc5vHXURMf+iV
9pHSNNyVzH8phjE1VQ4nxhU/oX2LKCf4xBJWwasbquBc9XZRGSUHWnDuN8a3g4eqFUDGYEuIjVcA
J8cNSN2hkQQUtHvZXqbSmvI3ga3Ns8GeCbr9jaadqmEUPARcvfhTatOomMTAPHMlLEUXBYHigqwP
lZ0HRJ8SrI7yCajwiNBylNMuvXexyI+sxkqaZkexJrfBo2gfrTNQoBONjZ97Wp5rZWPf5QAmX2J0
eM8bk3tL/x6r57oewGqCSfy8UubT8X9MgxlkHmwk6zv3iJUSkcN/CHZ1gsYb0E09f8JLYl7AZnmQ
LhacNRuEZoojY0/ux4DXigiPLX+ogiOiZ612j1vbTaD3aAWHgGTqMeUvI5o+5PaMBzI3C63osvI1
dM/4gKyQC4L8PTkAPnecv6jVhHOPmKHgzzF3q0WwFlcibaVwNyp/+osm3ZjccgK88oGF+rc6mZk5
dPnkHioHY/hKjPB/P8rpr/Wp5AseeaIpTqj4SeTj3KBQmd7wStms40QQNlPQXzqMbN2u+N3uC8iZ
1LSjASWTrHQoF36FPichHZ5X/BofjKKnhNAS1NSJ1WHAq7g8a2JyY/Ym8icGssDc1IEWXFhEajug
xJnqa+CMUBkUbU29j0j5ozEs8ktQw98WFekMDA8tX0PvZ4wbJzaAidonM9oz2Xlr/WEahD2n4p9S
pJWl0XMaZM7XrkKTYFxspVGIOoLITHTkNnuQPegYe0K05771zIW+EL9Koq2yveaTI9yapRKD1V5h
TCZfMJA5RmQ5HHZ5XylfiOGujFSPJs6T1yDVitb6FrLCoyqi8a4ezwoA13FrW6xOv83Msz2YraYx
BngMJp19vWDX8gP2lLOoFPkVDwiELWJSM1wplFpaRXzZ06+8W7PKSWUAcgAmBBWhgIVZaepM8fhF
P/Dv5hzWv/QAI5cbDbVscR9kO9K6TQTmgLKRC7QbSGMlS8fIZXbTbtI3vdBzzp4Gcv7c2tO7+w44
FjW6xL4X5ChT53aeckxB7U0AK9S+MjX7fZld47r8Xo8oFBKYohozz+cWpaKBpJyUJ/uM5J+zv/xm
oO837B2SrAikEDT80ZLnkVnJFBPIsA+G1fySeriMTaGj3WKvcpxgCQ1Z3NrlMREbG4NH9RI1PT30
0OyNYDNq107TqTPwb5eVpjeTNuhKnYn33MPDGx+sR0ZonKJ5687dFt8SIE+45kWVOUEp54vgFPnX
zEgWO2jAHybEN6QKUqRhq5+b+Cq6LE4AK7/JbQ7i5g7T9il59sgEY+HHA4OHWgikN+41lUY2YJ4M
nv4StGniyupPf32R30VCVyjQlpsA+kRLfW34+TkM8yYU9nXsmHPf10WirV+r1XiwCbGaR2izIHmj
cEKDLf9Sxto2ZP2V9qCyUmENczNOhM5ovPOH+R2sAST+v1RIjAvE4rgZKcsMon6/VOjWlUOe6ZUp
+hihHEAmD14I8ECMyIDus+MMpCuxrSrLqPokv1wPWSZ2SzMuyyPmfXpNzOptVH3bP4m/K8EWymt3
3RWMM2/sseGyl3G3XtNknrrVNnvOraoHe0ayAhOMb+HVvYSpPskFnOt9XKSYpevvC5wdG0PUAbpU
X00Ryny9iIPA5DyvvhWfxFnfqSeP+igTbQSFADqCtFCioGO2OrV9q576s99Qnq3EpUyouvzqS+Us
B/eFl991HddjjVLyUOHe6ggvT4PTjWiScfX9EdhRvOGaw8C2Osupo0Ijp3BlfvzyyoAZEur22g65
X7b+ttv+yrFJdBMGat5++AAIDP8OOkKFmQNKKyf8CcxNUDKtPF8RwdyfviipTST/HLvOxcPncYvq
z514p+7pewoopw6RqOUDfbry2EzUdIWY6V/oVvfbT6p/VV75MCx2CXl9wtGM/kOZ5H7AXxonQbxK
hHus6+llUcSmss21McHMCBXKh9D4RNUsM8UiBzSWlWe95VzU8qHAwqsfp8gD0Xv1MwJOqORu17Gs
tSDMAelFClO4J9LcI9pT1ONgkXR7c0HncTpPZRcVeMfQuyldg7c+k4lFLujLvP88xP+sELt/gYXy
qBVFd23OKPtPFYan582x/6AVips82CaeifXvx4efIHxpaVLXVVmuAwoBm2s5XCZ4CdAEdtNUT30N
DOL50LmtfyFKL0tjx0WZlk5AJu+l5pBOQJs5GcBnYR1htcKk7q4rMzEylDrP30W42LvjuRGBSDyE
X4azQnHRa1kAo9MMwikSTNozLZ6WmXZwV0aQMUp7jNwMi+4hheYkHPgIbrCd5HeHy0vIYf7E7R6/
1SIE4tHg77gyh83CzRc3kZ1gpsO2gHhTM1EmHGcBHjpLLTWuOmNIzKNGAJTKavFIWBATe2c3aMH0
9t9em7/9Oj2WVEYSpkAZAqeUVo1ombcGJ2i9wnLwefKwgwIGPeRi5F1/VMxSlvjE9s2vQN1/ThzG
Q4AZtjvY6oiBNYZfAp0PWsOk+kwC2vjoQvqdCSE4zbdqMRMH2/ARbys+QVDjoSqnlMlnhwXgR9rL
DypbRxBEqggHLgl/Sf5cPRBDR0lqatGKnzMlVdTmvo9QrBCMV4S3uNy0D1zE4xK/1HAfx6AXvzJ/
5hszmgAoDjGn8atx2QR9ZPr5MRa9YIqh3DndNfpLMB8/QOBs0NAf7upX0kIWpB1u3mgxFXi98Nir
bnnod1/P2eTDtfuoQ7we+isArdorUrffG+E+RgBNWcD4gg2378/MpPqMTq6a3/EP6zY4r/zpqiyc
FF/2lbitUV4+3sDuWwkOyGv5UL7L3wF42/jyWZ3eQENWNZyqnuiT0jjiR2gy7inPAUE9fWGadjnd
oIzozq2tIiwQrHvVvYpQBm/NDkCluSPZnNiMyz6eMu7E0eMNxm8aAj9OPTX+cPSwBTsfAkaR+WXw
fKs+s66H9nlhxreR5ZVmLsn64OqSwPbkQzko5ytrmqAx7NY8fxuTZpKHE075sWP0UBPE9RgRc0X+
nPPJtQB2um9GLz27uYAV9tqqA/zTiv+u2HJetIuPqXCh5AY7+9rWwcCSN0JcJn2wbvHcsusApag+
Tn35/BQoX9gmjmPxxYRMAFNN5a4lI2N/Y5t6YFgw/QOdtP1cd3+mHCjCcnaVEA7PxJOOzDxjQfFZ
/0oD59JUw50ySWnCI/CWbkdAK2pxmwtSr1X1weMJE5OwhzrI9rDCD7pxkXpzd2feRmL28tFFFGla
Y3ZZl3A4n8DeP10kgWihRp1g4CT+bw1R0FEyLy8imVcEqWZ7GqbSp+tGjIcSsV8syVctCraWa8MO
GzwZVLm4PzaH6Z/fMe5IB31gldIu9LVbpnrCQSxc2N/9TJcfUwAh1in3HaN1K4xisiwLEylc2i5F
i9OkcD/8Cf+1zNWw9l53IoYy6uv2ur4LooMg20R7khID+zYwnuvEqmJkDTDadoYf1xoSbnWEjvfY
RGkzY1CDCy5HXJVTbakxWBMMbndoJw8bkaiiIH9jdVUGF9uKNRw7KHbEYI3G789EJPYS6oquDVDn
0/PNYGAqZFKUXtQeSUm90mOrKzN3zUTTGIi3A3Y1K/pJtdF5bTn7tmRJroFGbLpR6vaFBP+P2f8V
5fPF0+FgB/jRH3VZiMW9B02PR73GRUMdn5ENWIlkHcZss55pDo7dUO56KJiW77ioi71IgHN0gShh
xF/bJI8wqVWMDoL2+2UzSZvU7XFVabKRELMqQLpqgqAfctrfs5goOhQti3/wxHDgNsUuig89DOPF
U/PTXfmEZmhB5oGN6ejBY/1QOcsJfkzH3l9iHB9QdGU2+Y1A84XHUK5ppLRljF6t+BXeKT/y0kTG
E4+NWkkFo/TOTngOfruPV48eVGxVgfMthjsat1z2a+AUzHzWYKwgHlfTZrBs5jH7XE0kkLEQcJ/Y
t4H42n/YCHjleRxVAOVLS7fY0r8iXsMnC6fMmo49eQWM7X5wwG+1CsafWpu+p+476rrwmi2ji2el
qdt7yG3gvv8w/XMbDVvzGoteFNDmfUWkhBRlbaKeGV58ySwrwY0mQO6xUhDUyayR0PieOmGI68S1
DvyGsPdLozX/eg68uBOMIEnDUQgc+wVjix+6eArq/At8CBgt3llZy1pjus0209SK3MXgCl4kFGux
3HOQAfUMo74ntKTQdLpXqppnZjLM1On3VmaErYgbVX9N7Oo5mPQo7uvi0EPQFTir4gBJugMoxUgu
EiT42mCbyU0bLU1yalTvhCCQKFy5vCVPBFkGo9exQ5IZJv1JkAhaPcY/PSzj4AKdeFMQ3OGkXw8h
6qms8Ja7goaNHIf+McJabJZBMugPqtKWHphT+0yw1L4Xy3tnJOIstg4rE72hqub41zCQuBY2VVzK
EWGSnaO5Sfytk3MlP5nEO+JGHDxUcgcwWW1OgpG0snazhN+I1xYIC/LeqIR7fNHhJ89IS6dGS9kj
f7u0eoA7XOesGesPddczpzPqlYLDy1jM3DNwXL8yTcTMnMdB+Tv3hukSgJ6xsh2ocl412rshu+L/
ArtuKFBY/iuzXlpmtA2UQ8KUtwC9E74DcCa5n4tKhpqKYjWJeg/jAVpEoOoX6SRCQPYNHAcqvBwa
9Wameb9Da8zRKQvXblf+x/4O0by5PVSl+G/OU/lJQxTxJrEP+xffG1SJszFaLZqD03ONDS4kbR8R
AUTMmwDBPS6KCsWcFt+WOy8Il7C0cqHhpZqc8VKPdDqDP2VYuwk0cxDBVTbw+PKNMa5Yx20bax+4
ef+vBOfj4omgXcqteQYjU+TT0CZJ6ot7SpOEKySE9LxC61Pf6pthtB1lmCa6tISrWB43+Sy2R42P
IFyfr/qYYt/5znfLS6mN2uPKePjiTZilG7FBYQsaE9nxEM3P1k0/XPvkj4LRQDFnRyqLRpibuonz
26Oh9nnqKOGGAhcKZA2jFbKYCB/4lT1zDQRzp7TbYVYspNN8Br2zt5AhW/1USKeya1NnTrWjw+uX
vhejQ+XJrckBV3Xm5HPUFvwBwJhAYQJupLwiN4v+FzhVjneJ9PHeIw+JijUeUrhtuZi7Ohni/I5r
OsISEjKfO88ILoKvUtUXG3baHh4fT/806cyikqvwzTUPMilUMQIAIofWpYsQT8pdDjS83HlLHHiT
DQRwRaja7oPdJbnL/4IibqKu44sqMoNX/+LjloFjFlh0GYb130h4cLI7GWCxl0Km42zPpljO5aib
WgSoIcYyS9GK/L+2tqdwGLgwyKaHizWmmcMr7BVmtVTTjBw0ycE84iPHj+WD4tWp85gmthR0LPXw
9BoPlVN3jsqkx1fT0wsAncPGy2vWIKiL4ggAfX34wOlF2+slwXwxugkq7N00mZ+qTkuKYfHzvc2g
E6sxTu8cPda1VBxKaQvm8nhRpHv1T0ortucp4lCfnToMfw5lDojd49tZf+VdnmY3egtOyFv7JSwJ
SiuhZ8Aibv3Lkzoe0/RGZwYH6cxDyW61wbZNK6xWy/+K1KuGeJmeUJ3sg0tHZNdhoL5VhIAe8d65
AKc501hbYcmenNg36hzMj5H1xCtizZ0a+BexjeuYVWbWzzsFLkpU3ppYW+jtVtav+fxZyeKwP+cR
QaBHDeXg8rbPELWQZce7Pt5AfJtHnrAfO86UcZgBFutRprAtINFPR131fBXbe7fKIBuDH7qfKnsE
sw5jNRKo2cuJ1ZCveW82LAI1dBC6+fjmgBqJpOqpaZCAtT0k76AG0CupePXCPpJ+nxloU2RpQrFj
NmFFzjgf+r77cMkFZlG7ygxNEQX56srG+jstmXG3ZGDm9XBjCoCsOaar00YuZhWiXI1VoWHedhof
IWae6qooUzbIkuXbEhE9dUPgqKYdD166uLwF09loiJ2tt2URUs8qm33gLunEsdGfp8uKiON5VGG9
paTtG+PAXHlteZ0eRFV5SHcoNzjI0jwgCa5N87Nu0Reej2reoLH+RQJj5ejJVSqqg0krDTwyI/Iq
oJZgY3tJO2ReP7HVNhRcyplVIorRBGpP1p1cjZTZ7IbaUt7CuzqusdLuatQO6d7GoZybqUvd3TwX
ehZRaAkxB3EoSJS4KyMpRHxir3n7/DkEPIsA3hLphxqjrSx26ifeQV3F5YDP+orY/zNn8iCvzeuu
KW/Q9+kaMiegNMU4/fDU2YDbaQ07LBVC3R9U1XC/iOX6H5FFKWCiZTFRpN3d/DgXlE7Nm9aVOGPr
N2nQRyS0oKjEwtM+fPeho7/80ZkkQN13r7mkFDLkXav/OBtlsdvuQOoDBDU1ig8cv6YiX7CYdYfA
3Dbz8QCwy2wFWO14B48kAe4z7oPBJjtQMwDueM0+a0lhLPm0fXBJdhZX/5E21Ezzpx9r23q290v/
V2P20EqPTFKXGX1eWLieK1Vr1I9uguMpHOB6L5m0R5pN4FZvVlS6qg7LNdnNImN7IGpOW9XA+bv2
E7HxviKEFPDjNxYj9zmenrWmMjq9a06VNHkRaIHgVdvNNZEQEVhJKcSRqGfvPcs+Mkl7/kXaJ0sL
Mcsi2h7pDxmRRCS3dPIQzqVxRxr9W46tBRPaeS4j043ymCWMrUDbjLAumJiWUo9xNebovLJ6L223
JHCAzD3eOx/ZHGPD1NOs2uUoQXJqmVBGBMZcKEAsR3BuzjNIQt+W5m8fi29s0t+KWDmeZj4lp3JX
LzYDIRbYZJ9BA2fifzaKLrC+Vcu3iN1OP0XzDs1elrgciofEjav/g1OtWqassBKTuJdwsrkT3dT4
sepsqcvj8N1yAHB6jqXsYUnL2gqOYqZ/a4AIcWflLiKvXSXuPFmnfMWTl5HjI+GrBTePXgTFFt/5
0lePimN3bcVc7vWF4U93GdK3IRtM2XCdUHksIinGCALWANQImE0LaT3Cz+CNzjXVObfwIHp13CiS
1k+lxsoefTo3a6fkNpLdDNvzuV3zr1PrUZ3NhkYY+eAKBMChoWY+LN8UEfFI/eH6O52e1HO3HbPk
PhizYfA/yyUB1dFzPvJDLEz3SjFNLhpbPmf5MBs0OxaGBdjKcVnLteVLuXoYnSSVGjxqEF5+9ejB
zg1b/Uf9uJhffwyZpTEigW3TImOZRAvSKwrw0W5QbZkAr75ASF06g0Anl19x//8bVSsMf5DKo15p
EKb7AnNfrvXDXEj5C32WBHuzAZZY5FfU13SDXPYJbtexGGI/+HJz2SNWujk6mCo6i7SF6TM8oXf8
8Y+3q09EJZLRKb+pHXoz9QQncXXktNo8vu6NoCCkeivraBu6/k6pw6p7o0T7NSf/WzR+Ycdwct0y
NaKwP53+ivZ2AvV971VDCxovWppJaGOu88bqwH0z7hGRu43bcrCaDZa+MtRdZuENcP6s704PswPx
KB2HsLNgYU3D/3cRagcPPJobSKB5fXnfFiDfGwO09267byfubbb7Hzjf8aXYe5QYrgvE8hCcBQAW
2kUz4ykCRMZgz+lqgaPH2NUNRmTxbPuX/vetXlKsnAMRg4aem/IoWNMTQMU/+gbBTs+je3YPY+EX
dBgogIztL1EG8OZxceC+62ZV1RU4czFOt9hRlxhyBL+Ck949By1mWfbb4K7wyPswELAHaXrkkmhD
6qPtDWgULUP83inTCwg6QpfGdSij6yxUfMm59Cc6GiP+D4+knB+aeIrGzVivbA9v7Xt3I6ghe2Mh
LyZiu42r5bbNDlqlx07ZNOrofFPOeLJ13YOFwlFHx5IwpaXoeIoN2n3TPE9koS4o1EQqaKVyzdSU
Desyfer+QzQ04EzGBtWqU4QGzq4JsZrdRJl6lbZGzRV1Y7VpYyWtxXXIfvK2AOL3lQrwXV8Q7a/h
qlPtZwLSuE8TCNy8eaavqhN9IrutSSU73iyqT/uV2F+YUiVRHw7p6t39oskKnvM96aSire0AvO0t
6ljfllcsBh5iXUxxZs5J0S1fTBdyAVazEQl4sf6RaCPyrAJ/WXz6CPFxmjVoR9sifljOUKC9XmTJ
vfy5gTpjngqaDtQ/aqGUCvZD43uHrX4P6tQrzQbQLI0OmEVokdOW2MscYadHgQ5Ok3yCgF2W0Umo
l7zPlL70HgzhIWGKMHJca75itzdDGlSca4TPrO/c/9Vl4w0DgzZeOPaEF3ioKgL78WrKZzqLp832
TC2F9FZOhpCx8A1Y+CjVPTJKz1WhnhJAkcb9cGiu+48nAH+tOfv5BdX2VxLnCB94Z0CvRj9X+i0I
b4RXVjJUSH4Cp5OsoghGozJKYytOCX8ymFZ1Co/zM9Yh55kDe+Iy4zEfNDHvAboRcrGzJ6zS3UT/
PH/ee1xH9uBicKvRvSUL3fuiKFYvK7WiuRqzlkPuELXLJ7Hg6ThiTM61lpncLy6IEffzj0mMUJ9M
O7N9gWYOcLSJotHPL380DdSPgGfdTsoH6S03vXa6Vr/LGX8PVsUSVCGpfA2MW4OWus5Kjj6wWCyF
XQ6x2bf4JFKojojb6UU6L1P2tTjdkSlLvtAuzWuai5NrdlrDMEEL5UGEQQe7VUKyNmosWLn0rBVe
mWhZTgUL2REXnjIz93fhumxSPQoViimaLAYQEvZH0VX38kA0/NTXvbl0D8jXbH9JIKhjLYA55hAD
vwac2pX0Gogf/8uODkcfK9I72ecjM3v/3/O8l1h7VNhVtENsDyPYtYNLRar4tQ+Y3hcGbYEC4not
WYYc6xnZ1uTVHrQzFmWULsJoxN3VOoVZoRR2QKpPlx9aYJ16hqRD9ms/Kn4qC5ByW9LOM69P5dO6
MT9QinzHpg2083bb3sT9SxHWde9fc+L+W0fr+seHYpyOSwhi+tgGEezWMrcMrag3ODuXhmF3e4wS
44I4HNiGetCZ2d0SHJ2ovazgQBI4itKv6dwI3IEMYq9ti7LjxjvLcJOyPc47tEZJzEjtw+xibAOA
yqar8t6dXMWLjK1VJ5zx/6gso7wYNYWGUE/svdokReDI9LHQqg32TeH+sZhKNfofKcVgt+GXKc7Q
qBGPRGFYOoS3vjXjBKHsOSgiYq+aDgZ6py5gyoCmprqD1pAHc1r8sddaAWtbn8spjpv6haN/HoFK
y245SMo4vR+ZTFzOW0OPZxEOdMIwPsHBeRuLrPbVwXREXnRFHfZ3a6dACsgXGaAcyovIrPDvYkck
fNqQSaf7mrHNtDh64ZcAttmo6wCLDlpvC0y+j1Rh2EcrLhJl8MsIXUH68SiEf+BEMmZeaiFZU/mK
a+Q5NU9tMjiSLoe6CiBNIkUJVzAdOXNc8MWSE+QmeNQSEE/9rmBN85cmwNQ3RBpF1oIfu9AitaI4
ZuZH5OEL+3LYWWtw0Nd1mGL9japRk0NnaJlmmdir7N+mVi2rRyoYIi9EMr0xMLjLgUzFkViqE95D
LcZa76RUGE9MOrOTAqHlt1nNj20Tkew8Th6bMztM8FGDRbXdKIkZBQ+X4g1Nyq68D2TfMIK8JOLx
5yErxzS1tDgT/hs7wCoxedxaq1zO0B2WpR/i1pGgSdqSxI3eA0gfcBm1IBUQryeqR00azAfntO7K
G/0Ql9KbahYES2Vb3Tvuo/kqKHA+yMQPz4h0Aey200fMlhEEXQZ4aMcyXwcAcFbtiTDuFxAbb8Q/
l/0g76ZSon7kTSX1dyl2aVC84QOC28OpkcpW7kGT3hX0ZMn6N99QZqsPTafohA3g9yjijlwIYzpL
iG2nEwvZJ+FXMrUqWPs7AVDkUhzzQz0iR/gU0iQ84/wgOijTdVSFYz019amNV1EImTCSSuVBJV22
a78/BOaijAlYGZR7ID4B96TyvtM/OyuZ3eYHSDS1/f2qJX3zGDx9mlXoFj3BuJZDanzlckgQeMqD
mqBs98kR0N7S0dj1j3pQxbcRhtDx6yOvu4R5e0D4rZUdeuQRLNmJtSOumJLBUd15mrZP25mvC+z1
mFyLE7jQYCl5HH7f5RSJkUgDoX7BLboozniFsDnr8Eq9LpWtPOytYFGAJipRSCLhyqivIzwE9wnG
hnWR5/RBwEnAPvcgcnZf09syzip2YMBgghh9aGPJiUGRXp9LWWJjymhUyUwHoM7oPB2M2xOKlOOg
7U+EAvGOs+WR3L8AlJufFWDk+h/z1wUst/mztVjyWdOytWFdDO/nHracMEaqjpdzyiyZVR09st8o
lrZwmu2w13XqvGSNo7jfcS6ABNjVHDu+4F+MxqhecEC6ZEtIfxvqjgwSfft/rXr13lUVOfMuG4gC
pX/nPWIxsEBlID7NGL4lq9/XdriFI4oMDwmw8KvNHDCVI+xoX8cr21/Wv/urUS2rA91wipafd3WL
WrkbNKdO6EFyUkOk7BVYIBm13AsHTGppM4pLYL3Hjbv6+rPIdr8mmHK6hn9Y7mVWoh1h5I0JiAP8
LrhgSjizYg9cLFENeSQqq5Qi76GxKe3gOL/96T70MKfHFvTn6i+CIkfkQxLX2aprJlfFv1CLKRlh
AYP7rRqwWtT7Rq7tN+SNdE9/VaIP+XQTZycTt6q2y5d4h/DE9FQFnbayyFkKmgpm3hflKv2mHHeF
+QhMPluUDdb98t3u4z5/sKRiei+M+f31xWlDtcpB8wPpjd2Dt0Avw5mCufhJm6gEAX9zKtbxIQk8
7BY7t1CmHUCtVQSs7GqzNwKaWRcEqGm1GetQTCLseZ1JH9GsTUlz2Ok55uhAgQwg+hFo4aXzARpj
a6IftLS07HU03dvOK8U8UwsnWtJUdUX52sVCAVjq7GHXCicpuXPxvE7Ems3el9IbbW4aWp5g8E6J
yMVUTcEMzyAbX/B0Wr95/7m1sLPTzOLvdDxWbxlPXK5jsAYgk8EuvC1UUCcsFbRQVLz9/TK+t7Qn
9rOeupioTkLyuOiPinoNbTsT+MxGqUBt7DbVi1l+mAFuhLAAt67x6xuDqszzygrP5q/WIzqFIpV5
QiGd3T6VRibHPiVH1wayPKaQn5g/sElsjVyWmjhxrjix20+1HArDAq2Ms7YJAOLC+fsqTQthjozH
TDBJh4v5x5/d1t9YLN6Rca0cLXp2EUvhDAylp+Z4SZodEawJ7dOlPTVU2mgiwC5SyonspIinQy9X
RvhTUa4BXqWkvlXuxnptjo7ZahYWYSNnf0Sub7RfPLzNmaC3D054O64wtSp1Yw8vMfSSPvPwpOuR
uy+OXK1rg7Xnms9smpjb1Lw98YG3oO6GWAgvTeXnRKzrNZ4Bax1oaV2LypcpKG5w2ngNlArbLB9q
SmZ7A03N/de3EDtqbq+qOVzRLx7BWFQLKuV3esqU0ciW27fEi5NLfK4srBTpiava3hUorYvwKUyG
ZYMjEn2e7BDI8bO99NC7GakVb6RcMRH0WSzZwFY+MTXGl+ihOljKeTV0bgk/yio4g7zgaCn7N2sc
mr+i3HWxPSLq+/+DrMPc6Zis3EDMP1mv+LOKMbGtUVPyZMO9nimAQI446cggLytLsjYDhBHiuCEw
0Ntuo3ZE2VgYAIFznAWsfDrXmQ+lKfioz0dSZprV//sYNnmQkV0AEeCFHs6c0ohpqhhcBtYIjaKp
BvLvZ5lQpOYJihsCGFzk6raNvww4elwBbSP/Wob7ftPYiDZWXQ3oU1XVQZ6qD8PkPm2xLlIq2qHZ
aIAZwHP5KezYB/pScwr0yAmaWDLGbm8XNk/7DZo9W5dHPKz3Z87PYoLfi+rYKhRCqWurZ3svSp3V
URJxByjQob2SnH1A1NQfSKRFqhzqgE50CYzPcwuoINFIxSQzraGrd25P3020zj37q8lM3sPphCzs
Krk9aIJxBaZyIDo8OYC9wo2td19CAK72AAlfM/Hc+ck9Aw264fOmR4T3N8idRt33QnT5sg4sjO/C
pUqEIHketF9GfRn2x7v8JQEBh53F62Du5yMFiVWGQaMOaedQiDodx5aBsw1snAL5IUm0QO0Clwoh
TiHNJpA9M2+LGp4wKdkWhMy1frc2cmjEgJa0EJbgzm5JDvSPP4IrXuyjQByMkr9VFoEaEl+BxGeG
27kjT/ne01fHJUBBDpfzh5fy+y5hBuEckMYWZNfSu2UJ3KTI2z0po8f7uadi6XuTgHLiJLjHFQEU
HTanZip2y0cn4qxLbkQAIoYDlb2fcmU5+Ky0sb+0U0i9QBDbo41zptJ4yMPs8zxYnqc6ee34kkhg
Mi9Q3okGgyAd1S1St/oqNqnaQnzNkqGhK8Lvo/dLYTNSqOU23C5uTKQkycG3y+4ZASh1hxvOSAIE
iDEA6v+nwSoVF4mcqBfFebgszT6iYe4KI9CxBBDOIRrwMWzQ/O0lfQB1jkv4XQkWUcdpuyGeSjhQ
5Rl+MvdLetXd0nCByenRlQCJ0LGum1TjXtmKMiUQzHyDZo7boL/XqRJ6CzHgOyO4R3bBKgomPT8c
pZSyCodvnWqqYl1EtpA22KW9G38W67G/GnOt6/6JF0t9sguOfZo/WsN+MZNdVnFh2x7P3wgC0caq
cz8K7Se4rq6W5NI3EXnIRxySzQWPgn0OGrb1YA/YiHI+n52rmS3NwG8YmMCDTSP0pMp3iQtGRlcE
srqVUJHy+12WqTQgoBfd6tl0bbvEKR35wYlLZ/dj5xgyT8tJPWDZLo/y8neSl+DBRt5VSChh0v4e
SSS7lKBoAwuxGh9evz52wc1AREawnNrGqEOrLhpqBQku6JEeVBTuGEKcOy5uNsOnNmx2rIgrEvzX
xWorgYGQp5+ylVklHAxLmRGd2lskzNoZbi8kz4sqG5bOqB4EbnP4rZAjQ2ICbhu5EEf3nnoZFQ//
/jCyCydL4DBPo/dNBJKutRY92X6fUSG6E+DX7fUiDOfFhB8kB9IY4J5JfuUhwbcxS6mbWg8oRyFa
6NkQboVuG8OdwTSreQIDCzfN9m5PFX0Sd4cA1ArBQF1Xy9LaMuj0h3NTao+28mqK9uf7QzPHm5UU
APinfCE7mq4naWkmtoLm1e0piyNWfHTHLyHKHOwMywXMMItJ37vLyygLEO8GiXZZy7IcI3aE5QaB
Ztsx01mvKzpWubQmkrGxxrCJ4wrXdx/xCbseUo323/R+EgBHK6o1kPnTtYjgLF+kL76tvennkQtD
RE3J97deijksXLgbVjmRs0R6dzwXdtkQ1u9BnSD1U9+x2d0RafCMPFkdkdzMcx+7KsQcGiJ01Q0l
k+Kw4P85LJViAtm3bgqyXNUGGzy0faayx2AhQyBTo9+ZfSoS6S7JSFI4rA43CqhGx+IkNkERkp+q
sNMfRwnyibjjk8gZcrJKyDpvaC95/egzpsjNNE7Micw2t4KREJTmjzwuARmCbcY85Jz+MMcdSAwv
2pZKBxWfisK91Oj0UikssRuQtiJDW7uPxnVeLL1oGTyWbJMmTYizk+kxrqKqdBPqrBtuvIG8Djpp
YSd3EA7Ht6ngI0ODhPWSWiwhPBDraG5hvae+1+i3gREPd1tp4zz5KXRPVvdxAe0xO89o82oAS/oq
pPhGQgE3qbJpB1/fdkFgFGfa+V5EY0lB7AIm2UEdnTVKaldq+4g+4ZZYGWGP8+Ize23Z+jWhrRh0
BzEuCD3T9m0iqoKUOlpi1fBdQpFoSutpJ3ltxqEXoFMsk/z9khod9kOQCP2h9inOs30Fq3mmvJv9
eGVo/DxIXPYUxYsl/AedZxj7fKS4ufmrM1rc6WErCnqpQtOw9LXYvHht1ZAEsPRlD3pHHDg4T9r/
UPyb4/IobKb2QlOi3nS0iGIucG3VngBgav2teYUYYwlu7RPOpyeeEKbnFeHttLs4JbSRFTEHGa0j
6jwCvXzDsqu18g3zDB8xykEhpD6j7ktNXsK0clTHLqe9siQl4rAOo0PayHt6LqcD+nmTWxgC6B4J
07i52atVtSsjrqkUbkxr6d5awjcZvwQFp9oH51GVUsfrukLEO5HECjpBTJoDv0eU7BTF9p2QNBbp
r92lhCEj+gJFuHPn7sAcXkHocg1caG8EXg8ZYF5yy+XUQgEBq4Cxd01jkPH0rr1mSVrdgiR3OVN5
2iQeZHW1MMy0TcxRC1rO4s+Mb1q68MYbcWBFP0QO4UbMSYTWqDm0jvI9WuB2ors0kgNa3h0+nhTG
o6EhbFkwdFAGxMyCqRHpYY6tYke2903o1Hznj5Qn1eqKJtgMtUWjNUJW5W3pCE0Dsv5G3Ctp7fA/
hY2OIoocEsO9sEwEm8XkWEmkvMDuq5e3qZLS5+tCdGWi3F3dZbwaf4+CTYuPUEFnuXj97TzsgsAq
T62yKOe1iNClYBXMqfkaRucwQjQXrpPRCsHXpyxg50nTftsBNOVxf67Mp45RD4ROiJjtk1OR67PZ
gtZDNK3dpQhVBYcwzyUzQMqSaLBF1lpbkBDbuISPRiy+J6yZrDdJIbGe/PdnmGK8PAkmeSzr+fpb
4rEoNwImOcSo6kq759IVVNyPqIstKXea4h/IU1/bSWFa7HCjGtGeifzA3lghXFnL9ZR8uLvI5LAx
0N60YVbuSVwNc2HAdBp41PL5Kkbgxsmw7NTwQFMOlLjDB0AeKtfWsRm5uIxdrSOmCXZ+YWxY3lNv
FroeMKFJEbas45MWIULL9ma83sCLEI9AA8NoRRVfmo0y71jdyaaBmMvH9dGvHDz/Xzxqo226O7eY
3WlgY4rDYhV3WW3nDvh3Daq3xeU9OwKUqphnJ7Yez8hvGkb6D5nXhMmwcTcrsOWfDDaL9fh3gfH5
eMQJijEvNiy5PdhMfNUi67ONkuHJi78s7kGVvw3NLug2/MAsdtY7SCi375ukfE/7MBI/bvpsiL2W
VOctFUO9FXV3zQHVaCogV6b9iPi5dkqE5NyNx14O6530Eg3GHxmrhGbCu9iDvKbMo4ferrrbO3ni
Hzi1gjTtA6yvCuEgonlKIf6tGGX0ZDoB2xE/uqTf24qkE4K5nfCH7FNrLrfAlcE/Xo3rG10mADmi
GvvjOPNahN50h1Ca5nm5QsbSHRyDhW+a0IfBLeC/9oj92QaQsL8LUwSGeTbkEOkD6kGUfY8XtBF0
1ceHXca2bIhI+3TP3SpcrUJUsMplT/MPPp9sfRVlvEKwdbrsUZg8KYhjM/yATsuXhm+KMg30fJM+
osmMFDiQ2lKEEPpNVEgEXdmy58rkWvu/rpzoI7YTppbddFolf3dy7sdW0Ruqag+Uar57zNn7Zl5H
jYku7lRrrBnJCQJxPR/54rbtBQ8XP6ttSp7LzVif7ZMdKhpYy2eEjFUcT8DyuGrItiBjdXo6ohI9
zV5q4WU+gNdDMDd1mnDrtz7bmL93iUl3SS4x63jab2MoqNjLfuWuDXmyXkMXzF1KRB9rUuSF9dKl
4naB5+qBoRJ6K8Sy0MwqxYDi4hVbiE5t3KC5QnSUke71INAYVOFzieG69g/bqGkS0p5owvOF0YLN
GLIGfLzRk+xOCNtJVZ4ttS1bJOHSzE0cufyeivsRu+un0A8CMLUzIFz4x4tZJJfBFbHkDLLhlp0d
/CIV3rUh9QJfvcUTvjjVG9eeAcSrP3DGeeYb1TXlBkW+sbsGjMFbsEOAej0DMKvQXlO2a6q7u/Hn
YfTveRfulPAtkDjDiY02aKXE/M4CvEnt/oULcYzxohqHA1QaMiT7g9bJMcRcM03iPsWOTUc1VsLZ
3p10iciPglPmZ//7w8GGHpipjuey0etU2EJYDNYBGuNVcQlSyZVs0F8ZL7dz6JV5rpHDIftUF1Z6
SqyT/8me7/EIBqcV0HSdhZvcfFrfY9LQMIu5fOjJofqdLcQFs38h0jyU+wg4bCTPXsOohywjBLSM
PzwcYQfflORRM0wsqG0W01ee/lytKE+M7Txn6hzyZancnKY2y5TYbXJUhIi55heB7yFMoF+UvM3/
mGM0RchbCKFUwiW87yH07U8xsMnfJ1Z1UHq8IwBMWMFCRFT2bsq6MKGewha/WEDKKvpSHOo8ecff
+vaWfJRXjdFHZLEawy7s6HfXEGl0v38eLXHx57Ej/11Ccmg54Au7k50UoI/lkSNvo2V5OGZUbUWQ
4NNuhl2n87WlQaU5qc/8pAVc4ceUuex56gQiI9dgB8A09z2ywzwDsXTgYB9lExhjG3CmiCzb2Fyw
b6XNcAVgpbEHHUhYuDFHFxyNHqhqi4E3FScPz4Fgo1+Yttu9zLMFIcHJtbpLcQDd9wB+aTSQ28Pr
GUR8Ac05jWqVJYEkKMYlLhS0erbRehlFgVI7dKNwZUxBQyfKNYdewDqe8WG43iw3RICIv3LlaXgp
Sir4d6pCa/ohK6mPkLzE5WeKHSkFniNrJTdeZCT9YFTqjrY8ejjfMIr2EaL/QipfvoDdGYgoP5RA
Q3OAFYumuUfJqL1MVbFePn4oOz0pC1dvCOnOPw3ddcYRBwKmd8WIrZDD/DGg4jEC3dDPo2iyhIRN
PxRl9Yeujz3ov8tahO+FH3DR8GvZw6BAmwb6suPGblIrE2/zmb1Nb/TTRBaGJdRlSMRPBRcZf7hR
RmlvzkFVqVcRf3lugEjFQ4Ejjs5FQjpHLvLg9MUZZCPNv2S88c1Fz7IoJrQ/wxwkBPPJmqOvPYba
iJ9WuG5ZTrUWLFi/TiMY2sO/AL2LcSVa9ZyAsumrk5unxiwF6E7HGzYKZfur9gJEc/WUHknbr1Iz
/op1gK/l8qg8WVdynLqYaC4Aet9fNMXLYtEYmVk3HmPxYYfC+h4j8Txwe9ek3pt1naFalvoaAxnq
2T3/REG6JKjqb4hM/nLMBgjKfaZewAt8dhsHOcTI4ZUuWfaMLolxH+8tg5w36BIYYQpx6aValTTe
4x5lbMvtnyKGPSPOuHSwCA9Z1kCOASnT3BacX5a6soInrcYvFqldAFdl6bkHDqlo3rf/iNjYygrU
guvbug07omd3u2zFL0H7b2CsLRm6R1U/ZwL+jW3aWc2WKxt5AhYYcXvz//qlXjKXTOCYA1BcxixL
PHXHck5K/t2m2qxp6sg4N/ruLC0n6itzF2p6pICbSu9EtpQ/VLtcW4IQeYId5j7TZ2lb8ms9WOrd
u1jRb0YhmrHaHUATMv5yQoUmxQk9ISdpbvpPU7TdEdedEzb0n7KDyKhMYDmUoYL2+gGdTpu9kEf7
d6IeXr90iBDMO0hTYM1wGAbwKHGRBbJEAtMhIH7pIIIz4Oy5dgMKjJxnnLYHU2ke5HVIQnVCf8ko
X+cklNzScJMu7wPG1cr0T5fL3UVRcnmlkfS4gLcLq0+UtHlvvMEPus7JckxobuhP7XzIk0hXQVxd
tKyhtXh18UNQxPpxfRhFXGdJRdf1z8g+AGKxTNRorEtpqDyaxmg2+TZmyG2DuFAsahg9bIPdolxQ
P+QO7XPAdFb37aAMgx7P2w6PC2nzCTTZ/XECMTRyxlNO40vpbdI91/LtBt6bcSZgBKRmZiP8i/oN
1k/mwkk/1bVPuI6tEzWk0WuIZveqO4rfNLfbXqnOflR8rpSoa3yPX0KOpv19H/wa4dK3sSgZKrwR
Z+9xsVbkOswV/vbjcZDncPn947ZC4unjLqMg3RD/qneU/V8+DI/sNGLIEGGYusNJcWe71XFry2U9
8Yem4JangogXJ61OgOttjmf2Htr+OQNMnh5BhK6SCxbCPrV7fu26psArkajySj5w/nJ08OwJzvD2
GOCew8TKCGcVfh5myUsv7HffIAmrC9vbLjmhChDWHVltCuMFrrx0r9Ae0A4wZZWHya61RRpxgh4y
WADIixMCM/JlDSWk2msJ3TAVfeP/h6rbOSuHhYH8dosCLd7LqkoXLwikZjxkRNxqSMgCaII2UppH
6w8Zd+M1Q8LQADQ3V7lbFkE/b8zL08MZnyMHtcD1kDNpnzFTJK45Nrk0Jaj6geI+LEvfMKnAJkFA
OakWNrd6ZWKdNCjM6G54G+ici6I/s/Ko/zFxtEz81zL5lgFkacp+UuspmPtzgp640XTs1RoBrczP
VStdkba7dkPvmRKBldSoLD5FBpugR0W3nklTgQ1An+9cSorWLmLllNdbJHCUqGQnWOu7J+T6cjJQ
mm4cY1vI/V/+xOA1wh64twNDTAYmET8S27ZFz5k2Za5yb4l4DG98wvkStJWgQYDYr/pHTeAngC3G
m3EyeucMBJzpKWPCy6AQQiQA8XbhuFwVjkpNkx9KZaIJZyvx4qSWxFVl1oVVpbpcuWYMbvRApIWS
GcQwOwIMwUG03Wa5bhHQxkHug+U4drrTXPK3/i+NLce9iXAxsu9csoeUhYrKhA2tnoS9zsc0+wND
PzKhHvBrmt0ahyzpEsMpOUCYtKBz6fsaW322J/6pENErLopMmIpomHSY8trmSHFJyVueCXG5py4N
O+L4chFj0/x/ArK7T4pKssUs0N5lnVfIH4LOsZzZW7XhFNCN8p9auzaIGG+S+B9EmWt+WVFkpl5Z
FzGsAlH28roYV0t041uoUnc3kmn95BrGoFiLwOKpcqT5Lgi8YFow+knotYnXV7V/MtSOxeyOk2WL
jPtviZ/oSxnZlA4SkB4dX6ZXL/dxnllF0HT6zFIe1BetkvjEDZ3uI73vnHpHTOIN5gCHKJFFu/5o
fJQnYINk/eJmGUWSgt4aTUYVuYsRaw8zuZujkw12R6K5tC7E6GlLEzIjo57DD1gglAw9V0XlO/EH
mTDIF2wIaFNNHjQQlbvAfHqAFzHJBlNYwobpls3hiq5+6NzG18WHQIejaEGLgDQa2L0NPoZCPJfw
X+8DLNqTc7dQX2GiVTw1ozZKKE8Yy1lYGuRxDsBYVcbiwmgPwxYIOlh7Of5W4IkWrMJtweujj8m3
mn88DbYP2VLt+BJAiA/yQl028cMNaykpBQiWbbrAH8FyyM4Aa/crqnbyUaaubcJMJHQI0kyhFJJx
eTEsuZeJti03FzfSzAN5GfqoWgGPATQWPtDmQBjhAcYSzDAdcnO8AxyyReUlhUli2+diAPSQTdCC
DRgnZts1ouX/ufbKDRcqpEsi0IX5Qx9KeJRaMKcVD3mIb4znK/DtPHwVzOgwrvYM8Af422eM3A6g
hSCRRbb7/vtvqQec9P5LL4YG1BnyoT/sjU5yaMcvt8btlsKWeeJOizyA+ZmSL/HKtv0CcIh4gsDY
qWbyUDrs5dB1RysoCDV2mFGf17fB/5Z6RSsWRDdXv85lFkJPN9EQZrjn9sgFM8+S1LUXWssxKPVU
YZKrrjWyBVV11KMdzmWImBcRcOVwMdYjMfpu+rEEQZcPykauElIjTftYwqBYgcsMIpd5Lg8SfHOT
vlWs85XDns+JwJAMzAsEmokS74DpMveLckGbjdo5MVdT+dUyXcaoYwinKu8Jd0O946shrY8pQABm
3OmNXGCval8uAgiRq1L9JexRPk/F8KF6iRaKuwdmYQ7U7Oz4XJ1CQNrLXKuMa0s/nzfBxaGTt7Pk
AeP7VtaeCzIHQ5+wGym53PFten5I4cJG47idaSwFExPpQo20HWdEyQRt3ufYFTl2ZVi8k/w6SMcE
J54zsTSVnd0e6zmK7WmxIqaFTmhT9NXtyFrvJG+AfCNnd+mJZN8mdFkrLIgfOznml9Myph5tbZXW
oYpV69gC+w2FaizkHoQJjqrKzIZJ0v497xqqgmFWk7+EeR1jm2XDHXPVsmtcew1/2SeqAUHiv4Cg
bsD6SM0HOBpQgc41MW783fbEECKQreengjI10gk8rccSvfmvc7kdbyHmq8tWDaXyLmauW0AdGmQ8
bxYo4EdW8QDx9N8pVwZRF0n39Z5/OS0b1RnkW70n3zjY6ksqRjzpJUN3s3MEiRJV8ewS7Zp0KvXX
4e8bYGg5BtoF3xqio/xPf7957okoCNTE+oqP8sOE8mEC906JoS/z+7uBL9DIFJmlLEWvFQ9Q6g5a
9ET9mfn0qi8Z5UdItnL+5RnyEugdBMmzLuvethvPnE7wKZiuJBmWU/3VVE5EdaVAGNev/PZUtkJl
P47w8br9azmFAY/+ETibS28GHHe9SsM1LlCwbw5LfMobOcwDmCGZNaPA0AjBiWVi6VeWGO3p67C8
sAeHsm7NaesZQaUQKzUJ/fD1gWSG/u30EpPhxJm3eS1CpCPCHtsrJx1FFKbsYXZ0ZJecnjvvr4cd
mHWnQJeDPEPOPWwY7XjMUWFWq9ebfgeCRfSPFANzJK0IOeQazv3d7QOQalmICSOB8Jd1gYVwy/qB
c4B2IxLXmJxrSUApKUAWBWIz3gl0Q0RUxJCYkDJh6FLic/o/a7M5MbGFQfK7VlIKMwuAFS6mQ/UF
7oCLGgLunPvbM0JLnbslz5uDhnm8PHPOlDkWqjMURIFiEDqWEsEDi9cZfpX20Aqe2Pe/Pugfvqgk
upnmqmWJ7/Nb9PoJy6ySjOZPgs0jyWLEuETPwi9hqqKhpXd8Scn5BYE3zl4UmQW1STKcbdBdt4Qe
cehXiln35Niq1CERgmBzMy8NnWjTQDkGPFtqQN13PFunQPUzNIzo1WhyKzwwAg4FgNZU119xBTPm
UscqZt+KvcLVqfSICcaTAvZb2GqnF9rqAC2eBra1QV90OCduRsVK3UBK7jmzh6UuTGgdF7mh7rCg
2Jfka+cqqUTs/OJjAUCRkX4x8ZOSeFrfZD58BeYI1lw+xeuh/1EZndsoHbl1y0mXB8X99jEtQ762
RFig3Wi4+43/JkJJ6bApG/UR3LSXyLKW8HaqFr1Qg9DPFzSeuUK574s7R8wtfR5qc7306PQbvAje
3i+BeK/77JIwvzGR/zYeATJZZuofE+UEt03xEq08vIvrtD7o1pB8pA7McGh8LpN33e3/PuI7hVgk
7S9TPsLxKdCt7AkxmuPjltDRHEdMtP0P0Yp9ejTlpHohTxRQUXg2RsOUI8nAn6q31+L6FNtpgsFk
FsMJht264QX2ImmxGJzqPpQ0sxlam8rEs/ZUk6aT45ZjkmoQQ+2Jvlvg4iLlr8ssNShTslbAX9dF
uvacJ4jrn/nscu1lDbSGMJmHWRZQE86m81naKhtTBbUIUg3eZkwIacDLyaSq6yvDaV43wCJjJ3Od
HpSe9x06fe7n67OFjHv+VKwjZXuJxA83jcjblUpXC1gMtokJQTGboqOcPAZAFbrO14tu5a5Rosx+
GSmhojWzw4MHSOnzid9t6IysSjaDAlV26bIaSBkYZ89MDtqeU4hl3H+yMuUYZoM38OayleM6LaIw
t5iYLZgrFCx+fsBaDBOQsfto92AbWm3l8VQNSe2jQ4ollQpqSsRDGN0rsPw0HEMZjLLkTgCliI1C
r39l3RvRJnbMKJTvaoFdNlGRwzx4QiSIJLLJMVOi1JKqL2OS5PRWh3SLl5uw0Hf0idYzjWUHVdDY
j3LgauHORzv07da8fqDIh0aOtBJ7hTp3xHFBeRo1EkYvK/bFep3F/7e2ArkiroHlNxVkfRhX0NF+
/xY8flN4MT3mi+JMSxrWbufM0N4uuTiFkkmdKHyaiwHpkm6heP7k8fijobUTqoJcGYgXGgBa57PX
/YKnr8QLif1uiCfbDzpyVL1CMjejV0/yxF4emJxF71tBqELDY8YzbdTn/tieaEl6/l8dIfvNuEq3
wjYGAczaINQxHk/baH9oR+5JALIR+gvt4WcWuxbRGwIkPNEoE3LKPP19mxsYbzraNJJhjh5EMo1N
2HiHlvbaHLbBMOa6799d+iuG6j6Pu5qZXaJDWPAr9yEkyCTcjkQlCki9o13teioXTEd6+FTcsN7v
rLCMxDJv+R2vUFyJh94040ARDkqlTWXE0fgo0GlqmkTBCYge5lc52g+64mV20LmG65ZEC+cFDIeN
rG2N7OgMNpZudEWjo0dMRJV4VnYRyEtWIkA4xDVEDwewHVC2LjmzQJs5nC6AXCl7TvICBQOqQKwd
8BwdyAmmRoz1VsKC5giZc9VINfFORdWSGJxjPRrLlssayjUtV1/XFZLiALtcLAzu6rS3aC7nQE4a
qr9Ptt/V8p4X9nmzYvszb0QgrY2uD64vfMFSmVUFKHU4nkVfbMDORkmPJXEHdsQyCXwH1bATADpP
2H/guOXYXFwdi6Ud2DBs4PevsxOzyD2iPDPwxhT1D+Y1nT+yK3ymxy3CgeqbwZ7iRLCLPKKWnVDr
Pxd/tb8c6+9iETXebMQw/VbXSsUx6Tb/edm61bz7Xa08TLtCZqP4n7MpCXzC9smRE7IPSexxb4z7
kRgE5vyDTBJrpzWSOfiyRYnHGWaJn9hf0P70FwB/dA/b4Ysm8E02IhShACoKLsoS3doE5YRQWAKM
p0rEQSUIngvuj22Hpy9TamKHyjct0pIix+6trx6AhldhVSLyWa13gzzee7qLsnUtzFMTj8MaoaXZ
ECUBo4NFFhuKSVf2l+r5WyXG+kgOvy9tMyXLfyJyNi7NEAeDWm4ISEl2v6OWQwATJbssId56zFnt
vE92h/IxXECuJy3jrcq8Kjx7os0ZHEAqmgoL+T3VhFNj53VUwQCCCSdz9T+GuOYih41GoLpeNeMj
b3JKDPMIA8Qfy2Gkx2zgzF4bZjiBSWCklS4ds8pdSilW2BkBgEVDx6DmJWPI7Lj2qM2e5X+Q+WmO
tuwymlRCfD+l7U2O9nQFTuYUfCNFy0zd3ehumU2mb4lfIYekT9WJDYf3b5JLtZse9gIgKAH4gk1m
T6C6hwA4/sSsjWeLdAWQ+b86GlLlfvmPn7c03uy+rqEq46jI502x5KhCBrE9jOG0a++X/JN5DCNL
WOTqoBXri3U9VV9sVtPWqEiHxIL3eZf/GISLqzuAJeJhYVUuarAxRP1rYejCIaejA9gd14Q3kz6O
ZUsw+R7stfXldACNPUU0x3z01WY47Q2tJn/UwkSdi1Ks6vV6GWQhVa/Y8hjuYHrHwSs4jyIU7Jfy
6AKmdoR/1C5aMwxGEfLbmLDoSaVTZZjbE57aneCRai8z1LTOAykk8J09gA4HDdwAy1nRE64B3zNE
jloVzciU5Xp8jaDA2KJ7oc4Ss10Z36KoJShjsI7CZP271rV+0g5198arjLv+kv+wnBVg5f4DkrEd
HfwbD4vkwlRZdZvbkis7IbFHN+z8rtmBV2rCXOiMTUIfUAdizFD25H+RBykyoWNjo8U7KSgOM5dp
Zy+UGB2wO2Mhvaq3jYYthganZNBU8AebM/62wq7fI23feYZLyB+OzI34jF8yzb/ByjpbOwlTmt3+
7f5zu60tE6Ik9pzgEU41QqTyCdi2TuGVcx3LDujC80tyKESbNd8kTIFw+fBANehHLq2AU87ULrvl
nFJzrqnbrW20ItMad53SoO9K5WNhrd2eXrdxdIP5VxMzorHOcIhTgULh9ZcHMPxMlmG67BfQeFAr
nqHpiSBkoyfkcxA4XzulQ4yqXUC0xibEyVSd3SC6dPSAJ2B8gPbZokhobVboateLjKR2X44/nfok
NbVSWBBIaFfmnON9++ayJcntFNDH/l/8j/epc/45fr4QzRtwogo4DuohNuSfxseiafiys9DjqxwU
bEoyx5Sx2alyFtOKjnjZx1EIWrAvSqKOH2V9jfcjcZBr1HP5ogEweK95xELHahmlkMJsMDK7eXPA
mcZMkuWoCUvBVi+KMMLzHHTIYT4tmlTl/OiwfPkXl0ew1Bmqr7LCz7FpxwclgHOyUPTjXqSQC/Zk
pQdHX/A8Tjtl/IvmNEzuriIrZmoaRV20uTAQwMTc3Mb/p1VyJaKCLWZQzYGcW2e1pil/NF3wE4hb
ZmnxEveLnx9TQNBtEmtHf5GRt8dDHaZD7Z5Hq5iCVlBKizfvw+P9qRnRWOoK3Z9I1LGb2PARcG9Z
RjXuG+LC8uWw/gtpTTfHGTSExt5V4E+jNPjyLRUsbMgnTd4IVhv50Uij8XAKlHLToAk+bWec1mWB
6iqFtGEoJDUo0+2OYtbkJn1D1ZPLMFx58GbK4Z37QAR1wu6wiuhwkZaDBIzxXMvfauCbCB4aIBRH
vpWDAVCR7CfIx9wMpflLKdArh1AvXpP1dk5BbwrX8r+PXbd7rnun3yph3ae4zQAKrQyzwqgOaDSx
c0/fAtOZaxDg9ARRC+wuAiyQdSlIwDh6QispZ8Fb+pMGzott+qNBqOCCvG9/9BEShf0N+i1qhnW9
iONF+xZkdqKBMjac+6Y2nBUHUEbXRfDM3e2M5zo5TPgXb8KGDoiqts3cNkZ/crNIFvbZjldpwRbY
97jo5qTV5WBlPCRnic78oaRvgnSlQQPuFM95nANeMuDO9Cn/8/2ZeKOsKs1SROf6Zen5LTJHVBGM
zXLFsltkwJOGEFEKFwoVnQFe4ppb6ggvhvoMkfrCyE6nuiNFdOv9h+SC9W3l6eAzPxBu9inDkf2J
IwIZpKqCF9MfwcZXRGnKiciNryAYzf+eVlkNc0YEWGKjJ4qWol1Bs1QYsaFXOmAZP2TbaiUwAPmO
THVj5LMbA2PfrL5idB5exwi1qMwWGPbER/xuQhUQXwjx9ukyT59jJUih+CoUhNbeB9kgk8D3vjWr
66WYrIgkz2eEqcjakNWGT6XJujOrSATI/eqASP2mI2wXWST4ExYA5OnaUQLm9/F6FAZy/tBlXySo
D/vL4solrRKFp14QwsQgPgW0oKMZloLdVMPSrGp+eIIFR4XERxblOzREjwkFObe/kAlRiycT3ZTv
uM+5akXolM2RhKEr36Hbdxk7AEF72jRfpk7SMCcEnQRLcek3VEMzspnfTkpBlZwJwTacebAIzjda
aAlSSo1rGDhe1KKeeO/HP98q5KqUK9Q+CkacO+BUB1GhUqh4JGRjNKiYTKJFnc0R08qmi336gY+F
FKdo9LGeB+a5W0ZDeT5hYTyWfHQXg2fabW0GtSIWnqVx7Mld28icrHyb92RBFkcd7EEyEgemfX+y
ii261OMq8WdjWAE5bsAD6Uw34K9bvPBzR7LQz50fYa+ijTspqTpXS6xIAQhz6RsrMtvwyRW5Rpdg
J64yroId+8uBT8Sz2xjH5OFqzVVgD+W/IWGoZXYYav+SeJLX96MPO1ufZ87MB+NnWp/mBF8E+PWu
VI8Pl3CCuRWBRfWNukC8Yu6RspdAPYMTOKftjXd05W63JVBL+iBoB10rvkub69SnZA2Nd/98E5EC
pr1BM809yhJUpzUPZIxv2AyRV0Dh07uYRk9xQ0pTCNrbWkmK+ZlPTghNZfuOLxDtbGr4X+57gPQp
FEpAGnlh96Rhd804UQ/LjRR27satyQw7nbR6XFFdYd/9sdP8T4m3gQ0Gtf1TzoX7cnTXL1KB8aZu
2pqK0mFbsTGoJD0z/QpZhiy21/ZR5PjJcowbN1XWv3kISbDxNNG0ZsRp2qx0HvUv091KvZW+Z4Nj
GNhdGT3VIsaVkknxvM87idyz0OCQhNGVTYolEvx02ehCPxUTLKRMK4Lehkg0J2yvZZmS896sgfF5
MaQMpSOnBsz0zZZXJFyNsFCJFXnLYZMk4WIYjQMAWS7SktKEsTOXhrnE5sTxtG1aRnASPf1b9XVj
fEHARWwH48GrVUYsVWmdNGhkak6AE7Id0UpfgGXJXIOMz45rppJPxkK0F9HSRfLJoWa3b+QTKO/d
MtEkBH4mB6J7Kksc7iCFlTTnMZPf4DJ2vnwihWes/jSlT8+G/Kxrx5LN4Pw6Nlh5v7xZF7td9WJG
rJpyC3Aq7ZhtwLR8TOiG9WU0dHiDZuP4C9+QErMJ0WNqkB7xhAyz0AZUzizLn2qyV5nzHXQ5CTOY
ljfbJDOTYhYSDeBqNbpV8TrBr3OYwQqB/7yDd6sychMU4iaH07k2djBxEa4eOdNqhRIoIOOxOdcD
xC6FfNLOa9s+dCxqOQ90p/l+yiNiV7qg/4RF0doXQTvZHpYvtj82sI6W69sMv86ipzSh+Gho7I1u
7JYknUk08iYagPQexmd20rOD/1Opb911w8g5AEr/ZKvhQqknArarvz8fNCgiFj+el2Zm3NR6fIap
wLFjc6WvuSRnnglHuSaZWnvUy5ASoMVzLlBpQr8mzsip8AvaCoUD3PFNkQZWAobc9EMZzJR5RQTH
82I7dPJ7g7xc6OtTy4kQW4BqmJeteeGVVu0kwDeHZKzkqnSy0EmlwQCH9Lv0fLj9PLFDPpX+8R8P
BXX1CEXQbuWpFeBDMMEFOOfA7Kx5jd+vTR5Zsf2Cl6XskHkCDAyAk46fkFfyMzoMUWpJ10ta2mRD
XLf/VHvgt4cK76jJM+9fHBKXHZnVICnojHOxdCP9+D0wxgUBvs334yiXB1pDWf2VJ0Xf4jthNE8N
KEo5pPZLydP/H0t0phent2sj9+EGIItVsdX342hK8nTfV1O9sJSwJkkd6Gyv7NIFDOczOgSLupLN
N91Wb0+5o7oWXoU670BPgStvKaa7Pp/j4fDngFpEEZTTcuHqEK5eaBkqW85/qEizOH8paCFJsUtm
IKCR7zlutOeVBFXYBzJi68ghoRs/+7bZPZmgX263HKRkKmmPO8+hqs4VazKnUTlzbfv2xZo2aT6w
nlwh7tE18IgDafOGleSLlwW/mJHWEYf8ScqGUm+3eOY9AjzoRr1JR6GxrSAU92E7VeiXHDUQ5+O3
bQKnXGe7yvHyyUINzo9Dr5qQ1cJvc3cz1eKVe0DQZomH9RbLTeecTBh7Q26NqmhpPBocr1pwwDe3
YZCbZYv0IEpaOijz3p2L1QgkOASkMMfWUcLscH+NahtBhZnL4hiCmcExqi3ml7J7oWDUthfr+8hL
2BHCzUXTj5mQn6sCgya029FdHx6iB425wIk9PBsqy9PNHxnYlx5Y7ELhNPGwKKb+lwqxjrFjw+IS
DjPHlo7WrqQXK8R5Bo4sCwd3L/iXwwMgvDP3YYxdjpi/0OAC5p+PeXyIzM+iO3TiV5K/bZdoPgnJ
TYRKuenhv2ztlwSVU8Xjy9cdL2SsMek9MuWFePgh1wL3SSQ/O6ncrEORvf62qT6NbjOK0n6opK6r
p52v8Q0osnVuG2UsyndLbzivPjkLzjd5wNy0PZicFGX6ZvbwizZ4rAxsFnKXCbZw1C/dEiaPt8X3
jPI4ndWwjz2KGU4OzlyTQl5Yl2f4ioOd9gUrEkfaLMn/rwycU0fjrZdJ7LLZug7TFw5mqbJrZLPR
7jtA0L8nwSKx26pWVjlwQXrYfND3LUyF32EiCE/DvMPyTLXXyHDK13jetHa65pBBiLjSRJ/AToHp
8Y9bjhLr+MaW9Z7f0lXkl10vYVsTliI5SmCK/wFh4AAp4Fi6J80imSjJrUtMVtGnmM9mj8q8w5Je
H/Hrzx8k49wVjf4lZzLNn9yI3ZmhGol2dyycuj3FhzhVEiamMR9FuTxg4SzUInCM7iiYqMOVksvP
K5rp8Fz2DtGOEdUj3fU6VRjUFUDbNDuH88CuEQ+6/v23b3njvL0QXC/GZyMIf00QQv2UyJXicj0R
IBDd8xTbsnuqkFNyvYhWkuf0Eog6nfBJ2+kpk29lh6H2qvsZFZPdPjRHrZx84zswl+f+8XBEjqH8
8IAc/rD3ilRoJtVVHaVewsPR1zv6+dHtEvDv1yHvcddVRwrKrMcZuLcfCSktVEsdbsvGgXC+Tz4j
ThHIfYJweFx24qgsAJUL3mp3oG03IkZ6WQ5lnbtCrseTb7mea4EqhUlsKckBCro9x6/TTdDs9inH
gBoA6Fy0+vfwjKOBL9u9FG7QHBNlxmwmYC2GNBbapOFZvgBtS3yhP2S0K8h1WSaF4gi/Fztpe87l
NGEwKh8F79pPcIVRX8KDbsb5+mlTDiaXlCzAzq61LEDcbUFQH3Qt7drp/aWi8WUVo0ygrBarC/jf
s2aEXhoEnPRde84e/tiAAzS7JdEM9Hs4yaKGqiEcmGcAup8vSX6chdfFpSXhFkWThZ7Hy4ElL3Lb
16FWoDhwKgGlIP8HYRkM7ujmO5HxKw0Dmr4h28IWIR0k0qcm55X/QvwpHQUCvCF/HZkLRcpYTy2d
ACo5D53WaHAj8si9d6gytofP34iUP5FtHh5GFzS96zMlt/fCIj6APkzjYQQvBN2vT8KE9d56qmb6
myQE/9gkMR7GaX+CHRt9vvfAUwDz9U7RnjfyRHFw2cQK5Cz56PmqRSVVJfwRhM1PYbHVnukhBFjy
60+4bdYRTh+xGFQj2wlLme4E1Nn5k42gjFXkLxhbrxGCNNdHwX0JfzDPf+b+/DVAWLEb5GFHctlD
qBxWfjhY9iCbTp1QHovU5z0OAyHgtXRpFZUQ0eBUOGgwsJwTpnBhTwAjiwlK9kHDRfJPl5fEl+2s
9LfeJZdutwPoB2+s777ThBZpK9S3TSdZa6q/2/LDwb4vxaAwiN+3T3YFpsk14k/uCkI3ieXse0LS
2LsEUw0MBcpx6W8cIANYKqVU3d7CZFw8kBJiY/G4ecKG71SsOlYx3mjoZASx7CXLgqOdbZ5IcDdl
qOH2vaxSRzmWVT9UHlXmh2z+1x0bFDJz+OJJ5YlnzAFmh5BppExtGLicIw75UdsMSOKsCcD59yYa
apeyPuzHtM0y358icMFFbxfV3fzkNOw5GSTFT0x5F2/NNUckbYKCLgHegoA+PhYilBDX16GMC+At
VCcBqyyYKqct0c6nE7qCY+fRbQxw6Jsx1ajYC9x0khjpv0aYG1MNqdzwH4Xwm97jrr2YAiNRAdkJ
5NW5Xp90oT1iy/dUf5y4cq1TAEgI+QdZ6UKxubczjcXSXF0izFLOWu1bbeXtXc8iOgD3nJOb3g0d
Zl1xGnCQxOrtCR6rbTAVX8vrFzBqXyT4R/A17VMClr20EDoyBItfTw/9bBECmme/X4MY/gfuhZq7
DMaZGM8Y2IcBEY1Dqwg9t2XjabLQk7fp0CBx8FAdbrbmE6LWSxCAfj098wQ7w9lgZg2TX2fo+UFS
RfLaw4MAdrJxZUlqikvH7MxGZ8Dj9KHZzGMD2dwgUCnzGMUi3BK12uXKogl4vDh2lMnaHHRHQHY8
+ZRxka9DZZgX2oKl8r0SwN2STKEKk3zqp9ObHpDwC4Yjs7IFJ2/RPstbseEE1p5Czkho90t3j5DI
rs/BqcTIapo96IuBanPnpCjPLtfKdZHmMrzV8+hV5y7bZILx/uNX6qzv7hH3fTA0Ds5pe3A2svxa
Qtw73VvyFb07JXZ1VbM0ISYQyaDq/fjcooaDiyz4vRrPyFwWZjwgSWkk8oH9BqHW6r6oxf99XtxA
8elhX/x8BcNNEh68W35wdyucWlI6f/QhOhC/ZTRfTdbr1cYP2SUtD2pEbl0T7Pf4zZMmRuKey8nE
wuWv1uhD/kCOR4p/q8sUkph8VqMpYw6D1rlD8wnWRJ4ql7tcBgN2oy4TWW7RslRDtpYMYQQs9R1E
hQO5ChJVqqDZaONcGXqMF1yJyhjaxP3RWNMaBz9rTvi9EnSKDACwrZDCELbvSPujdWirBccVqbV6
5TNH7ngilxWBt1kBuHvcZ61bd4uVupatlrdun5rdk9OiflFjCjF2hr3iBZzHd592KQyQ16BcUqlY
E5TxzSnp+t7OwRnGb/yWDitzC//14kZutiUOqDmxf5lToCsKeF6Bmpc6JPlPEE2YnZKvSLtt054f
pEiloQHE/GyYnPwSZt8Q2iOVfyMhGxjY8Dmp6gUvHQcQX84sPn7M0coW4j2kLYyTzMgpe1pssk4V
4ImYEm65J9XdYqwxX2fM8X6tAtIjlkGdE/x8aV6pe9eYNv622z4YMAqsbZ3hfXq07Wh02SYebCbK
Xlu7IPU1IV3FL7D9/JDimKYzgD0LVUSwPGauauLLU/UWvD8z1kScUyZONpEIJQ0Q0QxL9JAHcGwv
zLQXeWQhjtJp0mv8KWfIHFz5zqlN7onrYTCopYpJ0+sofGHYkpKo3+I/lWc1/J32kecW7EwtPf7t
BQT9MUICY4zFlw4EUciwfVG62Tyu9BSeRivDBJEa8trkrI7XAsG2+xkrJG9HP2hGp46pfMBILdK0
QahbbC/cBvqoQpL0bIR1I4URdXEMKDLfzQuMrFvqPVWXO05NKzCFoR7DqidT3gdkiSXqERlYhcKu
xNVLgti5UJFp8rvyK90Om/ugCKntX+U8Nps8AmF0xvm8L56lExk62UvRviFYStd8l+hTdlAmXLI3
fNd8FkMjUWm9HHGX7okbu5Xngfm1dGG9nS8tIZGIcO+F5AKxeIS/BSteCu+9b2BmaRqaRSDdLwL3
fbiSKGl6+FXZRpzA9iiUYkyFxKhIqg+V7RuZCSWL6yWalkftJUIaWW0miaVnRFf/Ol7WYWh2kVge
bHQaqRh/Q3qPQXpb2tNY/gs1Pk7gXgVBHJJU4hrhS58y+NbjptrUtb44Nkv9CwlaLwmyvKBkPeuX
64Y1MOsoVhNlMUmnXt+ALfb0/I/Sdh11G6wU+FEKLUNec/Xy8AXunTz0Z+Pd2l5e+jtFGuNb7V2k
pwToMU2LEtZoGnKHz/DxJ4UddWFyjN9BeL0h+usU034uH+9zLZcSUIsbN3wjUY4lDfbhnFz4Hu3f
xVORpfV1blmA5DdlHDQmLTblJ/GO+/IgUvFX0Lo8UrqVVmRwhIMdd+IJXnAdbw72DHmbDkuBCAog
saXMdHmqAKRiyurEdvpJYSSP9gQizElE5Gpf1lhSc9U7YsXZefGC5Pvlr11Z3yrVGpwR3MjkVatz
hCk/pBgp2i+76vm4+4t+QuFjkTQOyCU90Fgk0ybVct253wS2eY36Ynf95r65JQVi9PYVuCrmTAol
c19HuNG4+ltS8nhcxnfyOK0g9+HPPZEX4mRek9Ta5En/APoHiZw5bu4zkKRYeGvLInxTggv3/hU+
7x8jK1BLQeG5MX5CUnR6Y00EZT+OxXTBfVz+DSR3KZV/Oi1XbwaWu+m/SLGQAbyf2clZ1MnLBNIK
GLEDk6Y7IggajXRqTw45Sawm8h4KApdqWBYfNNACU10ApsaukykEz61lsVy4u2/hM1tITWB+NfFC
wheCkUnwVjrImS4VVHGucii+pX2ZTZq1A6XtsOn10qn+iOezuLbBV3P8peNMHdWskwoijiDVTqRO
OGrat7leONvxAHR+Ti4x7XFIbhPto6k4mfMCHEyYGtOFrMoGIZ5D3EBepaUikf0WGkkPqxUlTJOS
mL1nEV3s4kaJNhAu6hptZba1XyYq/2sOkHwPuMbsNjcTmIQVCSegb4hT/8Q/Jojh2i7ouJ8ui/wV
fT8AS4SO5ca/5r05FTYQg+Q48axINEVYi1Po3bLtBEzoUYKfbNhxmrqgjt13Byqh6tdFHszuXGcA
tyd8+q0UfRS586LtlkFYA+rwiqP+eIl92JP4wzKSLd0MBNodJiBu58yj0Z+ItlQGN5clebYalOHT
Ak+10H6DVvq/Q83T1duSfacXdJOQRmg3HZ5QbxY2c90lPGQjpYVfJenkQ+61BYLa0b6tVffz+NXf
cxRQ3okCM/L8k8QtV6dHSQIpPrHandXts+MBJaWj8xeX8f2WAuaA4n5HYIdpGPRdCbv5vt8Pd3+y
jOz571JHqG1JYdhmzXNqCh8HMKnC6cg8r0uNMUrhU1oK6PWCcXHugGdH3MnvPB6jjO6aa0qVPRhc
8lhsq0S4QoQLMTHYlt7MQ+LhX6ch59RjuLUC0o8B+QFivH0QEZII4u2gfJ47jFCBn5e7x1YRy4n3
gxX/vRmB+KfGc12+hIWh6cFc2Uf3/sCpbcXYZbAAcGHsI11Romje33VjHChQ55zxCSAU7WNnhaw2
GsLjn69dZKbkSl9RedC5EMjdSEkJ8hX1aMUvu2C9is181i0RJ//YC0ewfpdmOdhEG8r42D64LQgZ
ixkXTDNh6ciWBB2s3LtoGB2W9BX4Yg4nGAJQYtRnael5xCJ7Rt9RopUIS0Cc2m7IZ0+Us7Cjv1Mq
JxPsmHgoifzfDbyykihPmS1dKf7G01UjnB2fETckanvSjHEO6fXAMxzsAj0MnmjZVLpP7F11i4XP
KdGOyqyCI06h29prjqvsFvHZsNORE6b9iSnqTCm4KmOwq/P3eA16weCrR9VyvhoHXCU8UaxF982c
Sx0vh775nqWupWnIQxGC43tQSZeZMqtV/ehW833yHzzU1/afnuLngt3MtCbMtw9DWXg3kpI/Z8K0
kA6d2okH/agwArxno6MptdEGVdITnkt77draZV0DR5RkKPrTxsb/npWkD+AZSPOjG0uO5cCP+P+C
lQbbFY11zlf8Jn3wAMmK5O9mqUJy7iCVEdkzHHnWQq9zJjBCuDostH3iMGTCw5qzakYMdpVkAFol
0eeyWw6CrJs3WoxDSSf+Xr3Pzmh1/j5OMlKT2/FE1wh7tNaipuRbtGakLnXod+hJMAOEUr6ciNZo
w56OQ43a+JgAa7AD22rarNljXb4bL0E0z0xz9DbgMOs0nOzE9zFNULUcOGLyzWF2pb6l5VacLHcy
EdvTAjJZzRzQp8Jg/dRYA8uv/YcD0c7B0rFhCn38p194XEg8eZInA4LeN329yn1w9s8Lb5+WniHe
3afBJk+4Eircm9d7x1TUugOaN9r25JT+c4kCFaM+KMETudc4n3UEUV78Z+fuw71ASX6GLZQqWWQ9
7RibwsjRc5rtHZ2wdhIqBJlliJ2MQCUnzXTOKtz1s/9cDcVhB0Tn7hT5eSw2yYsoPnZAN2c/XooT
0Pt12kD5OzobA1HK0ozzIDGwU+EZw1WdBekWDTKOKzDGr7DVRjesJmSTxneZJ2s4WBW8K6to7XDg
NKo4KPc1cg0aqsMXkp8MRsxkTbQeCjPZVcYrQOWibMS41Law42h8EZzxqlRg+ZACetsB1fvg7OXW
drhP3sbaU22uDTs/DUhhBpyQK2gNTFRDIZSS1c6RqqtTtZfvjgPDzvg2uJN2FfP2OEl5IuqBmgc7
onq35H7lODtlmdwMX0TjuQunc29T3P0iXkTZNx+xdfbxRKT2Y+SsWY7rIZMk+XyYgENoKM/VLInx
8aboKJYD729dubEP9wA6L7Ids8jDPOrG++UdYVYQS9u8yGmBTeofRDUm45jPuPVqYd+89eMAxP8L
TSu9Z+IFZ+3uZODwjfoZoIlJ+vzAHBLdxoG1T4onlK1lacRJTz5B2IOaaTPh3vM4l23PDVixNvY5
Jxhsf23AcHl2wCxkPENTF3z1NiNxpxkCbYbICV2pJ8HxVy95L8o5/ltw+Qf1n/KTOU99NFxxTWBW
m9lg0iabbjUKNkEx1VAY9+ro+WQNHqtgEdws2FbkIjSv8XIyS0n6VFg4N4NI5Aju9f0HkIX26auC
eoIQJ9Ld7TMU2ytNCj9mlaQo6VJNQCxxIwqY3B2yazdFcxCnly1ZRb10y03St66qQ5b7tbsYClkl
KAl0z3NI4ebKKnbvPjg/sljiHjXhc8ymkgJrXFwSg+ypAvmVGKtn42K1kvGZUee2opWvgujC+Gjn
6Mlioa+dr1awp5OUzT2pFAWwRq39aPC0Z1RcC1IJSjmLIRAqSQfF5HlLe/lAFaeo6gzzHeruBjPV
sKB+0593ADCXlBMuVKdJHFdf0WNw0j9QQVjrbYdVLZuZjqnJrm2MANEk0qNHxqrnCXisjH1AqUal
x/QhYczykL0k27mn/bWxieihZU9bkcT0E7Td8X1btI0Yk+geUuSjoqUWre6lo3yMRq+Mcc1daOas
lTqmp8pLSEDI6nAWh/xkiLH4Vcx+H1UkX1Sn5GFliLbV/zKnwuwSaZXb2yhZtv7+6EFhcSLYgnXU
0PfnwZEAdUkQjsZEfENVjGAVxaTpwDqnIlZD9FQ61TaAkYakF+E8SZf7RABTS/M+JRdMkgXZ2CNH
KkZ5tN9+w4PVp0CJ9w3ePSMG/P5vasDICsbNb4KiBodoEq/HrFg/tFglXkVYAUdf8YwGGFJ61v+9
bTbG5Rsnc/oSqlCh2FubxlDKlBHR3XYhkdcLANzKlE4ogfuvLZqinCOol7cxIms7iSgRX2mKV3tc
rTqPZftsyS4GAnVx3qbEGV6UPkSx8C7H/poVYmf258cTSWUnbDqZ/Z0yRa1LauQqH/oFRvg7C1g9
9mOxZKqhLz31oA3drvMdl6tD1AfXXGZ0V8KN9QhPirut/Vn3NLPxcP4PXUAO3z1cfm2oiymev0QS
Vo5cLSfgYidQy4Tr0xESM06wp8KDsWcLke2Ntd3sLdIWaK7juWQPWhMM1sdgvuaD/NCk1Fid4+09
U0lZtnWCV740zP6rBmuZe21lBek8isinskQDtz/NHDMmvdnZ7hwIk6lZHxLku9zQk0CW4raz+YSM
PitgvpgDd23Eo69uiGdPZEkSpEOTxOyi/n/vjKIdxQsMBSrlr221ecTlLqYh5WMA7VUs6cyc1ZFy
CDZ3HmN284Zdy2qkCtjoYh7LvUPUyE38NymYLglhbh7gk02ydvLHtk4IC4Ju2lSNAg72inCghGfn
EY7wu5Iox2FRVqz0bw3J4sKMXAb9ALgwTYULYojiGbP6Q3JSnnJ3rtvFOupOk++7XBrtm4d1hscO
8dU81Z6yp4/7n14DtRpANZOBmmlYyA3fHtprdARqwhdayUMVFqCsjt5lWknx8m+xHDSZRlMEg8Fi
gPmtrSV/pFhGxPeJ3TDCxrUGNRI4Pny8q5QN1YEcs7Aw/v37TMHElLpRow2DGW4AB/JT6zNflQa8
q/hWK0Q1uqrs7y07nIK80kUhOtpKCCXUwKFXcTl1IChhtmlUqbXeh+hap9gp1cRxKe0k8LAjNJwX
b2GKpDzOKVtxE/Y8L4VP3qqCmwXeJk+bj+ZCtnNxeylp2ntAhqLgkf58vIO1rskMTOY1oJpS/ZHJ
lK+vCIReJ+5mRPHwSAOe3srnbzyhyG93/aF7YDGKC0rFVEl2eYwG2N6Nl5hpv+9c7WxMO/YoZ/zE
txsaFQH7/ps2PJid8XABFKJXNBi4wiV6J0qn6X++888xdPQrGzX70tujz+mcVFOqJSFzaOKo+Jbw
iDYc0l+tYWDdVORY/W0/Aa3e76eqciN2FjAqrCEKWUHsOMqCHwUcI1JGEKqEtdWj/WaGo3sbhnyD
nDsOyFuRCjRSY8OSpEQjUveFHG0o6ZPxTC/BZp9NieLla7TCkuYMiHE4FnOeA6w9OnBsPiaNQl9c
YZ/h7q+pYQON14Ek+6FmHTzr9rww+JvHI+BMaahJDOZ57jcCX1/2/YAPp8TLFonx0RIUTVX+ZwDo
BZe0vWXR6d/pGlbu0UzEOCYMycTk3Ec2mO9ew5Qy7hEnrLan5PQEvlWyZzpQkTBeNNTfrxkrEf5n
/uUWSPx1eogdWb50a0WJorEnfASyxlF5w/sc4FlocAWc6hNs0C7bmMltUkvZDkkbV11tfYcaIQiI
yPqsS6b5gKiFPN0Jj2dZ3qi3cPbg3/IYLuMH+lhoiKgCfLb7kAndPaaKQd5h95549HrNZZsJhmDn
eka5weQlPSNoMPJ/Y1XZI9dNo+K6XRZztP5axgnpEaZXwnpdBAcyJ30XvAxFu5XViDI5EZKguxfx
0TJM7aFngkV3ISqSC6H1ulBrO0R73VnEfTRA1fBZ+jTipWEorsEv7PcFeaQqXrpMHlFHIIimXNwL
wMFje0MBJn75fOwZTKLxdc7TZhUnBU+lFt6wHK73TeZSIlmh3YYDmnZHKBgVdufTPiOPlkZJ08cG
hee+FNDfVz1XJZ3+JbubXgkUyVfRe3m/6U9icgrKnWqv17KdnRMN0YRMpI8R2aIe4BiAPvAOt8dL
/3/zgtyxv4gYkZJsAzAHt/3eox5+kucpBbPFX1YRw7QncD33qRndSlQHn8eMTnIo7DmjWdn2TJw+
zeNulrU+hX/pHZoXSR2Fn4yxzIV0Z5DKS1DxNup7S3vB1CjrSafl19kxXIqkZhhc2kMnogwQzUbj
A9ZZVfYqBJhIU/vs2uAeaccgt5GjVQaigwqal9Z7wvFr8ybN5RvP0xzJXiiY2gRRxua4hBKsY5Ug
qLiiHQ98DqkrxUO2CXt2fVK/++nRZrOcfuUdVvZHIqNvczPiH6cNWCt2NIVVUWMUlDgTwwvBTaSN
6hNp9W0x/8cCZWFgpJP+GDP6ppb51WQOj8AT8V7GvogmZIVsRpGM5QB+zG5hawRy1un/3SGN8oD4
RFJf2kEbWCRUBd+ItWnvz9EV7CmpVDiuZePWvY9T2HgOD4fkZN/ZKZzzqjLhlyHYeHB7WhYq6ElD
tYjqGt87oMDMkTACCXuBBaSbewtpjo3dDbJ53dXSSBmz3g5uvc5qhmzFqpQ0eS5tGaI6ZKZeCzfV
/s2pZ1M8ikOJvKOlQ117lUG5fFwodX4SaaQTZWj78YGozzizObERDbmFXsETmfJYM/pMloKbuVv5
tJBfRUA5cYfpXOqD6oIfXdeO5gi0UBx7jXK0wyvmHwI3Hi3+e/t9e1gjJuKNd93cZlaidQbZwlRq
2J716Fv7Vdngge4JQzfX4aBGW2CqhXCa8dzAxYj4D6ixrkZ6u2ZQ51VV43ike9CbspShWlrEN7O5
qkcX6Jrj+LGm6I3YBACyWEgtE/TTuv8WY3J00wQLdacQvmyxv8LHNC0rpRUEBubx99TWSbXnvol4
swXwySrLkZWUWIcMPejnzCrUc8LI3iOvqJQXfcxP184s4lD519XUbOtDOy/QmjzH2ZCtTrmfPVXO
OG55Yvo2mvIinvHMah/M1Xjt7HsuwvW2vAX2jEDs62LVHCguhVYTD/KIWop9dcxp2CtyEQTqsylk
DeiJFX84VpFaLoywqxbFYopINIm+/lFcJ/xLkeDGQJ2zqBlC1xra5AluLdeLL8R3yujx5h2L1CgL
rvB6R4LelEu5293z43bzfNyK8LMqz6juAD9oBWJud7I01C9CF1pTFKxKtMU/y3L8k6BbNaEZD00V
L4Hbh+fBV47aeFYBPAvVxZnIgD7JXQL4fco2k/6qFXDV77yA5BnN8y2IlwqI4rqYtRVF4Dok/oKg
HhFbAgJaNvfcn/ZCnVF3egghq35DK3AfC2rmUnhgcPvXATj4K1YjJoKzZXIPXBkOZihjBjt4TWU8
ykTSpj9FClmmzdzz9e6BXozx6sVqkYsuQ7p+N7hE20hx0xO+6dPYpwttlCiJLTRqsTp55Jzfic2m
ZAxpNI2O1OAgGK1xaNscSlmjffMq/7nm4CEoZu3/UF91JGFaXIOZkfZ6E3MPRjbFVQaf78klUJRg
CEPQbQshM80lYQzhGFDDZ0MinIwFiY+YhlHoqRrtnI4MbEuxYE30e1SVMtsZCk7nL2VrWJbH1w2P
ViHG3/gjVulKT9+cZ/2F6ScqQsLICyzYKIFT/K/lYGea55yRI6QB8xRYxevYOY+zPDuVU+CX/LK9
arKVDWONKdDNUOd++JqBx7owzp9d+Sg5N3XMHRkx7K4UbhuDLM9ijTV8qvYFoLN0Gu1fO/LEJmae
oVPSxuR0m6EAhrZnZD3dVrTdXLNvU+/nE4n+7yav0vXik2egUYcaLQhE35wyHrvaE7JqUT1oyB35
qcFQd4XgCngiGSls2/y5vlG858uxoIKgD363PehU7JQmKdbSJ5tugTohftIHCe2i3sSeWDriMxsV
pJ+KKIm2O68HFmc2GGUQPkqLHYF8LTpoBjDxmxvVdl0nnob3FfwWFIebj40MCgfPpi/D/3dwGRiM
jjIeW+kZcL6AVtPj18K+c9mtcQC1WyHBoe1v19I6GoVT6TcEQubZxZS5YdFbJzHCRiSsuvCqzwUD
iDme2W+A9qlAXsiBSuEqeNoOjGihsPZmWaIZ5GtNFI5xXQvZqeezWrIhdYaQPueiedEXN/Gw0gH/
d0WoJ4f5jbi6y0Iiv1C1FYxUrt3tqq4MGg5mFMAcElFtG3fjEeNPQ3/3ja1giKIwSXuSJ1e0DNCy
06f+/Jg11ylA5iujAEodLfLKP0cxlRvbC1rMzVlxO1R3CKcih/PwLIfJDHAbvhpExC7ilBpCc5dA
VV+Ezi3C4SEkRNeMYIx9oocckkzyIuLUXDZ76QRLuFLJgKKYiKGr05k5BsAOQZJ2RGOd3NAMTrFA
kjLGy5pUsVxxkH1//yoc09N9kOc1ysAHPDZAHzjL9+ZmYgQzCwTTvPvh+EiFOkqip5Rzk1zTcJnj
FwHxbToWyGqMplSUbU7uDGqOo4YxresLbhfR+qXaDBkfb+oPjnTV6CZFUusOZ5bUM0W/YtorHjHk
EiQswesAtg8l1EGVt8ieEZUXouP84ZzZ6CV4fkZ3P2N8rZwakkKi9cJUdw7vIKVrq/uFOxCkO4UR
sjYDxjHb+Icfs+Hu9FcPFmFfk6cyKVEy6+m0EdWdG5SnIeTQrQCJPOnPzkD9Rh6r/YN4MZkLtOwg
Zd4KZ+pabv0kW2LATmTkoAmF8jLdBFYy30zsJe8JmkID7aSaFtyymsY6PAsVTISfUyMUTcErJ9Sv
YfjDG5NPMcS0PVau/OJtELi64ienT79vzW6vYcLLAV8+SOyOR+K2u3KflRQ2X8npCuldoaxXlpoK
aN3sznBkU7EC0hwYDsNc7arYZVOoA2ePX0eE8zgyQK74M0SE6KkmeoIydZ6Sp/tWVT9ypnSQO0aP
fcL2tB2M3FEp/QEBBdx7s1cG1YRJw8AY9YbwNngrBel2zi8IPlXwvqz4Omgtu4T+Jecc9hFeaLK9
ZTnAO342PpyaSPxAsuGXfpt/L0z6HIvyoxpDTzbtx1C0fjh2bJL1KE0IDyUZ2ZC+Q0KByEg1yVPi
hnKXyNA0IURPEZuetNsiLscQVCLTOVft0VFGWE/puYkX5aSsT8zeoBMvaIEaYXT5SW5W+3dGuVWk
Mn6DQBoFTAyzDMdoqxE4Nk7HsZCyKHwUJU0DXTFtThLA92SJWBGDIy+YV6USWhHLlkj+ZppG2jb7
ZMtP2VyfMj3p3R4mBJ+BPn3Mv4LMZTkhnHGsBg8OkEEGXmBbEnr/8ICydfNL1G+Dr+Ab4TV9wkLD
kDU8KlqAXYvQ9nH5clYF2XrEF3TqwYdOgV8vljorrbQPHmNcCzCv+3KjplloZ5wM8wRbaerN33yr
ziofUuU2oobPA7ShO0OUNG4Gdbn6K0lPNnyCQw4rylHBCEVunztyTJvoJ3ETSaalehN2U2NOTni8
pBRWcmt0IquVU5pNUJ4lroezijXloYs0mRlResrFVvhLmae9SFzMciVqbRu7z5iPiYMsXscgtfFm
ySdTRGqiMG0pkeDQiu56fsogU7T1lRzUXOq2smwRQ0MmZbksoPmvlLIBhMaWxFJTE3e3xDlYQwpK
/BeUO5h6sR9WeejeKtmil9A5A1do+xbBoNwso0oMv5CrPKRfiQ44cgPIlOKKDINgg2Drwr4AoRC0
h+o+Cc223tVJf2zhZb837j1JXChy7KXk6m4BXdSCqeb+cxD0EX3cVg2hEaxpdszahJWuEuijAz2l
KlElPUZjtuYkFtDvjeTFat1VyPKldWEO6eW+SLIZiJaZLW9brtOe2ul3XeZHUoNeLcc3eYu1J8f0
om3HSTq/SMbsKMr3GfwwTsGdfj/hb9bf8LkFET506WABQIQZ297c1QuXgoMj5f+iaC+tn0He7+eH
MvCFOJfP9DA1PoNmMC5qB8MP/87GS2pEuUKVlR+eDmdACbLIb8zvffFwTqCSMPvSmQz5t69ZVOQw
XWmQdqQpNvqEJ5A3OuOvqINyrEKiLtHDfi/eWL7uYweZ5te4798IRBoswgY9213mRfYx3Qu2XE9v
13IaE00VJKorHwQOxHGkYlBDwmNtZx334rkK9XIZmzsburd4J+uSZNRkbxFsjWcS6itFN+PWcxYW
dnnK37xNHONDC6gWfd+Q9q4yOD0fdBGO/oHK8NAvqZ/HjwTwyIZ5Lt63GXm8TBkUT26HSRayMevQ
VKems74YbA+Hw2uLGKBXP5uHFUdhBqYzTl2cjXgsO60+shxH3K0T08/BDInlaIhRpUzKrc+qJzYQ
8VfE3qJwtybRue2lXX4oc+Umqeri9MMLuBuLYro8AUeiCdHlKDCV3iGW+LhtCJ7xDPWmoLFEBdfK
4qhozKtAU8FTxnLQZPyx+n0Jgq5b6HUNIb7ae7kdaCXG267fI/dQR6FxJfe4m3lExzrm7sCSDwNZ
FqYx3fpOA6HvxziVAMzL04SK0zpL0TNqteOrs4g34PhuaNeW++UfugXtgYRqJmvuQJ1EWcHdIjps
R6aHDPojA8WgmE1iEjovizMUN001fNlPZD6QD2WA1NdmQn5YCIhSm5RNzXfaDIa39HiQ2bBt0uwN
AQPIfMvAnF8jidX8ckVfO0GVuy7EkbA+1wyvOdzv9LoDUfTFBVkgim1EhJiWISEWQUNrLnmerB/E
PkqUVeZF6FvybZK6GqX1OlnQqC1mMZuIhlFD1cTkYFnjtnIH3BVtrACbB5bDesL39rIs2nUG0qnm
nuF1wl8kPzHQByuhd9fjpZD8wwXPOJAiN+3UcYD7p4lzTGia1aTdp4U6luXlKZyz5BfDA4SerO8K
zhDRyodd7hED2LLAPBT33iVaT56KijeVryTGTetmI720a0h9Of5jYErvzyGTO5FJxQ/Yrw3pxr7v
tScXXrQRvJIMGAyboVs6f4MunmA8WDSohDlsL5ubw+20AsYDGO7Cg/KLGkLLd+joRncdkHEBi5yQ
LlWptgzLnk6In1LNFztzBizQyH2EBorcDxkXv6pfgWn1KveU4IqZVxAQ8yUNBJm2P5fdqVCfamgy
P9+X0nYzFXXl9nhwZwqYu7uDm6T1Nydy1cE+zLD+S8WTlTN0eW9tS2Vip7cj/lptMjvU6NoPAoOo
+4IP6X5NHcb3i4MHSi27G+qRVSEYA1LzU7YHWQKRKK75N3WKqlNHtnR1EKaUhNyEomu5tz0j5B1v
RqOif4s3RdU+iDZdHrO7gDbzNyOA+A4Y/UOFviie/9/PQSKVCHRBgu4Xg/LLZtNsgJG/jvHw+VUz
Us5lYlQGgXAKnzBJ7p54Ce5yyGmKr/3KsKlRdJMnPw/irSSMY/0ZA4T/pw1758WYoeBEc6XacmGf
00jS7nL3ly3Ijap/ZMPDzFowxmenaQEed6iCC8IUVtHhkJlwAFPCA0SQcnwzPIywBzycTaDT6scH
brzXSeqva+Nz6KDNY+Zk/7Y35uaSw3axCwpPppyjR1cxTKhnO0O9IhlxyByw60kJ57pWzKOcberC
RU6m284PS9g7cEA0RU4HUQijpstQL+RqE2z3QP/QHAY/bpy9EQmF9vdasda2siwYL9YJ3y4I4PsN
MKsHXV8FuRDXFCUPI9GVgy/1snysbRkotn9fwMEAenSEVgvIlIRf378obzhHIEbVEPmiGPMCGRud
B28LaDZVspioH6cO2A8e/zmIwMBSVyXPaLi6H72w0Zok3vjeMHNLayT5ZitTiN3b88gEIPIK1+PV
v4lgYq3eo+TTbw/4uP1gJc+NESMdV+IzQbgljcWkeW5V0tG8hHfqxP9V3cmE75lV92m2NakO8/jt
eIhty0NJGEUxRjhasgMTwb2H2HoVvCppwuhgWck70QZjkdSN+7r1jkycbQFyu33FOTp5YAnvkyDX
exOVfru5o71nLmk56B9tPVjWkQkWJtkKFojpdHHUPwSD4X4YI9fZ8MKOwLlxxE2ToOjp49kKt+wM
tbCfnZz0P0+MNLKizvfB+TdndGKmy26pvc7UYXjQ+FAoWky6E3ici9aSXP9IIQ0z05ZPM+FxZEJc
lqwePyH6pset2VePLEtV3mKb0OOHHLfqrmRSFT3D8y+buprt5ILK3eocMSkCa7H3mYYYOuv4U9pj
z39fle+NQmb/F5WyiVyE5mXEbTQVifD5cTGF5IODZnBjWqDAn19YATo90ZsSiNpugO/W6VYSFlQ4
fLGnrSRUcCNnESkc+sANbzK74z46YW0ku90y6CgVlpOvYaCPdmQZbdlahOzJiCH9bK7Hl4EOn/tx
pN7peT8Bt/qFH3rACvQbTCdhW1VUF2gCdlsZ4AxpO83K2CyI0GBeq/I7xe8SyxYE4LT2VdgHJXZb
JpqDKaXM5f6oZzSdXvigLdY/PQHnFBhBiOCPqQ96a/TurTK0TWZ8c8wHFbY3FpxobJizvgv2lDtz
FT8UBkNNk9Mvx+UTuStc+2vgZNKExLIR9PBPxbHzgIC8GQYXlFVD8fNW6MAHgW0qDmEXvaX0GZ4S
a449GZgq8qiXVrN/38N/NkGrB/UXVbNdRAWyF9wg/ZySBImVoYj9D7o/S1vmEnARE671dfIsNlmO
BUiuPrTSC7pTXRTmbunT499yk+D2NIrTjBsGfKxKK6qZ09E87l/kG2G/UowiSDDuoCTkxn1UUG/5
bbF6w45dIwl4/eoP+wd8pLLDnZCvGqHzfVyRvnq9soTh/iQ0AIGOjMgdXS50j8sE0bhlCFS/8A4T
HmwBBD6dwNa7eu/pp2xE4aDzpKBlzgG/MQA7XP3cdS2J6mNWLBrlfDvWB9JMZa2TV8gOtuiaOKyf
tkY9BnxyoesipR7LAl9e3SofdLYwXFmL+zqstoMh+YhauB1Lp9Bt5vwOyT00aCGpcqQTi58TYIdS
a/4N2uIbxRDdeLZ06blrTbgBlgOGJKy+fad2Wm68F/wig0yFsYWjGygzv5gC8QiqFxnWpxz+Y17k
HWq8VF5zZ/WJ1B+CSRDtEysta8oEqgvQRkanWwbcpmLKyAztTmTY0Sc8PQZv6v/6Q5/wtl0/kjZs
pElbjclTpyzcISZ/fsE2uht6KeunY2o5SwcuKmH2Zed7hT+Iga6cP0T/XAUoEU29RZuimIT40BRU
qQnh50QJ9OnfPhiyN3euV1L8U7ineqIk0A9bYK+/46pMrv0yaCOf+QP+PXVqql0cHustVioCJWB/
CiL+FA3HmYa0SA243g+ibzrtcaC/016/J+428EW3hbYB0Zf71GB8IK9ui/vepg7AS2Kyi5N30BmB
U8/aAA/H5qU6FqrcWnl4N74yf39ro4l4Sgg5TVVd1w/Tg/vzwaSyqoqxrWkcWKJZnaVdcvTtwxiz
qM+q3pqNTPEO1/KC4kB80L2N2Bf8ItHwFo4I3RgkHCwf4yeNvfNbeMtqmX8swrRoJQigB5bQmIIH
XqLArs0MUmDH0iHe9fzuR4w1c9QUxF+GWsUkPdD0qLGfdD1EMu8l+cfAyh6gJzh5q1uqne/ZmxFB
8w2FCv+t/2zpblc5KkHSHqnQbGGhY9F1jrjP7/fpgzXADleAl/+0+cYFZQSXcbB17AgNNtUMHkoN
GyIbowe3RDf2+snDWH4fkNusyNwucEK08qLn9nMNNskxX3tRfIiDMbrh5/jcMYn6t+U6hwXN7JB1
vBE63sz4Hzl858h5CKEjuU6i+ny3mqc4Aj2C/ub+ZIodrAy/rrrwIDM0ZHUlbnRP4P8ZopZqS6dh
xmha89SIP0aoLorXGQ10tyiuVUKd+1fC6wbZklTWoXqo7Mv6Rr1zIIS4MUW/Ku1gkazWylaI5chQ
UZttFIZ8OidNpnWI7qnU7qELIxn9BBgUaeZF6Ulb3W289oQ7Yk2gefnkpRQER+mOlAcqjSeNbdLx
Crf+Z6QGLYZrS95YkkOUgroHvWDEMgdfH/oQGEbqdwo4s8TtmqarkDLxGX30wR5dpidjf1AVovto
/ozOf68noEBiVS1y4gTSj9hCqItjF2rUqf2hSWIo3PQ0uqSIostVEmEeAjDLmX/2vfgE2rZEOnI3
7es9Gy8DHDMwo+C8IPex8nH350xpF5cCycSPjhbMg5/AHfDcPppMMAFySnVebQrHll/ZakycW8ej
afXmb3kZuWX0sEoGonUBZrYvARMfbKLXTzPISoRP9W2PUd4RREdflU6Or915FtlUV2PgtCvWPcKJ
34j1ced7oMNSIYKimeqzbmIYM1mzUeDpH8oXT1Oc/gIl2y/7tf/BkneeSFoL4H2+ngrtii8w0e33
NCjMM1g73GFsvAa3lNkFNH5K5w5YO7nhQ55ije5NYMsNOfEq3jhwy/CDs6GbsQGURVqr7sngaT0J
Gha6L5ZqWgXLpVmnpXIUTwms//043X01x7Y3jDPzWyQGX0DRVi0+vIhgJ33QTbNyqFjhAEd7mtEI
F2TVcoASqf3kT5rTj2cwVmtGZDAgrBJojHzovWBoPF5QcXnG2mQzrK3PGVe1JCaRcig7G7BSOdvF
147+sOYQ43y9/IafnJpcnCy3EBe4D2u0v0NChIugjaXDLaZrpD60ZK4GlnbWMd8qqHehtZKakjoz
gdti1eb+66zIPxbL9rXouUR9XnLcN3tHjhxbu08qXBh9vQuXaB8Iu5DhGbHjCvUoaOIXPyeayQlP
o2wY3MCWvGajRy4u2iP/OrvgiHSQQwtfnAJfgMemOIydSctGARkVUkysO7wQEW34rD1hTq79aKzG
oPKxE8xW5z2QHSgftZp4L9c8pw6MFI3JyzMj2FfNSBubh9vAYNWhl5kZeSQvJ+zR28g9kRiT9bgw
Yc+5xb0ZUQnBblZc9L76/h9YG4Ltq930xqigvfc1JQiV0TbxgK2/ZyQFiIoVWMlrOUD3qeW63C17
cRDX7F6SpFqJjn1ED99TnOieHThSGPiE6H1SMDMxjc4hkZ6zVkwQeeha2ySo+lZcCyX0KikHHpA/
X/LyKSsydokmUE0JPkUBsdFdJfoJGu4WmjafL8PfQ1dB1tUY71tWhx6x2vX+O3wiyVm2Df1lHyuR
YBPN4AnqGCl2rJaDc4yMXggmVu8x+Ekvan5kKUxu8IpIwZb7HJ0PRYMvpbGkpoozZlcLdX2iP7NZ
UpTLqiUyTNFDbN+NkyAjmxVDMqu9dbRzmybLIy511L2H9sGy0TQF2lEUCxHKgus9rE1x/rY8s00c
dd/x5W1tF56b3TgWRpach32Cahxz7efC7+fKWfY6hlWiavn+b1COT3IT5SiEaqd0KVwDDJUoA5IQ
e6XGIpXPhOqa3mvXxZX3X0+XYbMm0CayEJkQ8QFm3E6RdZIIlOeqyc9YqcEpjwlOB9/xOmix7faJ
t2zXjdZI8jxC5GrJ4cqzFcDACU+uYgMgK2n5Z23aBllLiOMYJF4zZ/W+LiU8quKkhAO6tfHw/5mD
yzE/ChKp3rgMj5s3e1tBbsRg7Vpka07v3E+5GBbBX1TMHR67lE4/4ix9vpRg6AfQ4IquSK2B+i5i
Pd8KSXyQ4EqroUGQL0+25iFpMwnbd70SxHp7eRrwsjhah7S1clXC+BbYewAFQcT5Q4K0fGagzvLZ
jFPbmayGcjga0I9IyqRZQL647m9l3s7ZdqGmblvcXygUniSE/qBMt/jxwe2Hc1fXcH5G6u1WTWSt
HWV7aWjvha02CUXUOAg3NPabzwfd0uP+94Y+mn2pqhJBVHAsr+RJlVfQeuPzhg0SkykfB6Gm16xg
SCPE9JHosZNYVZHNnhdewJbHOoCPTjwGwIYpxs8vnwZimhae+ktxyz0nzMSwT/Qny3nvrqYunBs1
4/PD1J5wpwyrZw0IrCWXJFD+sPqJhS0BYej5mXwuMgHHDt6ZaXIsAVRwTrpnbn7UV833sfIX0jqH
rP434xkJiESvNdJeNcTlJleYEBsOtX9reEJvm1pLgaTgSI4O6nshF3EzqPYwPIqwKU/Z3+N8dvom
q1MsodLFWyKHNEqfedFsL4IrheguDXIfD32tL8bLZjiSIyDZjYW9WraaPcenX9vDxbDSfjN2g9S/
zzXB7/kWA2en4S/G2li2hTF1OOY4ayq9q9q5eYOZWs1SEV/b93w/btxIimGQHAs7pFla6O3tzO7G
8ylCW763spd0tnkX6uW4iaKcRvR169x8FgaVOxlrZdX19ZEAEUrjzv+laI/9gt2JD8MfeWEHd0mD
+V8zhm3lIISAU9mX5Vc2HvdbR6BfhYJptAhbA2ZaEdvzFfjR6brfdWTPTd/2fKOvobYBisyQOgb6
4yEcfXzZ1rayU9Bb1K7hSlcI6q0IiLO+9DMeSRSfuVqK4xv6Ge/amHEDn3lAl4HxTvfusWXfTOJw
I4KjAI7dFmMfATIKcH1pNUJ5OalB5PWNMrnyoy0UNYECw8t6d+jB7M2rfEtQpw3XJZOLOkxL6xY6
iNSGv3XlRm10IP0/n+t15yONY3pCek+zowrVsVpqj4Xtnr6RZVa6K0EG+Gdz/R0Qf4TBJ7QuEh0t
thCLhWYuf1/bXsF9NSrcPUN5vIczjY37V6eNUjSnPrzqZL2N5u0BC3pejPYOAdUWMj9G19/19bww
VRfLEHxi/OJM8zCyr8TUxfL7roOE3T+p/FOkSNaM3/CSI4xDkB0uVEFbjzGgRVEkGivycbLYr6ET
T+FXdTHe2ctT1OcXdMxgGtleFYHHWU76tH4c7Z6gozpmvZf5hsNfMWf2YTLPLsZZsVNkTlKrJh8H
8cca5ZYXWbXmsBJsQU+lqU3/3tWgRBKc5QcxeYstMkGHbTRqLGXS1oGZHkGxihj5MWaoQCxeLWcw
tcDxAd72Cc/JlVfqDK/UCarnt0i2zIc1aQoNaukdy8HqlI3RjbL+BYCqy0UBxNXqpMaXrhcf5A3z
GinNcSY04kQyV9cTAJAHrTUiT3ZF/XOUTAvNYLRdgIgwafLixnUFe7isnkfBRDecFql7y6Vk21Lt
TH6gQvuql4I5ckqm6Lf6rcinvLKrAhoudfPMTUQ5F8DA13yu40S/Jqzhx6Ko/SUk4EaFBv47U3vB
guDfaYfOq5oeOU6dLCCEEpn7zpEAWsSescdPsXAE6EKoj1IwWOWcWb3Lp4MvlgpPY4VTccbjNzeb
nPGMgfNorZNxY/Iv4YX6pGSzFZ/fsjIVvuLJunqTWemdJbbQNPOPNLjisNmIt0TBqHSAheTwM/Na
Mxl0OXTiiebnxChnbeLmkWXteZmArcOeBXR933Zh/R7uE6kmiXXmcqJzQKuMrpGKin0hRXkqwEi+
RmhdjXXFB1v38PrOW+j2L5iOeENDb4OceVgBSWYMdomVLMVy5Nmn+U9zelMH0UM+qkbbTGb9wTQB
NE4tnLioTXReHd6eeLJe0UNkV3TfQk9TjSz3cxtX3Zrxipvb/6+MF2t98WFnj4qdhLNsBVECTY0B
DxLMkWAs3txnROY0151sFfyHxpo3vabhs50F/LGuKygS/X0FVFAKOCFhjVIX+rU/2KOV10Bd7Vj1
ocCS4jkujIEQEtIHh3khwefXztV9hNSgayi52bc5y7HqqwJY1tL/sqxxTbMAwtliGzZpRNqfCTfY
FJwzZ4pk8TlMknG2T01x6p3vV3VgbpffvXeMsOjSqSSkVBiv6Nt5ToSIcrPFPrH5eZn/1Mqz6do2
sHbbGVmPmBZBfRV1TAi+UoMnQKpaaFLd5qpakRFYfnge6jUGkaojA5TymXiFw59JNYdd2xncEzVg
VRDM12nm9waVjF9J7xJkEL+o09C0etmFWGQDTnXVimCcpkkDtBEk5hS55IvFgmZmZg1twY957/0D
VYwVX4ieapEKxdREucxogeis5VFv+rzI4RcQ6HUJSlxiB3vlZDM6/KzQYQWxySaXA29eZUqRTlnQ
jsHPr70Xbgxv8sWFIdr49xsorQ89rTeh3u8HG2iDz3kQcfMcdIb4O7BTaNJpWs53n2ejTyhLqXlG
910HLv9X4yBYVzg0WFD3pkqbQqPwhSiTpZNZyvhvWtCEStxvvtnh/Uug7zh7jQWzUqUGtmIxNllh
K4RMtrY+0Dulv+DK2j/3Xhyzg7h0MpulB92fnK1NlAwoRnW0ZnT9Vjgg+U/W619PgMpFfyDz7ekI
nAQR9Oupf1ccjUNWzFrnrPbCr9zpKv315TNIF/orfhVtEEYQvROMD8q6mwnY5nJuRXns/D4tH6Px
wCee6yfljJUX19QBIm9InAQ9nEJkfTw4AnV9PF26TmiaiEamBRGnngSa07wvQ91XsaqRzkuIuQ2u
VOXuiftyM32eC4xTvYAPW77/Nt1UvxdJI2GxFKlxRlZoe7wBtUv3B/D+dc+qQD+9uydx/f56B8da
Dp8UymX8JCADFoVM6Ff6em4lLpWCVI7sjJSIcUWjCyxc5lCjbbfkOjnncILQVcyO8x1rlmws+Tp9
66LcA8bKPkjlVKQHMh3+Q3Hj5vOqhVVa7QdKpw8nff0tdxZUQemvina7SiynEse4tWwuTifXE2a0
Nq9xo7P2Ibau9a8fg47tq5PXhN9DHUcWcfBtJ8SSumRc3vCkq7pcEfIrWbVFWT84eT960flsQp4A
Uof0rTt6HLG76cNMH+MUFECRMZmy6pA8jQihaXV4G6IFY6V9pz1b2+FGVJ8t+QXTVfiyRwrs5GJL
Dty7Ww/0wq3oQgZGoO+PxPKzkWqGQpWipLFIoQpp3qMeAK1/E+ilIls6iLBLAeGpcYXe3bdrbb+v
hFgs9/9Yhz+0NpTAEFBuBGrwnQVP3gE9aeRCLuv1bHa+1vgMjMFriWKQ7odGU5CX73GxQimLijwJ
1zyM9kVbFzFhmnF5u+dOhrOP+N9ApUfCtBu5/CHrXUou6YywUC+FwSelxIXWzfghFPgJGCa7EtKZ
Tj/cF9zy5sh8o7XPtvO+RV3raEPdH3hlaUWlo2nqIigUFZM4GjRTktdA54C3Q3ufC4xH7+p2ffah
2kqyPjQIbjNzzvxa1UwIsVAtcg/xy1pg9G6RJPoFw5Oz+f7QwmOgGeuYuccfHcn9QDWmc3kNt9AW
SSVyE+ShUUJUy8N68P0ttBH3HxmWdeuGo64AtVHhpm0emHGcld9yRznJFjlbrZV5XGFlBGIgfAsk
Gt3Lkc+opZfd9OUdUUubVUvN9MVITrx49wJdmq5+XIGG21IqK2pKm7HFaWvAdjEQk7ppLMMXXnu8
P1coCvPGal25ulE0sRKwQfoHEQ4c39GFfDOHNdkDVc9DqVqLPpcS1exAfcIanzNsbvIvldRRo3LN
m2wpZPP6K+hkohpnnJ3Qe1qGAE6wpBTGA5dng2udJw9T1b+JnqQVap7MdcnXi1S8+X+W3TqtNVQJ
sgIEkVY7kVvuXeIZ9Fvm+Dg9S22FCbfwz04P0+oyJfxLxMjH6auiCKpLsk/0EGtbatN7GoU8YAy4
w9iPApl1Oa0FO7c6Z56btgMxprVoq0D3pQnKHJIhfkx39C14ltdffz5ZzKykMtKiuv4zJJkmTPOc
MMiS+9zACl0cfxH5e50c+aI6xft/LxcTkI0LV32FlDghqHtJkbjA5zxL7q0LFrmThknIiD5Ix1WJ
GM+40EBy/3kqM/zpUkLOFFMfDBsgmdkPlIBZF/IobsH2Y4HeqvBXH5rJFNug675KcwXvkHsqVhA/
FuLCfHFRmNu2+F9ybUehxBTUDtbRP89vSXuIzwQnMmznCJ3iDFrYIis7lPGebK0i1vGmS8vqYuTa
9Y0OwTJkOqoTcz8HTtIt77F2aVRzswxh6K3PuRpFS5Lfap3UWUuTRMeReyhWgJ5xQox40TV5yFOl
O+tC/p2iUYCVEifpT0kkz3wdb0xXmQvxEKqUQEPi0obx2lKRuEUswBBX/gjOvAeGMihnwrhbqrxb
Tz9NvwZzIUuNYYy8lMWz0f+Bkd0vkHP4EDx6L62GB/sFIHmLiPZpVJBkvgPy9wmuq+Ew9ojS/YZH
GDoW8qqoxf3K4PwP0BRPWTEKq1eujV8a3TCnbQc6py5CXSKFgSrr2cQXs7PsJlcKsieanDiLk5z2
pMCYJXEbU6o7fdsnApnMiN6Ord13S3WnFsJqwtqpm2bcqJpthlqJO11dokvHFBsb0zNrIJPEFvoq
22nOsIAe8RT+aUd/a9DRF254G2mKNX3d/pcty/5ALJgsOWij9W+VC5soMC8Toofg/vUje2wIAoe6
DnkKJ5iZ/W0Z44zaWOGerEKhCi96gZ/ewqYvFgtlYIpx1iXpiWJagWMVWtRBs4smxZFLAEg3UcGD
J/TDwzyDoytNPpbxHyTK4v2+uzNbwgNfR1T1Bygaf9XbM/wB25jpm1BX4TiaYVzXvm9jit/3500K
nhCdaZXvm+lpnikkR0QzZSfgZ4qD63ZW7GUHJ7j0qSJbYHTZ7BwtmsWi2LBca57d7WbWbfRvE+0r
xoBpntnhNzsuB4pI+HidOFDLaxqT/g5KUb+lZ88A9Cvan1eoYYNpeWv/7S2jZeaV4Zku/vsCvz7n
jfGseFll8cycGvUb6iVRzb6PJlyI0zT8/A1+33rReQjdStQ086vx8vgh4zQxFkK9EEHNnpHz8MX7
XA6+uy2ffqRR8FqJrgeT//nPpmmmZn9Ibh8akjYPSLIZ7wRziDPama83vd4skjSF+yBHG6XJKW4h
kVd/eg2lv8iRFyJheaiXdHnPv4n7YjUrso1D7xTEcjNSf4W7wa7uAn2xijlFjDyalwA/KwHii/mm
58ZosjqY6LQdYOsLzZLiY3oLWzw/wO7391ZpFP4LgL2MAFrbcIkq9/P9K+J8IF6dgIYMN07KZMRv
RyBEw6Wk6U2nTa9kGnjXPUOCjAqJP9gAmuRTmooVWVrvMhbCQT7Kde9uri1sWuhzT0wR6YgqpQCW
FI1zNil/OFb1t3z2jPQ25fRfZE6k5mlCHePtL8S8zyYf7uBJZXUh+CaA0bOHcdiNgmOAfrB2kSXU
qEaetIeGtXhg9+wGIKATwXvdM5TlW8K19cv7W3qYtKzKFHlR6KAtffDmrW1ztxVYJqOpFy8VH9SI
/Q8/OSzKW8l9WmJHVEQXwREMC0FA3GwjJq5RdY88krC3aITy6cWupEr6Yd76/Uggq6W2JpMuNbBE
yhztVTcswR5pZ1jYDTT59oXBlZKz1bV2PCeG0fRa7O3c1ytO2hbc7dN7o/IEu+KVWqHIdKQjN+Z5
xbqRUYH3wnCMgcJ4Ri5nNPtjwJbxU8GXFWS5Z66jTWqdR6ej16B0FyYQUnwuS9KEhEtl9RxWuq1x
MvmjQs1eULaf/a0UwkU/I/jXwxe7XpBGmhLUs8nRSjv6swZ9GzJB236ti2faWuZJTLk3eGBfJevx
C1k4IegLem89fI4dUwz7icm2sabIciQKadVa0YcTUDhk2Kf40lglLquB2dmbKju9rMpQ+PnHoPHx
vhQLWZFcwt3EbX9zPOIIkGV4WTGDZUEZLExMSf4yiZ6DA4sFY2pGjVJ496s/yBmOLwjS7XLt42qB
/S7ecOSri8kcv+ylF2nvc0vMxRRWUJr6F6y3fwMoQ0W30uWqynWyh1EHm26oljuLc+k7GWeMciDn
NBDwCEyLr/wgstfyQ2RmFD8CMGEUrV1eqxLqQ1bsQuDEGJzTWsGrM2+dAWvDKyHqiTq584hlaJN9
YlkT7IcWXC3NILIwPjDg+JWhGafVk6KUOvNAo10q44HgWdFyj0ohZmbm0A7H5DWqfJyNKPtNERCP
uet1MK7iAWv0zo/5m6ryHWqIKWWVqVZHI0yjNjqtfUMxfvZXL/nJY36ibgs+KIOkm9makgDtfqTY
qYzyd6Q2XymKgkwlag0NkYbUYQR0ULLK5q+rueVW2liOxqTr8TFn1wkd+ZhnVYZ9Yh5t0Jt5cWPd
/YuiEERz873DAZve8k0CKqrovaH19pBskMR7w/LZOxHLigR9ZvPG+Xsz605bN07zOB4/jrd5J0Mi
lyD1dPPtyTZStLX706mPs+fbdtZ6w8/ZDMllJ9bqkQ/ZUO9B8twyimGaJw5OSTIcHq3fyxMMOIz4
P61GhGQT84Z9F13giudMOCpaICmPVUQkGOkaBl3kXyuzvQfRPBECtHTyVm1V3pxkDSZYUPC9p91Q
L6yV9PjXOprwT+l0cQlRPpBepMhY13tBfG7OoRCuJPIcWPcYPCEEYq/XPnyVKTBhJiwEfclGKZnL
foqNO9tZ82zRCCUIZ/rtF3yWycxLSW+nY42Ci3OFoIX1/kgNDhlH6ldd2KWHEo0syiO5UNUHp/tn
BC2ElzY8zX5JGM/B6f9/owVScPEylyDoCEqYWvqVYot0gAlwke0SUDTYuVxStzWpujOCPNMEMeZE
6NaP0hTaAbSSoJhJMmf4tdzWSxvewFoHlVKanQi0X7TC8dELJAcjrXnE+Csy1sheoz5wboHaqhfH
c90ixN6axQlUepFjSQBgVvIXbpAtUFOe8BNd1VtCQfOdzPVBtXlXYzK7OBlBL5o8ibYMODKOksnh
BsjO0961o+9wOShv55cZhRWdaVMq1ffaOnS3Va2t9nmguysT4BJYxevgeSzRInrhVLP9F/Yo6UwL
NFozP8lb4oDA9qm+JTUb1RNgIEJnvHgt/rmvIKZ/dlfVfXbRROEmA45Bho9QbHOns0OOgEUxqB0T
2wdzbNsx8pmqxqQLrqfi7BgB2ZgodSlPKiJxSWz/Y63Y24eAWOF90i9GeGA16s7qYSSIrxmvrehK
FwSQwScA0Fc0VBrhn1H+QcH+nGJxkjgtQwYaunj4xwXHuHCWvgB1R/9g1lZZFIXFitEiIGkxyPeD
bij9ZndNTO38bNVgSYEQ7AEXTzTg5MMsF9ZA8tZWJa2UGOHidYRcRftNb+V8MxiLtNxnu8ArUM2m
e9qonSwcQFq6Y/OaW5CRQlrZl2nGApWhmCMR7AmlCxdDLadcN9oGVickAJM7mE7ijp1YbxKkjLHP
CovlpMCEnCjspDJDxD7A5IDo2SWA3Z4swP81s1PJF1truO/W+L4UibIeLkdc3X9X8dcyj4J0Dxoo
BbkQs9wqzM9GOE9iG/gHnCwcmKwLWBvDQ5mhkRfTc8XYAFhsIDnjuK8kQyQSeF+fq/uSJnBl1nDG
8/vhJdkxm92O2To4CmEr/mwd9Q1PZeq51aOpfq5TXP8uYVWMQASRZqLw12k6VwktAclGIYfdgHx+
EUKVynr6zudQ/UhmtRtHTSsFbwubhz0N9lruaqvOlGBRMN0tqk776Zznr91+jvE7rxkCHAvVcjcE
fRb2GAkvaKBn2HLN26UOhm7YbuhgSw/Licvahrc62Tx3Y6wsP9ND7jSKugisW5gntkDWO1bIQ4Xx
yu/0r4sCYLDMzCj66Z74i7udana/NMnUzjUjbjsYRNZopdVnUSCsEtcsGjudn/v/1hRCUJarP3qu
CHWT+0V1rAGWHjzAtUUKGOUrnwPZb5y8AeLk9U4jU6UMP3LHTsX/YP8srfWDBTLtPWgXCdKX3v44
sXkORcE4AdmqIDSsfbl//P11kUC5My6N4B+wkExTX8sWwBVGu955WzG2LC3oMB0xLvvyJXir6zYB
lG4dMmhhe2gxSnltqLl5kfMMFFWSfeFXlyjmJR5aXldZGPJPmRSOFUFxLbztr94BxvWmcgLISXjf
VprYM4U/6h8wGEN0fHc243IkythqJY+XsHViNlONEnbZHjOSbgcx7U51vRtj+rA58nVLVR7jJ7Z+
Pyk82kKTfpMyVc425Hf5wuehT/pHR89NTutspsn9/DamtNF4+HExGIDUu0LakLB0nA44p4+8WCTm
3bOON7TqpdtI12KZW2HkJIDFbRfCKSt56hxlv02Z+iD2TVLtATOeLsKsyiDLZlByzNdH9XYiOTI8
s6hNsLTATrUbMTfnC9l0kuYTN13v5hQdsK/VVCRJuLkiyznVvZ1PZzdPflC3sbDdIuB0eevRbJ28
8fcjvxhIxR+wLHTsBjXYHvaQQGaZHbtu7enHpB+xEy9qOlrfuZDVyye0xZ0RsWTpeCXVV5zVl8Cz
aXSTL1RjFBvUREbEEfFY38olfIsWXdkeXC7er3JT5wrF2RdVxUA85nmc1BpEqioUHRLP0plHiBmW
GAwcaYIQZ8G/EjTrj62cBDuN+f7YGwbrOeL0z9VtIfbDxMTIkepBFoZszAeAoqzzC5JX0paeUpYa
zFuxdvso7atlercYjXkrkiV0PkvXtIUgruQTARtn0NHMKVbPzG0uDpRpQsMf0IYW90UNvJsooGP7
BUx2Voa94Ip+xxKU3o29oqhWZ9SXCVUZYo5WspLO0PsgxYw2Ig7aXV6ZPmgWAb7rt3bfQpK9mE2B
G7t4WXPbvlZiro5PAxMvj6CWNxyM8vDypAeT5EN5sf4NNV7rI5xFPi2A8+eV7c1jyupGjkXWWnMq
6P7MzYWeDR8g1Vj3xqeNRySjk8QA7H8YB4BmURx9HDPFgiXgD1oS3tPRcXi09fcPCAI5NRdR9fYA
KUIrBNMCVyJWaSHaH1z1o/zM7wvlQHSOftpLPwK9BF7rPbSbluVKAYwYn6hsXl0wcOX/YgNhEWAs
uHxFLLRhymjBQX0/JWuHgsQXuR3qz2SpemiTDFCVujaspzExTkda5dNgRYac6CdBopFUmTKAb9sX
ry2oxAlIOWGwBUwCVFTAGXOJI34I8diJk2xgOf1Iwv4gF241r/j3+dybMWgTs7/SjXWzIev5T7bo
hKkSYrp7GfJaiW0aCiMJjYn780OfpwIEiMYlAjnDCnOXVa6hHsaGa20HSE5Wza0iDn7QGXOoiEdS
c9BXTBE7WFeaZDkmsFk9HVqm83SQTlELgPSL4s86vLowW3VvBQRbJBkyZ5T+KJ4WSiNxmI5QrMdm
Gp8RDXhkrA/nrShECxqu8/SHRnCczO+FHl7rvRQcrRu5JCgiC6PZ/ihjHFGxDLyIqxc0gnXed2v3
WuoWPxi6XOvMMRNXwhoPKIeVx0Qpf76wpQT+3I4sSRfBJ02FKbpAZBvXyIRHsckEOE8Rvhu6oS7S
BZYqINvov2Jc7BkomQsaTX64gru/oXidT+WHnFsXTCKqPca3Zh6Z8MfSjU7yamg2Hwgraakzw9IL
PTJ/tVk3VW/cC9fcMlMoHU28UAOdZq0jSEYlAh0S1f5oKlC+TlbdpuUG8TXE1x2YPWbO9GCXMqSp
FLlMTR4AtE8BTpRzjxIgxfPQNc6jqauUTX2JcwR1a6sEx9pQPYwdsXpn3AOW7aoz73Z3xJgh6L3s
zPwUYtdARlG2yXtlOhtQt7s7oA+wuXV5FJ8MyEhNHB9K1NcxJuHBEvpt31HiT85MucZNa0ZfCWOG
+1BZxP8dqMoGPI+M8KsWJrpfMTTIoJe7By56RuOVeQ2Ipg4EuNqeOYLM14/Jwm/wMg2cEoD71Tdh
4QBJlMeuKZALDB5cT5ybtwHJzhk1mR5/lTW40h4KfwwzJ0mq4T8kSz7EN4tAz9ixz+4W7Xc1r7Qv
LL/xIZtsOyRGromtS7PV2aLl/owXeb0FBx40vkihEZcMLglgonxBjO+pnbw43Skv0VzFzOxb1HbL
upjp3+W5InBSw6O575gYIQB3ZgYbTXGWpGJMGmZ6Rj58ayCrbiNGW26e/CwSjE7K+/hWlpC7FGhL
oxJoelFDwR+IJkMOCyAz2UE3KnZ66+w/T/NpuyuJmK78l9+fdoGw3YAx18WKtQz+IGM2cH5Xs0Mq
hOeX7cpSQQcCg+eBlKR7hFr3LjPh+Ewt8sQqq4/7zMvN30r+qL6NtQ2h4DMYM8AsepX1/6D4sj08
hn7bw1rZp8CUbV/2BGKGloBuOHwM6eG8ORFd53PNaQ65kXvPHbtbVOvauKDsD8s3jtV4OYWoeyAu
3zc1iUg/XH0SlNQKoe0kbZOCY4+qZqjmWAQrIFZcePTlrfYLsJOE2JwmZauUobYh+dch47JPYXko
Egj5QFwGqZS1lL58qBmfKwaem34yI7R/3A6jWj2yc0hxFtD1tBa3flTgHZGHmv8cxCtqPqSpFxMz
CaFAAU291KBPwmT3+bZ+BtKJ0MUTUU3LTwjQAolyfNmcLdXCHtMUcqSuiiAQ+Cc9FDfj6zCYUm4L
EV1hTyLYV2zrmDZ7RoY6Y9vM25LANzMP4nFAFEjBU/G5ZFlZnB6Am4WY9j/yCf3hSzokNnoxrlgP
+uwB/FeF7tU28hroaW04aL4Nn6nRuEOfsOAHFSZJwKXyAJWRutAfdDsdV52rmGpAQ3rjGdIlezUm
b+utxZhNSPA/IIl9iCYkR5n9eCk4Ri93MmoUI31S9m8g2Nj1lOC5ztvruzSfgtcZSvBnZdXgQrQ1
oxRWRUoD0xsQ9YwkD6+12geGNylhesnjUUzjp7Ocl18O4b1rP2uzNuyhh5tHr8zkgPauRtl+Jr7w
s2rJJtN4Y8fmMYKEmDmDauFR17PUPABkbP6nAcX9PTS4M8cE/fusb0b1iplHK2TP0jI5I+hfPqeD
D7j1CEF1uloDO2YxeZhh6o1B0yB++hD5rg/mndvqU15dpyZMtG0klTdZntYXM1GdLv320nQmq8qx
EbVl56BjxBWk/VRPVvXdVu2GFnkJ5l9mkUVmqcaNz8oa0VcN83BnuTleCmMsmLxogIBYmZCf3zta
QpWgP1B3uBs12EPV6ccWeaYVDcVvPkwTAAi6maXliyz+ze4y5POvpq76xD2QYYyY0Zy5IvBVFN71
QrTy98D/1SWH6Uc806Nlc2QhFyzHxk0JFJmD0JeCFtZx2N5iJG9p8xf0OoHKNV9ZDDSkjbOhkMD8
NMZ/UUkWdbkFt6RWGG47DamjpI8DCGHWHZMUZPLjD6YtBb4sBgdA6PE+Ouacy2HtaFA4aOE9X2wk
RJVN0YQ9pKk1aRFPFrttf/PfwgAHP8IF52QuZvOsGiu3r16+R1s4ElWoKMCA6MHaH717mS+NHBLy
OdRnIZHNHVeI1OGSJffR/R4i3aidr8n4U/YP6LFFka29uExXRKQ5RJ8nlV+zgWo9mnn1g60GdIS3
PLH4yLL6FaUNry9AYfH4wviIF9UN3Q8OhQ6Ej/mbeDOMlkSjV6JbJ5CWgP14nDQaO/AZYmKX5B12
yRuhWVKn/u335scc8qqAOcfYDITyr3yL59s283iaoypRMV7B8MzoR4T8iQOItiXtqsUfsHG2x1Uw
+n149+TcLnZXLYKAG1H4zR4j3k16BFb+KHry7U8xatl5xNNB6ZstmeiZ+Iuj1r8kSvy6MJTO5Cth
L6AZybbZBGzvvA4XGC6Wn1+VD4eWhmLZ2dMSy9RVujjlA1T2xGlwvf4KTKxCCpu6+UIVv1XeEcQg
gl6DRwHs+uUC/FfXgUVt0lz9jG2FdnYMTfixJVg1LKtWfSOeNw1FaBtVObB1FAHGj25jr+Va8zor
6CsZd6lwf4xexoNmvAtK3TVcki/sEuNge3y1Dm0hu/LY6qZAoR5a7hgxAtfuIqAHxfRQMsQQ4pdC
xz1lKYyk1vh9V4lYQDJBEHXHyIe9p70laTT5wbf75f1CYA3fbcKdXBTR5ybfsrsRtc+UN65racE9
z1+RNrjCAtcp9dHtsXETvOyvdrOVpJyHI8x50aq0ALVsBwolm9Of3/vwsQC5oJb5TZafQXdwqFTL
Xt3zEMYIFIESKhzkFQLkRcD92Pw2s7jixBHqXjgEVSyLHnujLCj2oC5euJ0brTB8diasdQIna0KW
U8c8fujoon4CQ26gvc7wqFq66wSCzGIxfzQ4TCVLBE1A7D2isLaXlfYHTiCwfdONsLsKbAaQicr/
La2LDkdGS2U0w3F7Pedngd1WA2lCtnHMicI3rqVAF+2VAYcjqKA7mVYhfea1ZSxz93qqS464OU/f
5BR2+aGvfGb7EOPktAtJbzstoqv+bGU4ABbIsqLC3yp0mRChi9r6LVTN+Q0mlTyAokbe9eWgoRSv
YkvQHTOJJ/P2HFdCjCu8jAeA3ifdbAe5CNdh6JeNdJOjcka2M0fJ3TNohb6MYfAIfHy3WNsZmZIe
LIBHKpcpyqXBJpz1T3BO+uozLtiWIerkcp2k7LXOXIUHVIaIV8prPYsxo1AwciaP/L4AGLQA1nMX
hmm/JKzx9WQK6dnHy2Z8SmeHIVLS4LUxIlDgopGkw076slcwW6BfxOiJ7ZMCkCE4O6omJ2/giA2X
DffSfVz7hxsK7uzvciVuKxtlKbizcHDc4eQOVoXXBQGihpIdl45Yvig3c9pF7NS0/DOTT70buzjx
svMBYEtzYBb02mGcOfDDZOPMCRxW3e6rwdNkNIEyk2ToXbUEop8A9+wlvrCF74Y2jKLJ5vwY1PT1
X5AoLi+2jdOs3Gcxo/K1apSkLLzQSFRtoUn2Al4MquscdrUK3JgcY2BULEqBeGJgeYVQiHxKnW3n
s+5LXf4AwjnwzWy+JCh3LDpsjOeO3/H7m359lU442MEf7+Uhpgi6wpd8+yPzet/Y5McSZPvS+lj7
rVB56pbA0vrx2kvTUBDMtDe07PoeYoFrSBaP/B7uqJtCjsWY528OYvC+/WVNreS0lS8pwzPF9BUP
6D7W9YRCVVGMLa+kSxSmx64nhJXc5CVqxL4siGQnIO9TWDH4P7bGDX8mg54l0M0ozEH0zlbl3HXv
ErP6uAHmTUaWhtoORbZ2HqUxmIjDgqLDUD2O/4OBy1SGFZS4nK0tjCe2jj87Up6a5T80G8go/auO
Qm5yQoBertKsbMfasisXiAbU4SJxS53kuYAkh+JF//FCko1hB919oBA5f4HVSfB6PppY92TcMBSZ
fGtnsK7pzjy6PotVpKIe86ImURDcoBTAgTWJymyEHhDRPP0BinBQhRpproX8kKTE3hye8VpwFSZG
Id2DKzVnM9hYbytwAKbP4E36sR1LA/M1Sd/brToKeORIRxdEr2+4hYcWV9PLav7pnewmMKG+uuc9
6Ay0zWePdgBMHh0uELJQS0tdb4ZaQgg4q//mBbixehw3Un+AsoAZ5c7j1XS3UphnXY3/PIxViegY
TwkZd7DRms9MBXJQi0iD49QIlfuwCqrShxXl57zDCncQ4LP6Oiyslm4SanhUGcMthlNM09ZoPP4x
hWcH1YXOXu4K3vr3uf2gCwBrLiahaX3e25e3n5y2FL7TaTcAkolj9yw2V035/zAtU/UeGVf5KuxG
LhWbGaKYWSEBCWWCJMlu3P08cSkAIHsnysK7wuct/dwCQ5SQb9Fmcg5FN0ClQlULSNgpgPoc4G2v
vEC46dKpnJVBpnjobYxjwNoCYMrMj8WtlZHGIyJK6Kmnk2gJIJOBawgikCPm+O0T2dSX6sWzFZT5
KoFaQyQTsxh1RSL6ZE8LmgaqMA0ZVT5SvEdciuyV3bPnY3kHIsgJbG1bXDSPH05NmCJGBNT0RXki
wCc9IUz5P3cLm0ohzBhRLyy5CuXzUhh0BKuoJ/dmpRjo7gG7JbvcxYa9dsIXgKSZFca+XiYdlp53
JT9Ur+jd2eco/WzbtryTDuZ9Nh3hkPng3v2Jz1odFEpRJVayKpxCoW+o7/BJZ38PHuxOQSaFotGq
KuhdpM2nOur6jPwGclvCWs/6IhDOZ/6O1CQRCXsfnh/0l5WLAfNAXM68f6GWXLdi7mitMEHgsstQ
fHh06k+uYOxBeyPuPihp82TtDqG+n7dZiicv5H7l8GDzxWonYevTd3kFdirNFHX7fU20hoJwiahN
OHo/uvdFnOEgwzjtj3Zwq8edtXTD0VfC0SnofrJQPh1w7IeR2Alq5vvXwzG40Rcf3s0zSzHT5Y6X
huS7XT7zt5wPQtimHxSYRDwa4HVwRPoUfxqkR8PVxa0sIvoJGQSzsohOe4LwP48r+f7jrXptMqEy
5FXPz8ESKekUUD+G78iMOb8nkwsRg99MXVsJWN7f3BxgPfAaAXuHQ61KW1IOWadHLwBpPm5ESIqJ
gSWlH6jhXWsTS67xubKyZ4cyBeS6gz4hrtoWSLnBhgJP5LGk4HBF7fNp9xfQ9K2akAUFiNHrSpLP
A0pNPLx8sfwfOKfoXJyl1Yeg3C7+cN5nuZgCBK73kPMWA5I3dLhUq09BKkPSgk9zOc5L/pOjo5Ar
C9UUihPyyDiTF2cgYRCbGwRnrf22c9X0hEFKYk4bWbeRjbI3WCWo2TePOfrhFAbp3ZWTZKys5FfT
8FM58ICxFijZIYAErvINltrdg08LKg89KmpdfNzpFk4qvppQA71NxhI4bZm1XNb6UAFZKoPpALX4
cEdfE24b9HL7EsLKiWytJCCi+1OTCvL/AcUDoK8AqDyctqM7eo5KRE7ovKy0Q2/xSbl6QEhmLcd+
SSW3ZbkLpFCbBu/WPtS/eVeeRW6m6rq46I4oCSuPRzfpO4H0xs5rqHSIoZgms2A/h6JdfSu7d63i
OWut1SjalsT7cR9jLDFBwJMl3YB3u/MYsxM3SdF1ZDmNP8y6guKSsOv1sK7GgYJPnvlBaW2tUi7m
M3QRsLYDABx9+7/D95viofTHOXh3ZoYFGyhVCpxZTEUPx33SWxESNiKKfDwD3RGFhmlwa67bgp91
xua0YuxPrD1BnaT+jPlQw3ok/tdUhwytRO5CrRljLrzZBff9k/aRjVOrYCxto1lUNlMR+LhvjIaB
z8owS9+0NNHEhviFCmUZOjaC8RhMddTPRdmN8aKT9dw4m951vQz+XDSsuyOOEAWCyFeijKq2lBC+
9BDPnfXaUvl2YhyIZEdoFa9t6NOze0H1Yn4Dx9vg8Vq4NEy79EDeJ+icCH4avhfjj26hxEa3jI+H
8vpfkJBruSFEBazP8+JbM14uZcPutGdWybV+CTsgYxDqNIzjGhOthLLMBM55bNvUtk9GPk9G3qfp
ALLdIhhgwlusVNSbTr9cnNGTViy1Y7gIy8x7F187gX5/mVbh9rB79IEyevmZpuqGtY4giYa30bcB
C7Gp57TuXyjUMiatbD2KANoAsQeXbgZScgIOX81XS7fJr2Re8sfHOQQt7xGPNwXb35jWPwDbrF6C
YwzKvZJNKgShg/lTI6xr1euOFmafdsEC+1uH3Q2US1kL2V/UblhDKLwF3spS63YbSrZcUPxj6Uvr
5BvsvtvljgQ25y7/4dO1pw2LhO5wYeLD6765U2bNGnkfyZHklOWbb8uofzempruYJX6ikvMhGRMM
AW2PCMk10I4ZlaXLZUISq0kQxAjR93fdl0Uhagkkq/ss0IgLay3jotZKHBHEZZLVRJycR+wGB62i
DrJdM/uY0kaGbMZn+OcWL0NPsiL5LZRbH45n0hNHIYCxRZdcJcmfaMaTj06swNO7oIRZXfnjZMdh
7iVhVlX3/3x6+xB2kjRQUBihcQyMQMD2hWrOPeX6NjkQh1S8C+ECdBRflVvIeKec7YcDvzovQd9x
fmdD2SlK6ZcRQHw7tnYaTxGfwwxpUQLElyLToo6RrWVHe3w/CzBuTr6/OBro/pHn6AZisLntBkxR
Qou8Z3IBNtZ4+wnBQd45ULiVq99SjO/C90beluT7J0TaimKohX/tIT1MAbkWKwaI8d3xaAT1s5GQ
ffpXZS3y+yjPB8ET8PU01fr2R+IYsaPwkqHGDs9YbpbeF8arj7jkpTUajEa4dqGRWkb01Ooopb50
C1kaiGrh4AcYLv2EWBHto8TkgbHROQtNBz0S2XPWE2jSeNQIAKHdkNYCPOBmd7BctoP9KF5lSHI/
6LthRHuI3ueoEF9NmL6eiBGshMlIFsko67wppbwUd1weWyq2IRWEtkUGcQRXwtTXTK/UzxRvQgVC
zdBFc48QVCYIPeYM9MQdmaZgxCjNrOgqEVtyJGR5+IP5edFCme9YPe9cfQ+VUddm+mMkpSYVRcZr
4+LDTLkSAIBYl8WYasvc0qGZLCc80/w+NJBiczOlJ7VzI+jN1Ogh/1s/NaRkyL0aZAdPF3PYtIjj
GvGLqGXs/j9d3HU2ctj39dk5YLLwK1bNW0eQgznZnJAYYEo/SRcyqRkote0vUQN5r9PVlhihJPDa
l5gi1a2OpuPZtlr9WmLAWqzaSawnYL/7//7zyY/WWGP9WZ42qEWuqibYELMs1vibQXVq9p6pJ+Zk
qRNSfFSTCuDR1WX9mfn/pT38j52CUZcwHIiUWxHzAF/TLGfCtci04zenes7ZPb0TTqpuKlT3I9nr
LaMFX3JNXHwp4hTsV+kxn+llBC+UogRhm8c7fRkBj9nXTXdKVzKTgorWDJmJ6itX0LzH3lMf5yAp
mftiLgg9onux4YI9ZXK3HzMDYJ2L6urbldzPHD0P57h3JnIV+cgohe5zskDCiM+Fwh1S9EU5wmQu
hT95HGlS3sAwNtycoVfDuTOuqDT95g5SVHSpJJwz95BmKjMiGrZkmXNPQsB07OS7+NywlKJxcVZb
/Gs2dUP51bWDzipNhgFLq2Ewma0VldGMEvHll70NS0xN8sCrwwo1f5T/x6Kq3UOzx9dW+DManr+O
dYAxz2cLrf/Tv1ne05kYP8i8fH9VyrdM2uEcRu2G+IwFvXFWcfScsVuLBWnFohG7JqfF9TjMJ4nw
vOcxS829szHH9w/n9RsXCpEEu+yhAJePSGenVI5WgBndfj1dIvMsgvB2Qi9imjMLQC+bC2jCSvix
4+z+VitqGQqMvvewM6EAl2yi2VBo/uh2Rl85ytZDSV4ghomQLGueoZeuRx47gty8cL0/m0yI10GB
A5cCYSYMQINOPVmDbtICTrPMiO6XxAPhbyni28Wx3lL9N1GsJu1N6n/95Koq4PXkwcxpQ2/jowCl
jzN03ZVIHJm07pElTKfUxRJhkphO/JQ7e+tmAorYUilLi0SYEbR1dH53ZwWMTqbaYMT6tcbjU1iI
9WVZ2qo0hQkzZXA95U+9cAmRcbV51Ay9hl1gqB9L0vhIxVniUBRxZuylp8uXbIRCwnWs26FaKDiy
n5JCK0NolRyktIqCerxz7ukm/8XSgB3apW/hGHOIGkBZG53awnX3fwTGz8Ds+9VZsRczlB3noZMO
JTC1eR6OAF5mnFLhzVXLLeLqNYEe77iT+nXcl2MbgO715txDyme6KhKHlLirUEia2gpPjhjd8mYo
OcRuA9gKc9BPMgM3zXGP6zPyBkfJxcjVwvanTLpGsbPmc2i0FqVXoWiC7lj85lL3E1ffSC4wFpXL
FL2G5kOp7rhYUTTxQo1GBlzNsT1D0lNWqpsCZCozPLV162C2vDRExGtIA2yS4+msfu805Dfplb7s
oe+o+nJOr+cpJ9y+ToP0a5AlaSFjFFA/7zDhhMRWT85+sYAs2LjT5YJrRZL1Y1UJ7X2JKtqk4eAm
UyMooUUAGf0iwRrayjaGMBScUkeNgEAIpRQM0RqyseCn8Wb0Syc7Tpw+HgGBGx7o8zX3dQE2Gmxa
nAN67QgGNRmNEsHEzZ99Bdyr+04rlOkLemRXn1VMvY4LylTTGdnC0h+b9rltNk3DQm9pJTdRlp8r
4DClurzJHqOTRS77k00nh5h0t8IxRR3COn6r2lLnGVz1IyQEJYSf45471iWSNSp8cJBbtFnNwfvj
U8yjJ+B9m2YtE3zExyTEF/r0gjZnYVIQlVwzdJ+RtHjdeZalymcaxmv7jzUy6a/jtA3t0S2LMBMG
Efpbg/fUfJ79p3vfy6Pb21tAc0sJQcvHmTDIdGWVo5WguOkkcTQRN9d0sKOvEDBe+xgqRp9Rxd22
glutEmQ/e7TPTX34hbaamgqc2QDeHbW5h7ArhegFrSIbT6a2lrosOxbfTd17LtTYyBzK5jO/tEmB
taMgLA/BSR0KZsiE1jqpd2kcqFSRCG3ZyArqsq9r3At6YZK3vvUtsfEnwBZCY9awQR98lw0u+K/a
G+xCSCmFFpEWxCw5jzGBcKTZV1fieFPBi9Hmi81cPVHCJzUVFhgaejiuKe4O0B+dBDU4XZ3IxTjA
KMB51A1NvqIBC93g8VggZbR5vCGRGNIouL/DUmo/kVWMdeChjoeS9rWzBWrw1jT05crcjC9dIY9v
lNIdwJtXEuin/TIbU27zihLCQoAD1D7w0R6DeAaLe+VYOUe7xoa7hhE0kQirPXo+UcvaF+0qNum6
3wms+RUjBCUAJxrqYnNta7Uj5ZGENhUnvW5ZO/+2ekBVIhYtoZLaD/exQUYWDAItTWna8riAHnE5
yORJvGr4I6WC5vY7OI+zNQyHPm1+er/z6YbyCICq5XsDDZOM72QKGUsPLhsELt5RpoFqakcJp4Q+
Bl4LxKELdvlhX5Itjx0wIlHCUg1EZxdQtRIJ053BIV6VmKIlscxV+/nnzoHi/vwB51yviw1Vj2rv
E55jxNZanqut0T3b5Pvb8ljapc+Vx+T9OEfGw0tqBE6Jb4g1ptlFLgsgFN0gs6u5iOKlrFmB921m
XNq1xXze44ZYb51HCFRudFEBrSYo5GznDPWQGTebDg1upc1+PElGlbvXMtwZsuH1uMryoWNdC8Mc
6TzGdni2Rht9iIWy58IMl6cFaVcoZoTXS1VIIZVGrc749EjH6zkoZzh+dPmLM90bv/yPCJgO5X7c
CoHZFEsNTYcO2XcsUctpSLHt5VlSwUbmQ/dj+2CuOQldPHwNy6SrS46PxyVqsWk9DVVojV/0cEWv
CG3dL3uTt02fvydhYnwLzxPwYurxy3kv9crzSXkCdKzRJTeNMtbsIaiM0vLVcQNifngDl2OQwS4s
VwQeBB6uzSuBf5F1xBYV+NJqEbEljLeztP4ZYmjAA+AjlfYCDxXgoL4PEzz0DY5qU3v4AbieS3Y4
TP7QTaHpX93Uj6vtFANZKbmcdEHGQCRgywiQE5+otz4KBvUi0XhGNkFS4q088HX1XF0jKkcaXWQO
y4buHD9/d8Q59MESI0iv1glqn9rdnDZI18MUPmZuxFCfgT9wjAsHj4xZ6BA58eU5QSPt0iknZLOV
eOD26bOL7RetUP6xMOD+TdASQLltcCsk4FsxvoBmp0x+YJLBkb8amPz2F/BvZuvijMV5GgAGY3ZD
uW8YRQuzykbKKlOflmkwA85zJCzuax/5Vtm7s561e7dnHLKzVkUbozOvmcFb6w7QOf6HOCMcNxNa
Oh0Qt/AvwvaBw1dJm73B8GfrUoGaS+qmVAmLv212/AeXU+rXPkUWOd+EBfm/ZY820aZ1ZVddaeKe
ovH7prKMY+t96yh8+PDCbih4gv1ZtY/oBrAlg/JRh3IP5ALiT+b9u8vY1+2eXeimHlyhNnpA5sJF
sD9oZJ89vnypFd8CFgaQuEJk2VvufM+84og/pzbahtvg0EqgP9ZFOH9E48C7F1hnkWnkWdvEbzr1
edtwr7P2YWyYm7qDesS5SiseHYqQlqbWj5a+hsahoA/8MryiNG74uD4Papc/CUNS4hVuy0IWmAMQ
1RUT2OO+CSdNteJUR5/URs5cf9cTEnDDnalnYqwS9CcM9I2v2/UKMNyiEyQt8WxYNfCtvhaVglpu
I81D94lcvT3cIVXsnOxor6PHPK92Hsu2ZLw4mnRoBfLWbfpQLg16NmrByKayZPU1K3JRbWYJwyKt
92KxMyjYiaApNnskVd/M+yaNN8i8+Df01BrVwj2Nzjh9R6pBrap3IVloEeKDG5Ftcb2/i/8NVQ6z
QGddb+hUQhjqaXIyGjc8m6cqUPrWBC54C1w70uvdPr6ZmOOO+yDerwP6ih6bSJwTXYxRqIjFS4DH
P1Gtt0seoYgQy17bMtjra+ZHlWgPmtc4CHLOHhmRLi4cbHmDQEN+7+sFLxD3BEL1dZexTqKG+bjt
7ssAQYNd4H0jKye536/f6378V0Ul/ZAXKto5aYrWmXrAubZ8+H0RnRYAkvTKpa16ot9fJJZzb5jK
RjNJ/xEWW5q8UXc988i8AQPtcII4Gr6y5SW2xirX8iUUididVYSBSudRT1iW4ONQDHkokJsSHS1I
viXqdHuULcDVSUTOzB/igh5QUULBSVpJbj4ioiHEJD7qtsS5W7aBD00FE9HSnafLbnVgD45eDW//
hPuyYIU91ErwTrSZC0QcETVqhaK2hINwej/Sj1176M2JNURWw/dlPqyBfsUlkXz43IZZlpg0qaLZ
6CTAPDSuZUoLQ//zjiRyh91erfPXzx8IIg3C84VWs0ZTXrux0ZE7Xyudk4bxstWZGbGI85gDZawg
mCQKPD3fsRCoR+aXqZWdjGAneMtzHpjOIZJcFjloBKtMTK+mpMoptVCiuPYAyJ43Jiwu/ZxQv0CB
I960eOGwIeTbTGiBvDcjjMZxOx2bC2coOKHJoBvgXkOOk4Kye6eXEbNADTBCNi4ZzGEdlMYUHmju
5+B/jIIAOlUoVi4yTR70qM0g4zOkPhuBV6OtXzamOArqYRex1VKF4Z6jSoiaD/lJmA4O7UWFm47e
3TWhPYDxnyz1iwTPljuA9MV2J8bcDw2JUgv7rMKyZU34G5e5OeVZx0Acs9VIj8O32p+Y86119vel
hQpKCT2XN5q1Y+1wtbNYAHaKk7zEFzWsWnRy393z+FXKhGxMNcvMd+KhstVzJbTPY0UmJSnaS057
pP6Sh2dIw9KIdZVuvNaHuN+ua5qdoB/IREXnKK2/XbZHVo20IxYkYKvW+xMLnXtIKv0eklwdSIKe
Or9JrZAB/GhD5fCJn1C+YSXfjv/ijKHAPjj6wG4yCtIvybRvbaqiWgNgKKd8gRZMctBWkeUWyAnz
5udhkJALFfgqXmdvC0w9lAi4CzZhcov+nVkudOFjKcOnuj9kWtbZwCh39MIcJDw05FyRN4BFGNQA
USIQWO+/DSncM6F5mLuTwAE58MZMHR/OnvYgBZEYAVHPPUGq9TisVwQlNNbaH03evGTAWUSdgkRP
Y5yXtt5dq9D3v1ltjEEiHUDhluGFx9duWehqPTVf2heXUtTbPGLqHBxH4LS1C1Rk0RkO+9PG9JAN
x53mTiOOXcPtwbAO/YUI2AGt9A3iCRsTskybNJEEsBAfEJiA0zTOeFIiFEflx8DUrN2K8s72N+yW
0+MAzBQyFFyzYkomG3UjhO1y+gbaco/PRhtsmjUivpoZ+8QHc9EusCrbRTsgcYrDvQlgMXX3eJoL
blCiBzTTAhEvdpzdHuWhKZLFXJPZg78sLI2Hpf++AmyssJ3GiqyRrFs+3T8zb7QAQ9Ulu6DgOSfe
1ia3x3OTVSpid2lriBanUms2m6Qx1Yo2WRm47xIOvOdf70WAR01fIZXVKiZ0lhlVZTlrLjLUc8WP
7+ydJzvAfjf3nFEOzpOZ1r84JHU97g3BhxBnJWNCU2Uy6cDHAjvMK+FWWUQ8HWHKuTByfj9ZTXFH
2b7Vm6FBB0kUA8E5IC4le536/0dBstQCYdcLvhsyqpkHCa4JBIeS4KFYYjQpFdPfdayj+ruf+w0f
t5dhnBk8GiQ9beY9t6x3GsGbYzE3z/AJd+/O+HteeGCHOL3uF44axF8nMFCR9PmRSgVSA4cqG7O5
JwVh/2WB10Ojul3Aef8i/7FfRZDduClQZcr7c+kM/hiwGJcNfSm93C/DFD/t9Ltf2SdcmOoB2B0m
4iKavfvVnRsSmWtgjTF11P+YpN39lSm4J+U9Hl8FwHR18kxukS/OGxLnFkKf/tEeeioJapXkRNHU
G1+bBzj0R2JBDufMPXrfVxYsCfFzjIisUPTlAbR3z9Qezs/dwjLK+itCuroM/20ipj4kuHGt04Of
8wO6h89cTWnao4QJWM0QTBUXfsT+tpPzAIUrm5rc/WdCdAmq7z/wV8D3YGbNH7C700UkIeA/F4Ec
s3abW+ouaKbwq9/Zwy4Xw01TuMRU0FVc6zVoTPjR9wlopIgVzHA02rU9FL2GfDq3h/aqUETvj7BY
hT4CuqRyTKcWwxa7tLq0IDxCIt/JxCAD/BJHKyvdfQc6JlrGG/jOcXzKC9wylBzNuJ/E6Y/aZRuP
BynGmwQncQ6ITZBi8k5i3pijR20V84iLS32JHTvKaXOAa/Pd5JDwBOgm5a7Rob+3K65iwm4zWcVw
rFu+uSp8LZSR6GSaOWXwTbK8XHPXEcNYyDHbvu+pH/J37m7FU1owsqW/mTXQO1ObPgCW1H+deECf
dimdxjFa4oLYb951G9Vb8C7J3Pdo6uEmLZTLqb/s4qioQVDRfUEc/4nGYJaEU6PrOjyFk7+w+bGq
87hTy/KvtR8zRTx1V2+OWqtfoUMoqbzZAONz+/yp1rgr126TXZPrkwhKRyXn21bFmsB2aGcrSrFj
xmYmjOiX3tBQ4H+3BNdlTmXIEfxQOH//KVif1jmF857jcZIvIi+qqSGDnjt1v2CW9n8SbrOIYZjf
zfFLsYy5ZwowYl1jpEte8iSchRLCMwYU88iBKLlv1w5TfdCmzQc6z0SqetBP5G3XJ6X2qylkWnQP
/Y1zJ8QA7r8FxSuZKfP89a9nD5hisgdbwLWVpXEr7Iz4J02NPDQtCwn0eN9msXxJUo/ruIY0FbWZ
nZXlbaGg/QMEbj4cnwTyKoDK7USRH1SH1NGlGZn3u6YYchR9kAy9/X6HMsdZMrJsXsTeSqKxbJzU
F4As+iDuBGAFHnyrbXx9smZBZH0H2G3MSVPKcfx7+THq00XNLNgQ8MsSyKH5u+fEj0vAYbpvY0Xg
4oQye8xFOPflXloeCqFJqKuKYGMP96dnoNdIdTJ9fM5osnLLwIOkfar4NBZMROdbDJO5VGsoI2VA
rBEALnfDbpg4Fs8Xbita0GMawcWOMuTajmFIHACJnG/cxBseqeEEVmIxlBwCTw50GUzQBybpKGYi
WbbR7F5HsbICUGCeHwevKfn9kQTLL/hESOqDGQqgV4I6RKJvoVxCIxKWhwxgo34MEHBhzCNOTmU5
kEK5fNcOOaxtojuKrLVSfWWBCsgJ8JAew10A6fo+85/VSz61TpyKhmeMvnhQkcpUeSTBQ42rXyek
ZFDqWK5DYcV8jy17bKzASP68/XuBKV3OKEK4vp3kb49whoOCk4U64BtPDn9TpeMUZp5OwgOQV7hJ
3UBaeHbS622h9Ea3MVF2e6EBrLdIfuHCQZarCj+wgQCheQB7wwYeCgk89bF3nezA7K5VNOhVqMKk
+JiM7jRsaTKLTKgfL0Z58WQWH3oqcfu0/3LRLqmvOA6+gPjzfJnP9pBOtrNwgvaXYvnsBbzC8Tss
vbU+ZQFIh4pIp58qW8rk9W/yToFOeXc4Fa9MNfPFtuv1+wo8aCVAvmle+2lxqR7XGyqFlFC0U/wP
ZxR3sJ990SDgrr8Su4mDFeMxRwPTP2h66brrEStWLPu6/juKK45EVg+8vH7iJuJbIFw5Kdat9stJ
JFJA2V6OTiOaDec6Ucx/7rgmhghZI+q8+ECy1J9sm4ID/mxGYcoQzFrpFa+IjHcZ/tkSwrNEJKIt
U17nCq+NyHv5MhDqtMkiiwt50Wa1kwMFma1RVGrs1/Qt1gV3GtnaSwFx3Q/o2eqJHQQ/hVayMY5b
qJ4h8uoZllYO0qWIqXCt+d8Y01FMiaL7TjsRbaItzCYGXqWXhyauwmKPkYFNJCAOHx0l8dDRbFYR
h5biRNYpgO3IrOKVKZYs3NT3KXsYeUuZC3zLKeNXy2IUbmEZxSdGat3d13/2eQpDYG0FcnSzwflu
+bJ2ZUpp+gDOzB3a5MzytxTar9I4DV8tWu9MEmKRFoTpSoJjDVaomfSD/6VA6W8k6EM5BaWn4jg2
yTKjmVfNS68hsJtFPzPCpxvELC7Hp2bqqREHTX8wD1RNUGmeqPn6U3R/aBCWQyVoRU3PDC7QFfqA
/KMEd9wJ8lj+UoJPAX94QPLHk36M7zqEn0ds8OakZgE1cFD2snStw9vm7BF1WnfWoVylozYT+bRV
3R5ProzbMq/lNcSdqAGTy+9yRS4crjDWji1oNJzSsEZDaXSHV/wirFgCqrvSpGGcXgE2WdUixJTJ
L+m1Mvy1VYxAT2cnlu6wOMPBPGSD9aHOQYGb67YalGkeigl53ajV3u4p2WP/0WT0Sym83KwHfVli
4nsSXNCicQzy8HsFtZj71i/OAwRNypcA2KqKMTlSTrBABNN3sAybl4jLys3DFCubGHMFkKiwvfMJ
I475jI1dgI2u6sEOZQbIT4DunWC5Ha++NwlkaqH2bZtXv+ACQrFB/s0iEsNbnDOAhEDmuJy9BmfZ
wnutrRzRk8DhlVYAj47d7ZdwK9xvuyJsd+7QVo2XXJKU5oDwR2VLDVhdaZzF3mB+efrKRFAL/bTG
7LxckrWwmfLuLyVk9T3WRqnSnLvwChOUgMRl0P3g6sIFb0FuJ+Pa77CBxcP+CKQMqBg+gZYr3UBI
IPVOvgFeEOoLVMSpEIGVUq579ZPDML7peYP89tWth4a1FAqyFx/Cgucnu9qzdMqQo+hWSpphV8Tr
5xgF4G4sU2lvMSW5nBZwqLPaJDthRkzE14LNx6T/X+9oWQGupPjyWhmveHVmTUWjGTf6phfUZoV2
6W+PWqf124V0FPbU6UissgaGXMkkXMSL8cVNY+6LyukSj4OlGmXHCRHuUFU+m89kxIEYptuHJO2P
WSUpFeiLFJo6D6r8U9vSYVHxwaBaPsfTp2hJI3d3/L1BHHvLwI/7q25HQWAh5vHnFbGFlyL5PJhO
MbGIPsC+reebUB/2rFlwGNipQOOp2oaQ8gtmS9NI++q8ZmEcgVxB3zchraHEVjMSqDfvTYl0c/oE
z/UJMarhdbg6NlBcCvgYUXdCTnfVLElDfy9rskecRZ/W1elvU0YQY7Z1+wnH7k+Q4jUyQWrSX7Ah
GnQfprZHry/6MR4A2bxqYTwgj4PeD7C5f5SJqbR9IJy6UYy6xrKygAi/XD9eDCmilQB7G86ieK3b
7q6QhADirK9JSy4VrfaPJEyMfwjq+Fdau4oJ/44mzl46wbItZQR8mn3sWUEThbEflEqqFX/X6PvX
zn1Tal5t8e0dQxc2RaaapnxZTrbFsIszgamxYyIVhbw0gc32nGeE9vAbsVl+Ppli9Ms6UhF+Wncv
YphIrYmGljGqiYwxsy7vjJGV0o/JmQ8BNblu/sd5+Mh7ly1XvEfQar/+x4HxvVTI/iQMfzaXr1a7
zfTg+ypiU69qJYLyauy8TWEJBzjKbvmHm0E8cJslSTuEr2UGbOreUXF9Y++c1klSn4ncvENh/cIZ
jXlA+mYJI6IiR3AAEIN5fX4USRSRgvq/D7eVlMFJev6YrzriH9kMion1o2g4nFnYVgnrpW1nw1Zu
DRsscnRbI6cKc6soNAykDvnSfg4uk5/DwGEcc4A6tMnaRuM7vL32BUPoZoAwD2QwJHibRO2k2vca
LdF6NlFsuap0+HRUaWdOW6vjh3r0hRFV21rUb6UWO15kLuZEXEDf3EY97BxWUbT0yfJaTgB4byuC
ZDwQREaZFrhq0TWsEQ4BoG9A8S/CBfTTlftowKN0T1/0pY0xY7O8DMkfmb3EGK2H9Ed8AYdkqiGa
FmvCxuZUB/a+87hZ7O2ujNPCYEdksKbp+SXvucutliM20qLwlHJjKyaEZ+9Znn4yMWsyJ3thoP4Q
IVDgxmRsNZNgftBerFGK2jUNybF7uqyhUoq3g277MgZc55k1AVv8o3jbs/IENLvZEDQo7Np5REbN
31cNIssPT/+f+JmS/7u1mjejVuoecZelBoLCND4HSNoyTTZGkrG7DAl2w4qA2F8b6q71PlH2SWVX
HBGkwSqNIVue7/x+z6T5qESrqVxlmfdB1exbBOGqpc2iCcD7f3F0z5XjoLsAuZJB7+3s1J511+rv
BF70xBOR8PFeAd6Z2ZN1ppdyLsTqhHNp7Y+sAK8a1j/7lu4+1wW3jQghyV2FTz6YftHXN8iYkEuj
7R24BcljhNmYqcNRkeziidVKphDno46HyawG2EmAEih4f9aSwfzcARsRhMxxMwNCuM/6JN2sEhlm
JCn8ZKjv3/EqBfZSy4ZLLgDdrrcTKevFXeC5SI5hqwv6zYyVqXwiwzYQVxrVwMVwlDX2Va7/NL+m
F61P9NL+qxBxrxIi1t2xGaLyzHF5DQo/Y9Jua0kgJ4muLPv/21YtLVFr0iGTZfcVtj7kEIjPJdOL
3czuiQB1Dojh+0wHa5aumZKlNSHFnokw6JAPb2ID/yNhli9dCXY843o7TTYpjN1uhnf4OK3XZj3V
lPMhazm0fSTUelIikIoZld6fneXXE0pwspnOhqtSn3W4Xft5BT5/n0mJlAvBGpf1emvlzxi0Yae8
NGT1EPXanuzq1LShLQOm4exLch46Ozp92OrRRuQTKoZb9OOM0Oyax9vsMoUy0Sq3sb7BJxFXk9bJ
4WREr4q3TMs8rDntd18Kg93FGuOmV6rVN20PLI3JBDAmW7dqq/Taln964w9ZQezC+vvm1oE1qrkt
uzGb8RHpWLu5BS2TLYEHcTGEhUsLM+/3Ayv8jlOUl20vc6kBG5QILzCJ2BAAIFHZ1RQ2Y/2yf7qD
w73kk4iamDp3ErHltNVxvMHmkZ0sW5/CYcor+zVBvPCETMdBFphdX4dIPiL82THbSb123xxY5yuu
N9BeoQHJDLLhzOxS4RDRuC4wI0qhaUwrLf0odjxyAujCwZudZCulfYGChBL6yCqBVNKRasCCvnKb
oVpThO9kOi5vkfNXhNlhrKGYNHN8rYlfXZ4KJqRpLrncSIe11Ht+dLK9X/yAU4DkCMDgEUNYSb3+
EkL9qxY9Z8sWvkUiFvPHb328zPEdrPQwTaSzQ5exg5SmJKoGNaF++3KwVd8d3TpbbG8xN5bag8lm
gMuzxjivIRD7llywAxo0rUX9inKfHRYbdyIgYgpzXmWxOCY13rtNHftmVLQB5ZZsxFxMRE5QqDIS
DwKhq20EUkCX+rA/Uv0bRej5hf+32YGB+M+MTo/K/QlOi4ow1MNdHjM+pYjGQA8aE/rEfP1QLqkR
5DYL6G0eca8L2FN32yjMLeERgBjAfEBALIa+J3tE1egnDDtYryQAU7e9NzaIcZ1Go0uZKWS5wKZG
xW79I9tO34qPqMuaayV83YDd49qnpqCbav+muwV5mE1r7pZfITww+u0doqKXl101sHVNV8lKW/59
9aBRJzvRHwt3Bh1g2eg3KrRv4Z72E5AaPcBB191XKMGkVPBe9hjnAbqjkvsdMNsR0x5+IWvYjDed
9rBQO2uX3GIX/L8lLtDgZImLRGfv2F+I9+b5PTP5o7V4NvJct6XA7MuZdZ45GnhcYjYPLMgvqNML
slEbpLXaOyeGq8tjK0Pqcj2FZ1TEmpF1QgMPaKDmdGuaHDXgOp49cCgyljvr9jQLGTrBxsI0YMzs
g46TBLBV+W15Kb/ssuvD3CCP9jjdyrST0MLXmWmgNvKogqrjbj4bmUti0vfoUOfPfwkHpG6HLLr/
na1DhRDUmjYNXzSwRbqJPQ6Lgd/6bToXfmvmx3jnnJY/q4kAdAAB+HkNmc72MPRL1nZ6vSPgeXjX
38D3zQrgZMkxwzgyVTwTrq872kzo6qHrjXA/vy/VliV3gcqZbbqB1mbnGPLrl+ixOxJjj8HdnOYd
JoL5dGYHLhzXckkY2SIwO6TBL3tG4HzQbKfVCJNaWcqyodD+TNxx0b+Xj35ujdnMDHN2yZhvtVxE
AsNm+kKm9n750HI+TDel3LSpG54Tu+TCSiwuzW4P4otWgVkAYAE+JmWlccX7I+iAcRdfGHD6Qz5B
Y3l/0XYiruVsjzfP25ZLdyIQd5xkhJCi5x4fTubNUx4qu6Fx2edgaMc1f3ojLI7F+FM3ZBuiIkkF
C/AIyokRVOBXuCfNrL+zqz7Rb4aGKPZX85wVHWGvCzkuOYw4cRqxiE3dKtmQy8AkbrLhc5NnAOQU
V3XtV4cDgp8YkXUlgR3OtJ6JKfJ/auNIGkd9Lg8vIoAwbRFJHc9GziPeRdtTbtUk4yTFCCTXvgEq
LPKPBBXL9JSPuDjUymOH0geBkkTbiqQXB3Wl6DGjzmsABIZVu7HOl4Miw+ld2G/iIrtIIBSvnGoI
Tgf+V1nzJvIiHmKttndHbAgQvnLkQMkQAQ5mBtXf9yLItnnC72K2ydwxOtdqOLSASR+u6QkFua/u
zBXdp0ojSuBE7GS5y9lGkb00b1X3jpt+cXRbL6S9hk0xkeaJscbTYsaaZoaMLxJxSvUlrCKJ7Nlq
OHV8At2h/h+TPcIdyy41i0zKdq0EYHrEjWLPHbiIVugYg2FbLwcBFC55G3Grb+NZgMufAHVDEqpL
lHK1rFoKjCvj+l80AbodruSO4Z2H0hWM53mXZX3BSV9FMcweBrFgcfpKLEQii2zTk2lenVu6XKt+
nJxyQGw4Jfiv8+3LU4OHJED+cLlBfXnehVQhqvRiyL0CDGGz8aCt+mlAtfrliN7yLtLm32FbNlo5
5O7zJr7bKq22V9LxKzmIZoB3TTQEDeUERpzAJDz3/rYa3gE7zyCssmsaNrM802Tmfntb3/1LdbP4
ZA0+XAcVr/EqhCMzRrhiM/r2JHMn7wrQQ3KMvA9HOgn0qP3foEq2GFSwJ8ibdXBYtsfhUKN8x8+7
Y6Jp3RElbmOTDS0+4EbxRvKbbJGcUg2ytyHIIaUvH1z8rUNzZfeApWcu8OqycAKIypwDNrcAqgEu
VYY/DoOJTUEWzPnIyzWeswWISLBaQ9L0Q9cVq6RTzmPaMSDNaW8Cc/Wip/7jpZC1ai48e6MHteB8
BA6Qud7Y6+qp+EkjkpuNiLeY2y4PBHiroyei8UBja9gFK7i7/FxmxC9r1AmXYOHyiBNASgdPrkJW
X0nYqW+O0XwK96vejVz9P6Tptox31D8lNpHezcfxz7vJmVkqP3Wa6feq/NFbmND9FNRG7pJd9q6G
KZ37kO99yirL/9E2mKEXUlvTuLoKCoKa2KFbWpfZnqZCdygxm56RXOr3rk08DO3c5ttsVimXATpA
E/WMAjJHXJVaksbLkaRUjY4VvmQcCw8qrNKIzPLQOsN/rtovoxirBU2jLXrwVxvFpA2S9N/Esa5j
0UDiTAL2HwFlmS8qnGMAJZiGcpmkxSqGt9/Uk2NowAv1OmHQfhdUlmJeXbKIZYXO5QniwTnZjiYd
wW84De4TBUyIQcFbmRCIRVNNH6TUYE5Ie57WzCbImkGH6IORWfGPS/mS0tPLGX+mxC5FNNxOjx4D
dFLaaKgg9pezch/4ImdpvhrRsPd+s1+rpGR/Pc+uhkJuKnfyUdW2aCTcRWbbZqTJ/sp7jDQIWGPM
3xq9LN04f5uEZGH9HulNWbhofRCE+EZ4bnqosVdRRXSN5XBLpYBVK7X/9yJ1HlkFaX9MvoDxuLgA
updBVo8Kv/msB5nbbHAytV8YiL3A8WB9MsJVups2HlzPVxQQLPNQIiXf48R2h+I0+HMTvOVDT6N7
cGvWPvWPp+S2Th1muZJxaqYid18517XpyzB0HJKZDNTWnEHJcdcLkQY9A/rrdnA9rjNoG83yCjCU
syzytMcOHxJBqxulsotNjbKfPJ3pP+oA1vFUqDE3oIHr8+Yb6i/jo6NIsxw1jcM6YNZrnOKsDg7/
xr55ae4bhHQkVx4xNlaexUwfXdfrqpG2xJX/Gbd/CmCisJTg0Ddam7ERGlKtZHzKG9hdDBNV0Jhs
r4oo13BnjQKOKuxIzyXV9pfSf5jDj2gIa0wdPRdol75qrCmGPRXXzoARm+5jRuKTphJ3qVcwtMgl
cSx05BWmk+O0VqmKVsLc1lZBS0lV81bwjJFD8teXOopt4XFwLYUdBu4V2G/7jxwDck+ywUp7+OPr
WTBGmisxr/KxTJK50mqyDzwCa0PBDqI+ODJPqI2Gqi86obb6xULkOiyJO1Cqw5j82SH8roGcRRiZ
1fYRQnaMZS0/0UKKZXyaQ4aO+Z01gvWtgI8QrRkfAMVNhF8koFEBXa2RJPVQO2RV4S/Zw7V5Vkjq
tL2OLgu6u5iKyA7D6rLRz67JouAJ5B8aCV6nfRcSUZQ2A5Wr2Yhf4mZ0QjL5wYpAf15vvNc8LBDk
HCZ47qG0dKdulXc/kzuHY9VJZ9V3vWNY0/cd+24roBzVEN1rE5sG0xvcajhIa0qQ28fu9Iweew17
So5/9mucXoNc5yHLjI5ZjmMpLRLg4s8UYQ28voAa2eNpQwoBsXoy9dQm3ko4+39S4hz0IJafOgUt
daBwZTcQ8aZLc0l7CmVaU8k+J9TG+Zs/LkzviKdDwp7xMQmu9s7rvpoWL6mKJLIx3AN3SWDsGlJC
wFaVgzeIG+WebMg8WOG3qtJs6R4aG3A3fEcBkbUnqocnjDw47dOgUtF38u1LPof6cOtAeg6MrmBY
tpF33Ye8af53GbwyOgSwevXOJDICM0CQJmAOBiSiW4YvgJJJdPHpetEU1EJg4X5QGOoRpaVZ/VCp
qK6AYAsRfufV4d5NFcVvU7m5vycKxMZOXQOgpl6iOQ480BLjfjnriOFZ9mWvnQgjLc5Ho9EAbmR1
Bg52GtrAJU/kmC8605WkUs8B/hnecj+k4maS+d23rAFN6NPHzeQwyqHe82pQrDkK5gS1quwm0/1/
G33yfTDExMbxHv/XfwvW0sI8+U+3tKOf22gdJVOR8zYiNhiE+/tANZyiWm3fTMvBqrVlAKw8AiBl
nQHwd8l7AvxC5diE9MsMtm+iBa2NvRVZeuthZ7UMX7Llqk9el5q8gIploL9yA26QR+D4iLAuLi7R
ivb9CmouvuM/wlvly8RFRIiff1iFBcf2C4YEVx2F8AXQ+eUoixj8P1LbCy1DsX0U22wiJIHdVPwP
/tBnWkQTUlczeCcDsvZBo94/sbRogpg+fzOlnYqIV0GgapogYmkOdEoohzhgllQSe7C4xtn/+rrt
PaItNQVcwusGX7uWHCDHZcWVC3LqKrmE0bRBNbAW2nNWDYLzIFsDMldXktrpz0hj9fbFXM3oU6U4
0GQt55D18bXijhXaGxg8QyDOzzRKn0EZGSXSiMoX8buVRvMHSoBf3hYFBv5OKMnC0JvmoIXCFMMB
X58f+u+BdyAjZb7ZuyzOMDZPryi3AqhqODAmg/n2ZfQSCi2C3PCtpr67vTq5xq42OfGDHUoNJ57a
2aWn6vQjI0Yz4azT7FcBwbOC3dKljtzqk0HuefTgUSWwhacBbH3EVj3HMyY5uricu5O6o6yZVdCK
sgD0XHYrtStUFbfnwPXHuqFi0HTwt05sgWQpVO2ijDKfifqw2msgpk5Iw6xjEQh4vBqi52B1tqUn
VqJ3S84dJXj7cz8Px1fNB4RNvtKyno1+jpEjmWqr+xWF+EmgyRYWYzc8tWl1ob2jDJYGYPWyELTD
g6OKDfTxzZfxsy61PxKe4PB/QLODgJjN/yb+3Gw0k2goczm8PmW7WNJfeROzjmd3pTTjKX3govba
jvhxxWVKfNU3DT6wixunjgfA3YP/W5DA7gIllS5viyVD99kaYQU07TKFTTDEyIHBvR6rjHT5DCAe
FXpJMycIWbEsgCbzOrooxTFk6t2l8Ac268R2/N5VFiQNPKkuzoKc/YZg34n9nxG4pY/0L+39Zm7h
A+UTgC3NgnBIzO+NIDCjBl4ndp/qf5qVdvVYo/F81JhaKGWiHNxyC1IY0P0CqkVnIxnAFKxOCpr0
FvjK+/XSjFRyZCqjvtvkZfrlGAxQvnBHa3AmmTO9jv6y2ujMnCWbhoOHDGrvHufcwTJVLVgFaFvL
lBB3YwNNB5zXMDJKMd62p6L7jBdrGAi2BVmbGBjT7aJwmhcfqRfpYdnefIXBWAwswbaCaeZcY2Q8
1wZqDGoAFFJezb3n46PZU1p14nhrS6WK7PGNQZ9PMzdTBJLQQ0mr5hrBauLMpr+YaFSzHu6JPDuA
+ExqIuotWciE8PqNCPFEy1UoJ9JAoirABZvWTXjKdBAmDpFbFHvfbgnGPpnFebY3lAaffzEr2v/Q
7Y+/T81tb8IqVUr83ajfwPxKtQ3AMkRIaUZhgkhdC48LyKOt4i9GrP9J3pBCFcJRU1CoJ1J17TIB
dFvgerUtfGevIJwqEri5BHnMdWf4aC9YH4glrpIyelWn3XaZr8BwcYN0S9Qff5l+m4hT78OG4LU2
wD0xRx5LmgiFe/rjl0FkYJ6iI/38lauKYymNxXEAQMMJX2uU8AOKozt0YNYIOg9dJS2A/3r5Btsm
gbkBquywUi3u4rRSoRMpSqPO5EcWQaJM4b7aLqW57SjLPmsJRRS4wZqk2vzRBfWcmQGuzuOaY32K
hNOCBy9+iNNUxemrjcNGihrpKg+zNdoWl8LsM2AxirAOZG6/Lrh2VzcanZtsm8wSvB5kkTIvNcOh
zaTcyL3yIWR36OHzF1fcSlHZiBvTxkQQHqMZK1Nu8IQ4wRzuPlGkAuy8BfED+AZ8tTOZg/8XSrqh
ah31feMefdoz9uVGuyzMfZkCzFOaRjgowHB4UKuO1GA2bwd2b6q1H3Ma6NX+f94EvUJBsxYKqwev
IDMPvcGHik0AA4lD2zmXWp4BULXb7cEkPgoDw7s2BIAc0+isImAmM+LPFnWzest0bXr1PFKc3p2i
YEAIjheKO4elQK+qqRfd6kBAAcHGNUUyB0DZxwgC6ODjChWNBydv8r91P4nEKbM1ar5sajq1XTAC
N24uWPebJw1+J/9059FjFvEtST3z5qwIvIYkH9ceqpV4sf3IfFR9GkfokuVEHQTCSp3FvsG3Y77U
p9cfNPbW2+LZXBzZRMEAm4WQBerbyhzJi1e5/yVuBKYN7r1j4F/NsD4lFp6RLboc0eM+zz8bj28J
OZFfQk4dqSotrslZON3TbC3cplu3ISrDvlk/CNV8L+r3nxS6bPz3oZEmmGQi532++eQrezjPqKWY
jxGUjQVdRT3QVDZ37HN3hkFf2yfRIL4SP/XrgM5t7EJ/y0jIxO9zhnDmy92Xdb8hG8L+yxBiFfts
LgX4cY04maDmWyJ3dgaFECTo/6TTWvi7IL22HBefkqAzJqisTwyX/BQaUZLZN//KvZtxLep7kmMO
3vBYlH+5edBqYxjMFT+Q2iqc8t1dFXDtQu6PUyf+Ha7EY95RaaLDCAN8IDd7ekTDAe9RsRTggAlB
1qdFrsVTnvop0pEbl4l7rBcQJKIHdpNt82haej3a++mFsdBVRyhIK0wUFZDUfZhmkS9kJQdEltS5
+Lh7ZsPsf5DvbqUGnLQpa64LJf1K7tw9Su9iy8urabZB9yf5rLP+H/VtkCWE6QR3LELa6pEoovqi
DDlJgNHy5iZOzWlvpP3ZCylDuRW2sl0iAhVjXtnuuSYIqbxmjjIdvR0lvgMl2FBnVyBa851HOaHC
azCUvqY8hJDZbqKyzXYh46/xdS6n/qMYrZrk31sOKIxhsnfrfJdsIPms8UG9UyJlEnG47oybrjZR
vs5QDpJxCjjgxypGwqD46NU0us/jU+nycBsIqwiMyc3B6A7MdjkcikoW2zaTNp0uzo6Sw4n79UGP
PKQRLl3f0CASbHN5w7zDFXz8n7hDdnX/zeQq7V4hkATg5ty5mvq22KC5MuwfOrjp7Uzgn/luBMDY
eXhAmHH4FjE0eVcgBwakeG3DUfOPEd5YaZQn0rRodF21JUvti6fPu5uMDRMBi7Yxt5kMXK5pSTwo
L8Ycoi3dRnVkZnWsDPGHoGGICJ6jWNGh56P3P+NSbDoui/SM+hbpiOmrr0Uf46kY8gJspDDT+EfH
5pSJzXOCSjRA7vwGOT8lSHECke/2EiNWxI/100XAHvhoQuXOptO9lqxe/ZWZP0O4WBJ/uIhvgBUa
iznRSVrD66EYFynhHqocZ4XSBD9APra5YpzXhneIVmeqJyj+2h5HoHQX54YA1tZiZRkjsRNoTS9/
kCsD6AejeYYUpbzBZHSqMg5tKlqiBR+5S5MhaNtQUJZdodaNcGarHxVIu7+UJeZT/YfZ18sgGrPA
2sha3k5/7YxaV36Ti+9cOlu5+0OcWOioajTD/Q+HJLMprvMQMrDZFtOrQUiEM8aJwbSdrpGBd6FH
YVaGQBFD/CCYu0Ck55F6x+LDB+/0wRYkUTV4LGrtAtRFnlixvQOI7cEeB6Pvu2TZRwgHBoahMk7K
MuwkbL9z46Bm0CffInFSyqy8g0hPcgVDCUlUeVJ8e55cMxSS5QOwJqIBGirT6eEyLGO57reGpiwG
NBLr1EwBU754bSG7Pj6ip1pP0dAXFuxKXdSM1OcxQZtAtPt89zlpgRZ/NteWJWAorkxn1FNdDco6
ydX2xK8NvEI2hbudLOm3N63CsBUd1ujD2TEN9s1yadBnS/YE1A2CZnydI5JSSkXUoketsa/shKAw
NQDSo9S2d1ORl0NAS4fkvvNqfeQbdsykjiTQjay9FIwmhkJ5wUXBfBnxL+JJKcEsHNkbKHq1QGHF
XFf2lgWKMx5DfKbHY58IVyjCBkbNbRYkH0qQrv92EzyWcSePvfPf9ACnm6JmPIpjmbsXBNisiseF
GwIXL28wde7pEf1K79I4tXUoflT0XG648qxgrbTPMw+KZMDd+zPpNIzllgO4/PR6AY4XBurSsEyl
bMhI1moA3NkOOmD4lXbABSnQveF4YethmYK/1l7byeFK4jsFw2cMoLwTk6GzTn8pWIWWfqehxA5g
4JV7zyPL8lEfPNft9umWeQzxv5dhljp2RWIj6Rogqu21cgCQWTMB+BNiB2eGjfFBIFwmc9eTxYgk
Pokk8MwnbWsHNo7dVycH4T72GeZi11YKSntHA92RhumVvFNi7ZA6mV2gw92IMzmv9WwS82dNEsOG
tWqvR8CHFcfkk/f8V4s7xPG9heJTI2oRk2v3ZOWi1Xt1ycXTXSHSQu0ExGuHuEYERLEoA3TFrhDW
A//7qNafhv0CLKqbpDTf7fK4KI0NxfONMiQy5ZCfRKMjXU1JkoMXfGxt0OTigeLx9CAh9l0ZR67X
LMBK8ZAwnEE2LEAWOH/pNTDerJ+7axsIsawzkvAqF9ICAU+NGvplFEMNFxjomm6OgHiUCiw/b/Mb
X/Ly24BtH0jwfHO44Im4Lx2YtAoxl+fOa0YsNeMFjjLRD9r9WeZkfh6SUdnPQNQFo1YIOAZNDOF6
RTzgEx5XTv9s5CAf3uTqogqjpy/1Ia2YdqqS+lw+jCkfcNT9uucaadX0zgW/IrpnK20XNjuHtoYE
7XdZb2TAwMBgC1jem+qaW+reZ6PQtS/8qkBk6XrEkBwu6xxLhVPJlamoQSAymb4cBflrP0rM1LX5
0bmKapH2SWYgSet+ksshlwNi9L7cQY08+52jQG8/i+O9xqVfM9lk58giR6qgXMPYsY8USqjoO0H+
J0z6gDY0S6NX/Ov+Bz+0lHki1UTgejwcjhoWWqMh7HXjjjRQCdp64DUAg/RCdEmQrymPsko5QMRD
gdloqa1puxwIXi2O0AKLLdMEYzUV2GGge0ygqjdDnx3oo1+BhZsMMWi0ZYkjaODrKijpt8Z6jjsY
PPYeJ/cKKsbZ4mGCMt0qLOITt7BNHc/PTSYCHMdrEJHJqSD7C9tjYKx3f07cebrHwSwGmD/O+8/L
0A9pVOya3s0wcpBtnaHMelSqleBjHOH2ZPsU5kbz72VJbzPveTMx+0hdQEzU0aUtX4xUJW62FYUG
eCnuirRIid+qCyPxyWl3mE/lxfoKh+GibB6eTT8K0ogoSOUIIatlZNtjA2guJCsILnv+1J9Bh+ni
ziLxeuXL49aKEQIgJf1NzCDuJb5M2SbRYyoEwWkRXv+xJhvBPI8R7EYuqHw+txZJaXItp6Uod6xl
o2cIeVMdoSu46iV6KvPxP1bAiQqp0gtaC2eM4zXeiJXsPCMdVvtiiIy6DLzOa2eLMKzxAL3YqpVt
ELHkL81XMSuEbPTK40ZYbJDfW1BSAjWAxj8uoc105lbBIstdlzs+uab68iaX/3xYMgR15nFW1ULO
28/1Hwi1XBJp5Mwtt3NJViC22c5rXq1zfK/Jnq0HYKTPxUaSiJNBkXTojDYTfqSsASTMsxlBMozN
A8/PspcJStyEXzepP9a4vS1UY7iaziqlvDVx0R3bBAYl1EVgjt/C9aSF9ksXZ34Q6ON+yQrRDNQg
m6QrlwhTLdkVTdNssaG6txm/TWepy7yWcMuxw+6JpdUzo/oKXDrpBcMqhRUCbdWFHluZ9IrASvJ7
cXaq8dSJAscNeMDCfi5QffIHkm2svPvoT40EeoVTPEZ0QdUv9ltW+CEilylyLKGFmbFBjzWworgM
DXCBzK2xU/q77pmnUT9qsZ4CRD9IAHmW6DofdkHCGojBKusbsDvqxBFfn46kc0aCQlX4w51Cdfdd
BXsYtgmXH8eq+XaMmJ8vetzyCoG2W8HlyzcWhmH9uCHsNtYZQpXRQ/suO/NJndhHd+CsfRMkxACf
oWUYAREGAKgA6CpxXYfErs1LaNN9F1of7BUYlTu+g+olJvFaVf02uau8ALaOJSDUIRyV5xUkH7U5
lFEAdHSWzOS6qqSsalUh7RNFa1X2LUGPZdgmkFR0bTVRBVJePOEYfE7woXwjKQb0tA940COucdTz
+yQlRi7jAWTJMdI5txDAgqa7ZyBUYHmms8kAAeXAodRiPHMeQ6in0M2z5XMOT6nOJQPmEM2Ad5ki
CcyQJXdMjoYu46Z/PiOWYhrKgYq1mZFSVkUZqvkbggeZdnYsFStYyp8guusvTri4bEKnQzsArj4b
0SKjasXwa+E61KMn89RD8Ov2YfdesqbWg3E90z9YQbRPhck3YMfaInZ1Ha8tOJ/cJp8qWozQlkJB
YCY/woaownUXNWipPNiGGoD3ozsS5nQntMqPeUR2GJdM9qRqPVr6H/u6rAPyg0ztfeEuolZJQkcN
QJ/agDP3TAhPjC5A6sNp540sWip98vFsrsIraJ13MNciQFI/mYA/IkYgllU8hia2+aINrVJFbo8Y
iay03BAj47bLFPJi4tShFpfhc1Xu/8bEvulTq+StpkN+6ivRXZXwJeA1SSyHFva1uPPF7Tnx8Ogw
Q2iUorwNjzNzsyE29gSyvXIeonLC5/tDu4sCgvPKsKhN44U6BkdOi8xA7J/MGD+TRg+67Ng2Sxnp
IJSuLUoGZYqb7tf7j6cgQNVVMd1om8sclGC7IFf+X8OP6eqs9QemDi1W/KMI/cIsMtdj0AsojkFd
aYLqtafYlOgzdZ6Le6Dbajz+XkkpzHPF0t/reJv+mkhItTQbVye4wtExfKYGd5GNhkX9pope7kXV
tRCx10fhmfG+A7eABaB2qxfGIXPDw2mBIZJ03Qe/VLsy4onTuNrW4GEKYlssyhp5rWmhdqwmzatn
vgu6Pz+9I1ceBo/E7nkFr7CY9Ge1LqHqXx9FXP6R3LRIQfMC+q7rFeTikax00zNwrU4Ez/EzmojQ
jItwJKFJwOHzb84R9anWPhh58vXL5pgojRAY1Y83P/t8xK+PXy+KAtG0OGtgTMaRCuBtUs14IVrh
lWTYGexZXvZabw7l/BpdH989yJPbGK6xPyZD2yKoppe0fh7NYWs72BF404HTz9DEjyvKWRk6132O
pmhUXmALPqWIozXdvgnShNb/P7eU4okDWFptyBu2tbrqvA4g9lup+RgSQ6/ak2c5o044riAOK6Cj
GruW35jYm+8pR3IkZJ+jOG1F3y96Ys2OV8XDRR0qJNUsrjS9Q8KDuVJtQpuhR8U/ULOO5BXj/LKa
4SAAnapGXFIkoj3kWT+AE+OtlgP6jAmhFxKtb3MIHXOzr6ZNZVcTAlRIN3jYwW/7k5V+wFsx0uxC
qU830VEnPtGwNaBVaBD7tCsOL0GFvISS0A/vvgOYCaRfKS+3jqFTLVhjRjNR8R2KvvGhTa/ZGmp6
p6rezu/Dwy5vcMuBEurVhviQYPPq12Du/2LFyrs++xd2DxJAnP8G2zImMeeQcB9dKOn9cMykkNLu
4CVU6HS3+8sTtbjMaUin0T0v8CakOHQ7J80wsrcC4ocH5YqKWuUgOyb12IdLUVqq6IxgvwbaUz2n
JcH1MBVBZeyqu0/8QojmM/meN//3S/2uWiM73fuMKwC96FyITFfJ9KLrSD80qUHeZgltd76nDZZ1
dM5dLL3y8h1KSPNfWoTGk0FT9TukMv6NTgPFzFuZDH5rWC3YAaB+6RY/sDaa9IJCHYHJTAuII2V1
d/j3rxUOHYajxdkMW9zOMZjuoPxlJL+DahrGZjM5MIaJt0a85M4WaqbzWr3jG8XCED248eKMKTfa
X7ixK4ZXGJumuuXN4kmAHDSu1c/4Xh57G4rWvok18/iFzD9VhIUAQsP2rQPcz2l4YY93mm6qaMcL
INisz2MY2kQyliz+v5gzD6gwkjCFgZEyGSyvC/INHRp2g+LK2FN7guGGbSo7/KmceWSh5cLXJAD4
UWa+rd84Lc3apwP7kx3eXi4GY3+1/VNQs5MQ6smrOlCTMDWyRQ6dHWjoZEdQC+mUxPrxa3/YRtai
YnOYCe+dRVBNPXaRcbOdqUL4ftE4WB9BAZ6s1X8jLSHFw9FTic+zFY6mG7RmAJF/Z98u2X5retaq
c0k7J2Ue06oyFCzdimt40y1j+MysCNm22CWo02I3CxQ2yj0UWK6pI5X/+Lw2FTGp6cTYYnYONqGT
PsaSinCVQWgvSoSHC1ovvcfRGKdtfNQmlrx0FHQvXYVhra3koi7lwAWN4r89lhPC0+DoiTPz0eRR
1ottAIKNLdSIg46Pn6alq+GqmZ5Gv/Kkclv+fs34cHzgyESE8gUentbkuZRtUNTaVICn/2fdE0Cy
6ZDvnhTSfHHtVaZak90yKxafg8LAx5om94D0mI/g9oC9OuQihpLQNBq53rml5KOy7QyAiO/ZDYCN
ocTmOib6Mg0QODMSwxJXlXcnO/oT1mGbaDpP4GYv3tbpNv+GwShAFqjseN//TTgQsoxqJgwjrfRA
tMy7TJMXX62N8zrNwRGxtAnWu69/HiTDLCY9xS7C2frjvS8BqAAM/uZIpUAjmZpJwssUV4tNXn0z
JA1wJpGKto5nai8q1vZEWO+Xx595ZvqIDLLVPKQbQhzm7yQ1KilahRB7swxTyBd+0+CIR6wpwWCa
e26mJstaxI096+94tKM1U+lsDX0ig/kubseHcoRyU2cx2VoTgkSlxsISAK9grHVhtollwF9t5+ye
0HpeL8FlR5xvxBtiGPgOqdiCxbukmEZT8/HgbCpSgNMiJtJ8E0w6GAz+Q/Y4MG2XoNcNyZ/4VabA
jx7WI+soWlytig/jCUJN0pTox7oabwVzRYGw2EGijyCQ1a5MBpR4IbEfhbkHnK0xIqGlnNiPR/O0
KoPT3uDfJqlkvgLIsJ0fcOAD/pLsrLvKhiWcFa/k/Cf9yhHtGOhcr8ZH+G8uHG/rS0yDxmbz12g5
0HEvlivfeO95vXzSbqlMKs/ILqUlwRpgH4SbM10yOqoj2x7ItI6WU38I2HF8nnENGp/0S4/tDDv4
j/3sRIcoI4yTwZYgRpZP0Yk3NL1JmP+C4i6TyV2qOFEdQz0xTcp8gkERtqjNGsT+H3elBbTU+ubi
Woz50bwTobQjBWdXop/SrQ+Q94bOWR3j2uIEx1goQxcHh3PyPF7cOQGhA8M3YLSx7Unu2auQcyQi
emk4m3Q1zbJ+IhzZXw1a17IP+LjcZK2bn/Vapnx70f56JzllxtWQ+Gg6bV3RDOF8siqjUoFyFNgQ
CYsuN/Bl7Vh7nRE2zkhj1yfHfnZw23zfU/dX5GZLvwGA/by48b7BUHkIDir1jx4CmTOvWbkdLPyB
SH7sjY4bvDg9LBiq6beL0kSnf1Q1fZwAuD4fpvKNjZ7XbcQsMfcfRDoF+788zUr4bheyQrr0bpSJ
Lhk1092j0MrYffXvaPYrxblz09mXwugoFhpWpMq8SkcuwBY9CF0sGTUsUQLojIvg1bSrggkujBJc
TPxV1BjNDpp9zJQTX/df/qEOlpaihEr2zkksE1haUDv08YwJe3P8a6PGBGg3EZCwjP6uMy3b0wWz
bZcE9CltSdq+cGTKraDMBTiDwmbyjaK5c2CC/TYaOmFtHN+NpQn259UMJ6rVs80J550nqqEEbped
0tTvDaU4kX3UbLj0ztttZ7qsCjLEJYL6St5lB50D/054sH2XUAyDq96aZZQ1jUhEHYVK1wR0t2vB
lbrnuV5MEJjWj4yOBIK6D2i/LYZAGaHp7TWf0QgjeEpeE6qRhldSAEvQUkuO+bnBjNr5ZeL2DkIl
rRIsMdcFkUhajhunRryCHwv7WURqbZdIaCQNwRRF3atkEKdg53miYyJVRn1yPfyuTQQfyKMfXJK5
tbOW60OGCavyrW659X08NKbsigkkDhhv2UNAxj5vhHmG+QoMk/R+IWOrVJB/D67fvxcU8OEzl0vo
etWuzQaP6y2DGErpZntYMrbklpt4MSEM4fAVSB2zMXV648UW+Iphy9+mqKn9KUc3yH1v8QAWD/BB
VHSIOnZ8ku3AdW9CMUvxYxCvdwmuAoV/efPuwU1xgry3aPr82VU+rNFmdf7KOT7ycg0ZOVCgTTQA
55xbeEw38nVFpEfp4/9iEAbzISDfCTAQr/xDgn5VXXLcj8Pyk7kIeklgvchYJWfKJLme7LeA6cU4
XGsMSLwpdMhRUpQc4bKYN1mzXqbXfJn7lWheL/yhB3S/xnNDBBxC/QjVPxCDJ/I72DC6qxUMFM4+
wh5ilqnHFHSvRkjXLqTNfjzsSKBTFyIh5VcyYEZxmPj7x7JoMz3bJvRLJqrfbUYVlBwnIE91B0TS
V54YaAIBdzU+PJEiIPO/yG4QaWmVsg4PU0Y6qPvqsAvHY9OBktkqs6+XvauYEYHQxLjfTSLXB/Ti
SUJsdnBqUgRMnTiQNvUHQBCSJlAWic1ZYn9LpWHaSjI9yWHMZmXOBsi8WdUsj3P1fDsaWb9glv7N
zqPWnY6LSmzIZKCkXjgiYxxUiqrVrbUAfbJK4289aKZ4KLSsvQSg6enPJHAT/b4j/MPls8lB+6+l
/SRJyyc1NaqUThDbNWCV6GWFkB+QLTqthjcF5LuWfbkWbpAbGlR64rjD35T9DV8+PDizaLBJvFNK
4gNn1l5T561Q5rwuCtReZYM1kAAWRXjBUHuQr4kd5KrX1fSW+PY6lEkn+sGP62/oj+KuzWP/uA2H
ZpiZOtniTbTyyqj0/06Sw4p2TAz9HIZ5BAZVT7fQ7wXKS+eCgTc6EMVIaqV/Uzphyq0ucM0n8b0i
EZysGV3VtEDFEMVXeNbJpzPBZZfGTX/Lr6WY8TViMFGYYJu5c8irecgS2H+0zHOvj37eO9721gb/
hG69XWBAj/XOAFiRdRgwHLLtb3YVK5EFET48UbU0a+tmGxkbRLZS7DjKyWeHFzvQ+mvI2BllDJ+V
PqXQHltmdshA1ko5wsONtUQ+zGLzv7N+A31W6Sm67ZIo8ljJGLM+cljAXR+GKiK3AWIFghoWregI
SmWFCPITSENEPyrlwVK9IBjaKZA4FCyawzU/xYDNQmM22MNm3ZhvfmjN7IM9P3fJp7176hl7wjYF
6tVRksM5e4FsrTlnCEo/Wac7uvH9Jmh6KcQ4S1/Tc2vqUmJo4nWGbgKYB47FKRNtt5gSRIjSTQE9
F93IblRwxzIXu9frwNnbaZLEDTDPxz7Ms1hXwX1pu+SSl/tnMQBdN8f2n4LNgLleqJ1o/B7yChB/
vQ7LRKqa3UCmrnzK/x/CSXizTnrI2cTrPyXgKkVGIuCRHmBsKWmOj2EWJKV35izYs9/VXD2xA8Pa
PmF7bLMmlUZMekdIZ6YRSp0zJgdgFnW2ifqsCOODv3MBb1S3SpubK7WCv6l52zRk7Ajhcopfp3wj
gZWUtalG+2yEZY9SzkkJxJLA4PVr83FcGZjMLvixSVrkKUbRkN2WDnFtyPbjA9iyYXARskXjW+Jr
8quy21W+7zLNxXLeD5Xl9tgIaBezCycMey6aS6x4d/nkTB8Jx6++GRuaIQu7Z4vr5H+WxxLeXvyy
ku4a3nv1lOhoK9oqEWKl1v59YFYXL46J3CUbAiignZwzXOVJyhBzVJPdLEIrN08k7QqA3QVPBnQm
rtAe/D/I21Yuyq1dD8KB5qfblUJEW4i+Qvmj2VrultQlEgH3Ar9xOCdaE4ID9orvJQcZw5+4Hjmv
yiGvNR1OuLIT19KXJO0r2CQPIMdEWYLV8ghiuYyHv2a/Hz1j6IKBkOAZJ7UH0ruRw/erip9a29kp
QpbLenQ0Z7qV3s5r3YNx925n6WvrLl9G3cTGOl0A5+f3KBxvPY/gb2DRoi4slRHEmPeDfjMlcbLX
2tbADUehmi8IaXu244rcSytAYuFnLtbt/ZYDhmZGVNV6kRqx+7CgmyURWEE7GYIOoVvTqfYiyF8d
zOPIsCbl15s/0D4IxllQSrrlR+n2xy1+YWQL3ncGs9d1Vc/dBcqtMsBH2Lq/vNkWmkVwLeeTlbwG
IgPip7TEAvPcFBFhXtZEfZuzpbiu/IGZBI6M3wvUGlxEWivOQJGgNpyBF7Jbme1R1VOkWVdgpxQX
EiNumipUzqIE83slnrIuLxVahngXUrMm+PPa7qz8C+vxdm+ApD5yueqzxj47/8QsdjcH53T9h4TB
U9Vq4hvHPsemCifVXMC5ZS83qAahOjoERZa3hn1lmvIzWtrQSWUkw2P8BRH1vXU6GcbiO8bWvm86
JyoGL01LOn/6ywln7OO3PsmJydi1AVx69bF/7M6zGQyjZbGWbiX5/ruDLk3lcuCGDpKNCJwKWwpA
GqcMSS3EM4GLcRvVyiJXS0525tx31tUEa8w1cvgFTWeZyp8Vwr1kZq7aQMBvAVBqmJ/i2u1+CU6N
GGkSwprTJOFk+gJsJu1GuP6hq9gpDHnEKpBxGw77Jb3q/RaffYu8nkj+C2w12of1LqabtkvNpOyd
gBztvRwZND8P5DRc7pNQPkCeXIURJ4nBciAivmztBmGsUYE8Po8QCHYdhen2X4kQw7cHePUILGbv
uB8nE3TopQHW7f0un4JTbLp25yvVAQdEdWE4C6UVDIDj0VdZdLfrw9k/Rl6yPD5HQk4fcoDozsi1
RUyfNTvqAG52NnOnROQt3IPgAB8st5SQ+93ssKgapEI54ovo4DRXatyH6bVMZN4qceDbe02A/7FW
1viDbxu8VQ44F3RlcWhPl0kpoRb+P7br02vRK55VOSfoZeHHXu03qBmP3MX4R7YT6uPe0XAgyhwC
LRaPoJVVPNwhUpcLBpwyp0XF6kMxSplc14+nuSYLtqI5wgkN9Wx7LUSGwTxx0uthGjX4MEwavzQi
QEIuEIBj0zQZgUDHbtK7BwWi0WxHMbpFqa6nC5gWv3UiiI29OMxit39icZLZ5lC7EscqrqiqQgc0
3lT+0JnhXkV8bhpUYK7EjBTN8P6i68BIXvrzu0FEPNPkt9pEi2YPtzZzi5oAz8N1D7Dcc69zCVgl
phXtBslJLOJ85aoNsseiJ2i+SujUgF1ePzYZrt/fQvCC/byB/8Mvwfk7ILUFUocrWBc0ozO//fEc
twmB7dssXAd/j/lDEZ1u7gqET005dCRVbZ8HuTAbVJs+7u6ARKJ1jKH52CpqBPRsBQR5YIkoYeVL
ULfr9Pq84sjZiL6s52E8+HyrcAYp8hfaisNzLCtMctPh1Nw9v3fk9qqpDAWD+P5VfGjyoNgw0Fu/
hW58XHfPq2wK0zOeKt7eZo1qzKqDrFk/W4BSFj2xBwpCAb2Ed4L0hX3XwZJuNN7dmLenVWDWYruB
Ud/J6e+y1s+XWDqoCARdtmNoc/MHgIGanm49PLrA/82UsPJUyIpLzh4L4gWXCxeqDskt0xVRPGW2
EkCUUY5FcbY7HefKWRVcLVTgrAVNpXVngdCgu0xvUU0zzSg4DPG6EyKA2kAxHaORtxhWuU/lRJS2
vMPUM9LpnaJXyjmhD+H9GDvMDuBGHymPpjaYRE01f4/aX81342EQdUq8A8k5G2/xGkKoNOhlUAq/
vSjULrMF2F9BZpHCiLi9a03omvfJT8VDR6o8WsCAO0xUs56pqOrXxKRtKpxx2YMqK+rueeAXaXRA
vvDzGH3k9orSob+yVNIHzj/y8AtG+JLVzQYBguzgIKhTAhGMWdB7U8x008SBUUMwEmaJxp/uA1Cg
ic4ddAd2xRyvdFNlliAafSfrJarbvloWodiZm8DIgoOx74Low4NlSY1QeHiG9LADwz+KED11mm9I
jAhaJ8+xbW1RbD4B225jSaADRitf0DeY6LuRWlteHoA8VmcjrusnmtCu40Q70Skmsa6TylMHbWm3
rH5z+kDXFi8ZNStXbMo1HuX7lE+b/Nnc0B0k5Spi/pOGq0QelM3rHOyjVxGJncTGS+yCErfbr/x2
QyGUqhEYAmDRe1zg4lhxyLQmqOeaBXKbxVzVeK62o8wGHIgfz02l8CvUtWaEwaze6IZQDh0heNL0
z9RkgdCWWFMtmXwQ1vLHWUSbBIAxyzb/wsf16DLdrKzA+Pm0tG2jh8Df6gVvqAxH5fcUJJXbiE19
xw6v7QjlSpYsm08TkvvgwsJ3SChKOhoeqTOB2kKQHvOJFHCDfQwPlrjMqMn8HbCrVNCUwji+yJ9w
GpOdHdsPFFuP4QQ5rP5zeXW4lxRffSyBhkplorrTVFkCO/5D9xddoWw3hAWROt4W7+Iqlv5rqHf1
HyFjKGn9jCpOqigpqMmA5dzsxEA5o7Q02B6p106M3DrsresHmWwkszEoPfA3/Y4eS9N1cw8eh7sT
3OCfeZ0D1BDzyK2iQ9knTlIzBWa+C69kajl9wnHZMwcEyddR8HTgLG7cNs9Z+/NrWjj7WA3TGUoG
kyEsatS3b6RlzIJ1ggoh6tLBldcVHT9nQcikbDXrIdPnoBRzRed5YCffv4rmQvEIheM+ZZgsvYVA
574CguywSiBABgL9c4TbP8LPBSzE50dxRg/0xmfsXpG+p0f3TPU7ddf3+gYK7ktmfSRroNg6a2uA
huXPGAsn7dobufzPDs1aCj/01TtM4WkeXwbKHqzDYb2fCjGp8bEix4e2MB+bjL+wey1idi25zpV0
4H5TQuWvz5ZX0PnkYDtKnQw42nh8ktzC5eG8l0cgZ4tdwogWryuLvLV4Voxi27wb3VXMqxCv1wBH
5qP3XiHeA/ySBhZIOxbSL9E8TUXRrKYs3uWYDRt8270l40X9w9HQT+1MvE/ZrW2fT238Vut1uNY+
B+79+VEBjnrv5H0z2HJaWdlvLfBxtYcUek/Ga6ot0M47rLIssGnz0747oA3QhhfBV+QQg3Hq6A7B
xZEy7z68xYB/+dnSlm4T9DHQejJlCV7qb2Px/C6ySrFE+AG8GNuVW8RQtB11sOjHziRusUAYpWS+
hXCRL9aBhLGWqfAtr3aDLdj5373JM3zL8Vf092bEwG7kGxiGb1zjsMTztWZyMcKlFOESOAnh/wd0
47gIg32YrAPz/E4799RNgFSJ3Dl8/AbPAFD/9xXW9/HGChcSZVKt7p1HpcSWzEDl5gnO6gCyAESb
jdJhw7wVToMiJ/TlWY7EUXjYgLwMz1XyYorNoDs/i+0Hk1iwTPltI1mysWIfvTM3KF0p6/ir5bSJ
CXZ1EkCsUkLnhNsA71c/vhhv+rKYCzfE6Sj9uF5qWgKFubGpVveOVWDY1M0JEfMhfGWxLMbbiamU
IeqBLuXb4icqmLpaWbuDGQoiFjje+8T/GPDpWDJbKEDd3iTRR7Q4M9a8yljvXvPegMhrADdjbXKs
kXCJU4d9eCNdvDHPlk2Ntb74L7vZa2R3VMdx+a0VxxWq8BoLL+N2ZQKeRTvK9yBQNq/pBtB4dVkA
+eybN4PSkLx9QayTnM0fMJOSekzCiway1RV3N8tAN36MpsNDsnJtcUgxSuH12xHO7G85ddyu/RFg
UQk6WEDh3NrcKncowjyc6HC5RQJaxEmpOnIqZWd0A5LWtpIwCT44sv4V5IhhuePHrO/cPyVQxiWn
iyzb8Ulpal4AzQSIK8YV+wyS5UfafAEN5oF+nP2PT7D6CIG5u8GNiJfN3+Ehi/Uy2XIdrdMIrlfY
BlXF4jnRU31GJTPGBfEcjBEelSL7Q35d4ZA5X834uFQJYmTetXon/ib6Ma2OOayhAXDMi4NcdN+N
VOA8yuoHRbDx1WylRVnGVLO0AcynumlL+neZAAk09fZvYhQ1Nft0PKnMYxGdyhK5WejlgKvpK86p
19nWL/dsV+hnlynxPdrwlgxEG8ss/M3qgcIdAFE6SPaYS0ES72/dTXzJKRduiH142TnLXy9wrjZR
24/OwIH3lHkRARNHXMyc+kzDEDLJDGPiMUPK+CprGfMoZ2t1C77GjZI7vEjpyiQPl/G4PJSRjvS8
TVNBaZyxoPoZZAlBKmPoOPFswc8vvtOw1X/VrqpuWzIO4vdedH7wXH5pRxCT51o5ecznMJT+rUID
ws8J88BMbFFaZcsyhBPsWzqus3Guit0sywEW8mvQVehPJUuDOHcKwMdUVg+/2luD6owUCd0+vhmL
jspz6p9UfyDVlN7RjbnxTIvsAkrgnNecuUsSTw8Be9dbuxElrKbUFlX976mXGkBk8vinO3wWyJQD
9W1NwIeU6oRvryIa7iMcJXAcXadr6+6nNqxuSRM2PTms0cxERGNrP1vaAD0qOYCx820R3oJZDRhG
/UqkPKVIhGSz8o7mVyHvCNIEOGq5Q1edV7ch5HZkjsCTrNLGE4O2ozudN+8It9ES61J9K9VgiRqi
OnzHUrIiT+EyRH8saPr5rky96FHHVbTgllYMpmiUBm4456d3H9LogLx6iDGzI1ZPxqy83x45RRcM
gC7kXayonjmViUh0vjw/eJZ0C+OE7/IrOSagR3jFj6ZklRl/Z+1WNeQcjQGmQoUC7S1RexTGn/BV
0Vhm2yzZqGhhZwMLMSPN4YdWuX92cHE7Hd5+u0Rg/q48No+oMKMasFtO/EFgGSnSjxTW3Jdyfh0n
rAaFE7YNRRfyArZt9eqfqrLTgoYnypzHkqSt0Zz3zrUfiKnRPex06TAYO2mq9WOeOdeAP4tplbVc
mYt7ERlsSVBo9zR3QlX4LFpn7p08sd45LNlobJc4eiAUV0mj1Zf7FAzOpYRACdRp73wK6XGL5nnZ
plYnViS4ypLAE+gBmi7W34ngnc59D8sFw85V0PtwPZNY3vdLKJRguxJ7/HKS3JPC7TvIqrVOHFPA
eEg3bYWzLY4uI0HtZdrbDttAFx/55+Yt7KJDecV4EpO1keEOEKjOij0Y7mf0oT5COVvlsLCQYfUT
t4+czBz3cnT9shpQ0hZ1bNqeKsE9cQUVz3vlZmuKbnCeJ3k38ByBavQsbAwc7Z+o1nP7UIVzpuM2
/63qP/8v31gjIxD5lMVua4B689aTy+P/10BLvRHIRBo3Afryo9W0mNFbwAwjI9phQZZkSaRdUYk0
Mxln5R3vNDOCjP348uzawlFXLgwMn4NGBWkPaDVx+fkOcaZwSMeg63c6ip+UIgLPVnINWxmzAHiO
hsDLOx1zSnEE8rkyNNnDelES/8YWR6zfaGgSAHV5YZK4mRVZXe4NLsglcJIAWZz7OyJqBJXb1Q0S
dL0uXqWGPrROc30NbC8LIc4xc1LK3Wd/SVCgORIP835nXT8HJrI1W4PVTjVhBcJSx8OX9sTY7x4g
soQa2d6yFXiYrAhc9wVJdeI2Wx39juJ2LPFJVx93k5KnT5qqFTgUyWwjle8PwPMaYHlUZjjeAo6E
g5IY6ZDKIhAe0PidUZysgBEYswvVgTXoIVPqsOZAlaur+w6N5yFhFRtUa/zhEpRgDsbRm9nAglqE
fQCJLP68H3w6mr9LoXYarS+URPn4KYB+NpEcCp9kZMxlR3koY5j6nXnGIgk8VWP6guWjav0u7KVI
sw64NvM0tsAaeM9ttnr3Q6UjcMWMYzwYWvG8zO9T5A9NsH0hfqHivhHcUhl4fXsmmEMM3L0MQPQS
mxBxGm8YM7atShaRkrdvaYfCOXzi3l7QVLukUUmYELSC91ymjSN4gdQwimdHDu76PBfZPwWlp2i6
fu9LEid7/EP9gZ6Cf1+VCSEQtN+EfTfj01iyXX1McWd1sGtdRKc69BTM7rd6i6ORievIqu2xY82w
3XRgW6C8PLxOfW5Gey4kfjzrimKebs1m1ZZKC8T+Ky/wSVV2th7stORP7Myp6fQbBsC3+CXRT5XH
PTsyJhwFMkHtkc/1jPOcFpxzpSHT1dprVdA7v8FH0Cy5NDC2LIQ1n8f7NrRinNAvetfJDs6+3+j7
6rUrRyQRFofvLopmvK7xjH2H2vZgqh9e9jh5HDaX+XG7DUATQ4kmLWlp1t4gTBrFfJdzOOgxEhxE
kMz+gpWJIjl5PRO4L12Eg6YQpN2SKpTzt7dO9Kl2IJTF66BVNZIUFRnvdljFidF01vY0lsTSH5ru
R5wIXiKZ9yBFJgQm2BgdD1+D0L0JrBEeTxKcKeqTzjahIjIKpMc1RKD7JGY8oaimG9ry4W/yBhAr
O5yRhs7ccDMhCTrPscknoXP8ukAb1GLCfYDMUuzN+7HhwlZLjkNnoQ6hEZNioELfp37jo9xgnIdC
FqNfchgTAtqAtWWhQcuKoifhuAjDZNLKTHrPR6kYGs7IU5xseRGqyF+h52k5JFF6s2WhoVj2NiuP
WmTtl2Wq0dSPAL7TuP4jbg+9Gnn9VFYEt8pqOwbxlTW5pwcBWJYGyokKqof7CNBAbMTOc3RBL/kv
bOJhNObIt6CWu+7WFeKYAL2vMpmTbgZ3QE2548Sp6c6MR47X6y3ix8130OGlPt4gPBpgJ/nRjyIj
yz1MB8TBX8H/CHtU5lX1HNBlC2YWwj2UaAspCiEoujcca51VknvY6r8UYmzNfWsS+kFiBkRh7L3N
XQ3SwIMBVAGpz+VJR0oErx3tHXrBYfY4zwGHMCj86z6GPYpO1fG8pfUcYI+wvfGDaPcXzwdsy+PI
CkYFQOzd5eiNxsje8hD/JM7nuNYdydTsWzDYK+GiYZdG1e9jS/wh9F2w9DdtrUjebZ/BbogxLZiD
1yKj0VGZTF5uLCb8l0f4urGEF8s6cQYWJqQCXEst47bB1+8n+xLAfPSXsVyj6KwHxqBkmihX1Wib
8SoCTyeDS9dKgLmDLrsD6GNYU/3pWiIa8fGaL4ueGrlu3EkpymYmFTlVsP3A7OYCRcg/dHgqELof
4US9dmGjj8yzK43niWtxst1UYWVbc7plMT/LZCptzaTFIAAOhB48Gyj8MzkIKnOXtagRTKe1cOMh
0vpjvmFi4mjQdWA7fJILrcBfptkNGPQrBI6vQO8PW3VyuXEdRhwiKNI7VEQAG9dqLb7cIfQhib2l
2ivhgBcYXAR9ZMJMPhCWz1R6NfQrQ244PkxOMuxnTvA1eFjJMN3+piApBygCPDhwxuOtOTYKcNDr
/2HiaqaZEggUSQRSvowXRs4U0yd4hNnQdlzy4fFmV9FY3SeYIMBe3A69LDinl518M2QUg1i3hBCY
p51Qqi6I2S8xLX34vItHUCAlF26Tu7thSBpia0Kp8FmKp2tbAHogk0suGBTdamgzMord2ENA4Qge
tj3ZB3x6PTbjvCXprh2rRCcVQ1HR89QGKEbu02j18/U5sZ3K/J/5HsWEcBkgz82jWQvKfa1rb8XR
omXSGr9+VVkcr9b84hZxL5cDAPMBxGY7/5qCoY7tXRCE0/r9MZ8v63lcWTAsOY0YD6EcfIsKv+eR
mN4Wm/h2G6wMq/wy9RnHhTLo1WbbRZiL+Lf05WvIPhXjUKqFOEFbxs0yFfglYBNXWkoDpNHoGov6
LBDOanY005vGXDFgVW8lvlSLPxv74l1KHFZjJgbLaF51HAs056NqrlDwHrMe07Z6JQDOrKW9kU1B
8OH5khKloS+UBl1aOcpcqwJYk0cfow3v7zR3hRV9Vo/yqnpteFRlgzM2rlWYjMxGs4UpEZ4diIgJ
n2LZOuzzSPHYWe6v0a9irz4tfyXnmlRuDupfNxmmjAeaiUHt6uzMi7iHlxCXV1EstNDWbzW8N68k
asQlYohuwzXNHodCCSrLfGtR4tdKYNpzpzx9AoqaZolBY1+B7HibopS4ZwnRusnufGz2FX/CNwpG
wbFCMUmgkt2xNfVshY8lmML79pd5KXfG2mnb/bXMP045ZIeHKxQTGPHj5M9pR4i9T5Oz2gS7N6be
vgq7Jh3R6A3D8JhOKuBLQ/tEbV2NXsh1O4WtxcOaA6H8Z4U4ijM449L4ZZu8C8cKVNbf+ovMw2cN
Y9UdvS6+ZetdqpMbGGVUTecgzlGGtPyCU5t7YthVoVBnTUtkFsZ0LPdjwWms/ttU8M6WUujMEWZx
zZoZpR53O+9oW/ExL3dxb1EM+X9Cug517aLFvoKa+6uUDen+iTotCVNjoAmQVFFHNwNa4S8fB6Si
1Ojtu95ndhtN+ps1plFRNuLziIw8KYdvcKUEdL+y/FMreJdBpeH8ByWshXckXwxt3dktCbnjXBA8
ZNReAD+KPFy5ve1RxLFzsEOD1g5nqoSJI5FL66se/gvsb+NtaFzpSujz+9wty0v610IBgF7UDHT3
78GmYwVnEeHWHYGEXXmSLsHQOFPFMXeusEoqs6OGdl2YRkfgFICHQqlMaJs6Nsd6XfQ6zmj9Gets
EAEKETbcpdZcMjkwz/Ujf68cngdusJXY3zTHzg9vnlg4YYTKNMincAoe2LsdQqd/DaWSs/ssxTRv
arwT2B82drU6fhn+Wlxd0Ja79VEOmSCPoDZytx7w/lL5WW37E3Ab8kfk7UUQ2Am3wxfZHwwf+lw2
4U/GlNZn9V2dfJDCBzVOtvXl1HuRCNxO7osw/mOzl4EGbL79aHre7UhubObV12LEdtrbZPb+LdiF
MRKT2tr2SOCCqxHfy/Izse9CMKZOTo47Pq/VOMl6SNzzCd5XAQQVFhpHAALMmTGzZ8WLUAQb4b+W
B2I70ErnxejftxnPYT/mP1Z85fRHuci5d7ZngEIyEy44R5e5r0sLCrDx1CPDjlLGMwWddPPhB9nv
Sei0kacEwU39V32cdaxRWIuIYusRuHAb/Gomf0XtUOWzLNoy9cd4oBvrqe3bdBr1AV0Vs5VfLf+/
0/k4MUsd/+xr9Brvh13sPoCmHxJgVasXlBxvO7jYINXPGJSq50Sz3Ka/YxHh8nD8QC/oLUID2Osk
jNuvmixRMs98MnckEWaKSrFjnXuR6aqS+EFVUEBVB/88yiuvhBtMEQ9DxD6N1t3NCboCBDAuzzas
llLrg0IyHoYXK+GHARmU+4SCFi114wt3KRIqJvQgGtBC2jIDIDhmMgVv1PfspI/ogv6Weoe/O8x+
XE4KWCKoospnr67Dg4KCGQI4TGqr/vPE8op7+bU41W9RKuh9bh+pmKWcVDwgy9aiSxtyFoqn+1Zk
UnpzUR1uZJlwX+XfdQIQDJRO8qGsCO2L97A8nOKqc1wEphpc7NkntTw7jU9kqeSCBQotgrgBNphl
n8wo18AjI3u0Rb3ZKDpa7bgTLj7XQGyJsIKyk7XzUNJxgtHCkIfZpmk7Dp3xl2kytIuX0xaOa3r0
TIdDHwlOlLvRAhB+DnMBZFB/Ak/I5zhjG+x9iVALChLShIgCDdMibuZ4iC6AeBvO/YzAZLtmfF8m
AvaxOaXJf92V6yYOaGDc+/7tEiWchT9HG0KJXPmXweSUn1DxJt5AUwJVQhhx6hAKbBEkyZV43c8B
Hi/7RPA0Pw2ITOOfQ5eLin9Ny16XzTzp1B3QGvFO37LrLa4TtldQR5YwH8BD5n7gD32tgPzVoa26
oac+rEDGnCmaveBDrlqE1NnAo/lWXgqheAdwxOtnHnhJ+OrxXUY431+OFD5sUApd78f+D8BQgVpa
5dlQRbjP/O8fvHZmUDhJdzv6TkcygWq3hCws1YsR7Kg9kUYWfwl7bYgW6LYYsVOYUaytNyIZnx/p
MWZNKi/oM2ent5RxC3wQUF4jJp4nYiSl2dd8TVAZEFjHAFIgWhLaups58bMLehO/ow9GhuvveiLF
8bfjTFgGorsXqRbEBq9mPpYhsO7zu8jHKeo+vr5odF0TjpBeQetVCM7Q5kgyu2zQGTgezkfky3T2
ZcaUP9QJRIIwP7QDAA1ITwzKsQ8WwS7UIhLWBCQD467bPmWzXrbSdII58Y4pXr5PuQNtlsGEoukX
PGvPANzX6yIvXr9Pv6hDzUUEPaVJDZGD0l6JGNqnMvsIwx5YIUsUngJnUj1ggOi/zw1EhzK3TTWF
NTjslFi2MZvVZY/1S1sWfgvAMo1VJvIjzCojFerTJgs6lj2XOrdrdd66m8CVRpvnABBjjSj7ahl+
x4g8cI8Wp5xCp86GuaGmJFGqLpqiTdeWXSG2fHQPnyrVlHgWq/pd9AMHO+R7dYaY9ZKkdT6gOquJ
m+rdztUasCo4AVBILfdyTuCRQvBoBPDQUTrvyNCKRQFsnpu+x1XaMMxrs0x+ZqmV/H7T1kg1k4jO
6KBMXtOkGus5HPURpu3Q4cewBuhOEajIOA0A46drlgHGDzm768/gBKVb1tt1MK9ffYfjxSbHwEUW
RK3mdWAPEMnUqATOv8Ft21PpAFfi6LiNPvpxHoRw4RP/tkvJ4YcsnqWbqBD6VtdZuivGi5qHy3pp
BUPArYcgrLb+toBbcDK6BoR60W/ocM/mjAsLVRrXj3YZkvYCVqxC0m6MAmJX+a9CpvsasvQ/RBef
lLSArnsGpgi2MVv6eJTWCpXE/IuA+IrRecb+Scd57kafnPZdK5FWW763YGL8L/X9C4tv/mH0FZ7I
DElpyA7/9dm5IdO7IxBI0EUgIZObRwqyA+f/3mtR0TqBUeD1NvChQDnzjICMn4wlK1D2xnh3tyan
TgbXzCEuxE2Glo8bLUVjBZYNixdsFlIm6Jspddg1N/kcA0cmWfwnVQvmgaCY5Me2/H1L7Vji295C
IvFRYPQBhdj8ndYQ5oDIFWWJFAwRAe+1SLzc0j8+K2Ppx+Cf4XNepQUwA4YfRfr2sRECtzDvRnai
wxnh1roj65j8bi9grbJjrJx69IT91q2/NCNFaVxnYwP0T7HuAD+TThNi9pBpPDIudsqzk+so0PCe
fL0yvpe/eG1ioSwjuHOPLEV5I++FwYtcouON7nxLsIZCYYTFkDd6wQ3ZE4n1L6T2RkVciDAbSMbN
q2nUnD+lkKH9JzfMi8B54i79HdAG9Dc79HKvBvs0c7UqWwG1U0DrbNwUDG12MGC64id+Jh3gyBR1
3ajwd6R0pxTugC3ukHAk1LTfFpm0HIIzFjb834n99V9vlU1oEa0SI2b5nBCcHjgPLAPmOdzQ2+sx
pxoPdO3Ye5UWnZKLXtmsV4fLRZKvnZluLQA9ZgSQmQnds1ovrpoZJYfUf1eSDj+pxED7kASvq+cE
J+qunIhNY+nOo4bV2NuKiwYhnweNdZi0HnF8DQSAAvX0XAzaSVcMNTt3Zz1gktofRha0zkgSFge0
+oFDvTgq8f56T0KIarYGFgA2LvAP9nfAsPx+rZPrFHFFkjuxIF1zAQPsqU610aCEg1f/nTursH/i
8Yu9i3qik1PXrBFxnDZ4gjncK77wBIHD4Kfrgm/XeX0PLNtjQXf4++J9gJJSz8crJJAYRIFpoRgt
I/NfLnhzmBZfuMPl1cAJkimNA8RYEj1VwvLUToJVeWWSsXAfQwC687HMMbs3kps4rXZNYFxApA/T
zx2sybSPpw5TEv5o0B1BpXomXblr8wTY1K8qENlR0hqvNEXOk82cywLkAYrhKZqsDfIadKdfqIRb
cxYW2da9yZ/1FliWe29C2qNH86eIeOTcNALT7qfAB8nyVcKx2zu1fO2UM+CR533GQubhHbCAQ+Rk
LcqmIAuyZJkf8UjYyXq2rVzPx/gpYsPJO5XnlN184XZPcEsvfblzIssJ5IHiGSepbgFZy9neFaJE
RhazRAVXv+Kxwnf69GKDEZ/HCPLuIaUw/osgLSGXzXvpr65hdxb3wVun/uA0px28y9/T2UrnI0mN
de6fV/0Clcuz6h0ip61JfUIH874Xe/bPzyktE0Ei700QUJuZW3Mk76VMGiO9Sp4s6fGOvJzlvF+/
yVVUNSw08kie7/F09GjcyylyN6JpIt1k2kUnIypr7k8aCS4F+X4GBt8WjN67h5sb18A/dixDHFO3
DJny7UhO6bL2aIP5DR+RySBOfqOhn2EzCv3+tLa1FTuIIQVnyzyWqDLXOUaFWRx/EoK6NNoe92sK
5EDhugWzlMtwKRk2PJm0VCxs9ofe0z47NB6Dh7W16q+x/kN1sSVJskOJY9hdckfiudh0//Mgb4RE
gtMWv0RY5Dh6VGAcXxpvkNY09wg5aPn9JSq4qKE7DzC9/CucMSQXp5RnQ/FjUeOVRdOQXgy4/Zpz
VzHmj0dAaFxfrFt2Qqz0Ddxx7PdWxG6SnsHwHqOHc5QATKO0qqXGn2sP3Y3tCiusCe5HigwDxqK4
MQn4j8cVWnaTL7d/LRNuo7cOdYew0Mtp5bLzTxdKBgdhd/yjwnZh89Zm9HjuPMKFPIY3riOjlyHV
50zAfPqH87FJQ+tkz+ExxTvISamRPHyCoZLXNOWXIK9N5TzxRvoOfFjMmLvisflPYlXzaaH0gwMS
WNVZpBHsxY5In2phSJvsSUNhzrYgHW6tf++1KG2ls1qZoUPlUTNAR+sD78L/2jM04XL4zIfClJaP
CEObk8HlM8HX2A1ToJ8p8ldpqu/YXz5pAlqqr2PUFV/sqlRKUb02gtO/E/qHoSXUy4kt1LoJYb/3
NEO+AQoH65ZvbWwfAFqjo7hzI5U80EeoT7HwDS8isC7gB36PYG/6HJX6ywpKgy5rUtWjKAo/QjNr
3TYa/lKDFYkmgCLD+KYQv3LWLfBKg3ALF1Rj8z/Pr8EcLFAdnK/TYSK2QO+D47KmgYjM0WtJxtbq
vj7ywStVtFlfBvU1mssVKj90H42yeK6xY+wbdU+vY+EmxY35XycihqmeQcNuJSz8Vi280BtWRqyG
tD06FAn12cK1e3p7gpSGCfsjKaWGFqThd6scD8FxmU/mPrdEryhAidxkAEvFGgBithM0oJfgUrm4
SHzoqBfMcjZ3K5kB1fM2+7vpAZjxnLo6KMKN+qf2sQgsoSOc802TcC06A9GUrO0R7pv1DEvUIen+
+ur3gkJS6WpD5qZLUOq1a3En4ny7jCgElmJ5G1yJTxQTD/+cDQ/ip0Gt5E1fY687VDOHmzn0D8oi
lV1nW8CnkUKeiXLhI8K3HjJ6sIF6KqPrOjpR5PKIO3x9ytSL795d+VANzLsjpCTM//Wv1XVsGDG+
fD6APqK8Qo/wxZL9rGo4UNttCaFykq0j/x8PjmGR/kdsAqy/5/K7/LCzS/7St5iSbrTwLmETWPe0
j4aO1yrj1jWa7ErRGVo+rv+L/Ekp9lwVTLQgMSec4aI/4dK7qNJGtYPdORh8A+1vgDnsyWpc/5rj
oDfZWz7Yu09Wl5NBmU0WGWrBuaaRSLN5CWGW+pTMMua3nV7rW5k/7zqnzWFIOoMqfhsU0Q8zNz2y
jgds65+XduxWqwKiFuLua0RG6Hv2uqWPSYaEDtfRmQpY5XVjxjSf6r1pqg5VFXQvyjD8REUo0ffP
W9s5Q2vHTE2CG2Osw74AFgnssblQdy8jIIuk49tgiQOCYIfXVH3A+gBiWCsUULGTp6cxYsmp5egt
VUczg0R4OBOx7ug6uRY8Qm9D9eH4TMQChh5C8xjlUXHeb0d0JKJ/bqHgvegF7UB57SPsTgprLUXB
paN1NW/ApAkV9MKAIaecP8bDcjKDuXdPv0pV6XKnz8YwGMJBZ78stn5PLJE9uCYMQGYi2YyURGCM
DtPgIMSaFAM0g/ekiotV/5iyfjI9i9iKAKqNek7crER1uV0rhxN1H8efhir3rgZevizZrOEnMGqq
VnJU7tr+Qm7HdwiH4p+Du6PP7/KqK6SBi98V7rqGW4t1nyTdTXHtZxjEQjC9AHaqCUrVrqq+meXj
MTzlMvzvuHQ/OMDfgAICY46nZF3loB9M8mfwKL759UvkRCOg87zwlhJJBZrnnzeJjP0V3raSPPMW
5RRLbyHhY1Oh9rkw/Akv4fHe08RR/RshSn1BYMAQX5OC0W6cGz4Z3DCD/xTxtForlXRgXEz8YD8V
ovJ5K/GwrwVSlk1xCGrEartgTObHzLmZfl8Kg2NpsyN/yMNRE21JGjt/bDjZzL3fNnc0EJPzl1S1
ZTkpeOFHKfgJCVU73WuWF7tN9eiR7/dNULcM39UMh5nmUbPEZyOEzUAtP0+eGCr4QIZeJcoXApKP
AorNZoPSp7apGcE6EXv1orL/zmsG8S6UVCRqx5/Tu4//pCivZPX4EqWNCotnm1IG+JxZ3d93P7DA
t/R4+uoFMk+9rqVvh9Uyv5fn+A42wSyv8RXJr0dlYaOMhxuGh3sKpxra3yEWw6V4O4DTH0DsicIK
6la3jM8Qsq9oHZhZ1ub8J0xnQKIIgN90NKGaxNMwaboS1/S6ZX+wQYzDzkRoih0CH7coGPG8KGwb
cgB6AMss2Cv3j5yURvC+VC1ZhUZIzSr5/MOdySOscZA1wg1PzbN0jUbCLYuAH9t/LtjC/RZhJ39w
fgB6pxrrBBUSxwR/txsMGttVfUuTayLU3yrXOUT/6spck/qEvHjSrkCp7Jg1Q49oJiJ6P8zFLLF1
AgTx00frcvbrqaMhuGgjgUBznJSxOX0XBfEcZGGH8APM1nORBSreVN5z/SeTVq1NTYgOu6ahP6mI
k3DtJecjF8cVO1Thy7bTfeM8v2P1+go9urwj4v3Ssxwe3Zuqybolreq6ok0iqPKUKW70dqvIqC+J
l1WSA2zykVc7iLswjcZ6dwhmW/85WTVZ7DleErQcpFEGEmYqnmrfU+6thrZ0vZMJIBN3KZiDh6oV
xI2058vRswXpRT2IGLDeyJGTL9nIo/4bRe8JKznE7sMPM65Jrd2v4VZzpPDNVHAHcgkxEGyIJ48w
W8LFTkVpg0Dm1ysi/VPscpVVFwRaYfDtLYeOHXzkfKCiidSb1mnBcQ0zIuf5N4QEM7fvrHWkM+Gj
DbvtJkHUBY5aYFFA1wqKjkVRRuBZHzVlbWbPhPHIhJE3KNO183I7AH0zcI8oL/yr0z1wh+Ja3B6j
5In5e3YYKUQoEcu/4oo6z8EjFRNuq8cl1hmp8PH60mS5AWc9xzFIY8MQAwH2TNl3fxocQGb0ZP8z
TmWEnAtDoH1mAtk2KqzuBL4jeyO+IRrsV6268EMZsuCJYpweAMTFdlfe1piNVDhj8u5+8pcKlyOb
+Z9PxamNyoLEMvV32P0K/5HGZtXPFVjI0g3NH+9EY2eXUKrgsGaafGC90NdKjPRRIx6PCDOZqDs+
MmjhQZGotj3G071ASSVgok1bpqcgVSgFhqBg+8lY5kl2Nv7KmwQLQUO0MtGZZ94Fb2dv2tFFOrxE
eypRD2ZrVlUTZsl+OQptCsitWcgq5FwPc78TUHYcWTwFZN5HcpNLJrhFWHaNjAwZkWnJi6q3FSCm
72Dxi4IhROXPnIJcx19aaul2dXqmTn20+GQ813+KfXl8BdTsYpyJt0CA5TpV3KkAR8ipNr6scVyT
C1TBw+hQN+NAVxQ5FERKmJqeedOeiTJda39OtJ6Fl5LncuSSC2gVskIRJYMPpC91oU9NuD2o7MI/
2/kCPMXlaUB+wg+SeLprni6G7sqPcElqguOYmYfLeP1xdZpeFPwfBeNmzd1QtMU7ezuzMKq/PVAq
D8ewvkFy8n4lhNCyaTJbBnyKwXrEm5vBm0wZoNUQHHnDJTnLLmC9Fe0gKRNcWbyDd7BE+zTW9Xxu
IE6nE3jOLId+70erl/FiR+eJH/LqifuMRoG8o4I5nvBXeaystuOzarkDwhHDdI9OgCOnHr2TnL4P
JJi+H47GE/4wJNjQorCLmH7setPNXOirIlHw21qVp8eOm+sjkEoUTSl3UN+q9RaDVE00zbwe5ulN
AnAbt6mUY1Vm7PzcNyDJ6mE5rQx7o0Bp6+SV8E7mDDImQ7yzOlvrZfoK730tePyZafsSuAVKSY2H
5Q1VuAc9Z+vTbXtM6X1TFCehijlPiPZ1YCZHIVpt5Gl7h+K3xnQQs0jgqgU2Yli8Orrf1ZwMuf6A
o2oUsHbrFkksJLUZCC7cgyXrz7VlcRtje/rgK2sOGmK9eEopgi8o0wOy9Fjy9l/ofqngJE8yCRVT
QdazoaVobuYalB7K6yE5rt7DND/RruYgmZuFKIYRUryh+PHB2YtLLxCULYRf2qyyUXFYSunz4CZH
2iNIVadVgkKFAXpmdt7K1fK3rqXqOTuz6VbUVXfV7oZos21AjyDSsODx3XklX5r0eByqyu88dxIi
8HGFfcFZG1xNVgq0p/6yRaurUtkXHuwvlc5lImf9T2NgDGERc7w0Jiv0ZoyKFFTM5b0URHKZQy6k
SoLCg0gyw2aPdTzV2rFbyBRCqeYHH3E1EfwRav0d5d6g63kA0oBgv3iFhRQSjG79i9cJqSW96sT+
LNwl5O49/uMibH5/vWfsp4igDSnZjbzbcBB0mnVapudx4YSysxHFGf9Y4pyAEu8YMw03VopfSNUl
Nj9IL/5J8zxLeq53QwqCeW3wgHLXXqUPSfdpLWJlGOZh6tVWJdc6yPn9GcIOXd/EWjdabjX4ZEC3
CaC/Sw4871NbLfXYC4MIM9wBR0QRh4T2J3FEUsBoy9DXOoSUGVuneC1YoH2xfoPOh+lD9ON6ptyc
zN5/KUqupymj2q0skXb3kxFbb+WbWF66LM8SW+IRrWUejkErKlr8AcL2+2S/p9M7Hdr3NqzYTevn
u6Xxld0R8D4BN0EULaRf1UHUhaa80PtqdRGMQP/A260I3gbBGlmizMU5JLlXBOng5uqUHNuKJ6nj
VfL3cOUi4mY1EpwL9KCdWdCyRdxNP9c4ICZEFN/gV+eUvK+EVHCwLpQ0iHJcrJW6GpjlpUyCjb+L
GPf+CWsf5cf7ZJ5Tw5J8n4T13Y8idvW0qY7rOY08r+H4v75xB7GfIjD39HQFPq8+FKoSeDdqBX73
7/wHFycawTkdQ1hMHUuKOmfyDt5hgnmlgZxDkEtvAt2I2JW1pch8XGQQb4d26jel9aapS/tvKgoh
RG67ZpYPSTI7/cxTa7BhkSXGkzkhl+lngBZQNdsAbvVyi0LB1tQUgV38KS160KWFjnoZ17FJsEV1
mEHUqbX/FmfMOdB5MrLT7zqYMHaeCdigiBwOkqLXd+UGQX8PeCV5yjiDcUfsaWICXGdQVK/g8gmv
eAojox68CKhWWkG3pqq1MEb5C114c1e7EQiJwvOUD8IrANDWnrWWqU/tf33NIDDpUXTQd5jTTSHE
5Y2RaBY+bgmAMvr4KOGAQAYyzfpqJRwVgEpOJ5t5EJ5u6QsuDoopf2U/Gji+YEUvfNyFiy+xoBoH
PgcWgRjuFnpqftnL4guxUG/9yCyo2lyRlR2MUxmP2OjqQiUez5IAX0FnCpKXd9J24DrO6P+3LXbK
2h7nxbEM+NCAfq4Qmo8GN/8uQwN8otHaJ3QEU6UbtSa2TFPcHy2DA72+ul3KEE6ChLwW5eKVtaes
DZPDk4p3RrW5+d0w+xz3NbEEE0AmgFpYyEvWTjb6gcbbRKwAMgNgSgBGhbdoVc4J7KeyyuK9KnCD
39ZGbEFTE3LF3j8sG4GBo4Tw/Dw6VqVIjL9pc4Sx4F+GoRv5/Cddj7BeSp73dWKxvA6ryL5qeD0I
O+1eZ4tTlAog309clXWhy3/8CTHwod70sHoYZOV8CptqyE4mshvddFUa/fpzBZYavDJ7yI65QVRD
V6mxg3NViQASmmkAqSIGevX7giNpgHO8o3dg3WFlQw9VT0/3F06uQvqkxIUGovB1NKcJVLl5did/
tdpCD6qmZe2kcT5lyrG2q4SJA1lZJW74H1R/KzhN4B+Mgtj7T/yTFTjCgrYWFyNVG6Nif3ItNLLp
VQ8I0kaRCCSIAsD71U1XKAQbgtKCqH33NK6EJFrmU2mnbyCoNbZNUfJGZpKPK1wFfn+cVXVMRIpa
LlBFHKj63c3oARIZpUaP7dBaNvQIUBMFyCPC5Cl2tMl82cbHNtABpfEhhZ2tgPEg1AfdbJGTTqI0
GLuIxzPRqTuFn3NMF768s+QAaUbXbV0WFrX5xVj4QqdB6hNpCN2RrMnhUWXTRXQU6kFl7/H8fVdJ
2JlIGThhYFhk1ZHftT3aEay0mcQTfDVssDpDUSfasRmH1xVY0uWEeiyIyFtNdpKy/7FFHLMpwVIY
p+EV76fiHsc01UmOcu6tsydQfUIYVNAEULGMFlHGC7zJHxCb6Y0CGwdsQ4lhUSmkq8yuZFlVcrW0
sRy2oK/uHJgMCR0xKt1CM9FDTktg+mcFdVDUt/XcnhcG1x9IEBG+y2QFcJU3J44irCthUVhQ1+hH
Hz3i7mFMxmu4JYS+NyDnipXLyqjaEZB+INzfGj5T4qFcYTwW4PRon6XFciLtJwGnaOpzdTsTYN6n
g8gfrSJqa6hS62UessAV0PlrOUYv1wc1j4vJNkGjCYmpr6keTuGhXui/hvpEeBxvXf/uuZ73v7rl
i+ME3xR39W+WLgaGRC5xYCbP5vVfvggl+37d9fuGfzIqvYWKnXqtEB2x2PFh8rLgI668Y1iy1IhS
GtwvB6mLjHK30CTSCq8fHrcRCn8mUeHBDOvhnX8i+OCX5Nlmx5jYiEqlpxgZwhooOjxhun3pDK90
jSH9TZbLhNcS9P0l9iB8ZP6kr0TY1XbhB8Ta6Q1bSbW7H8A6jkFIbFtejyuuGt6KoGLv+c6j3Rmc
syuCxVhHqyg+vvSTK/oV8i1oxCgT0ihYiRUwsJ4swJEJKE/3Mqny7Hu8UzrSpeSSHjjlJ/Nzg9dg
7/FyhwPyHP9mLSnkw7A2xuqZvzNQDPp23xgc4E1UKCIS+xzzVTbxoSjM2HKADVqBcJRikWDlTDdq
HMKYPccadqYWRoWCtVehZiWszjgwg8TWb85zoyqBXfQKUH1zwEiuhCGy+a/vxHlGJjwuTe+7Vbjy
lumxMW/qaf5bt09CI/Sg7nguOJb8OHrP9pnN1We5EhoYN+VovwBfrFiAlchq3DIfFsQocpFBNu8B
128AZm1sOWYZQAwV/7m/qS21nhgtgeYwOaCkpGKkVEAnJb0pGhRQ6qZgL68XXoP+DwcqowabBMch
MbGbU/gUHi/yNs2r5/PepfsKN1lTpfBqNGjzOFXW8YhQZOX3pQj0rehb6rChnkwpbmVYOvRDewgI
5KcuxzDYg1qDjA5EJRJGoA6y6YLE9+eQ7A0eMJ/3eN7HajNa9qh1N3etyIau9vkVa5UAklSvwuda
ZJXSNjrm1NR5GeOT96SuVl0CKFe1mhOA4Sh84GHflMMqI51FbRSajOowHjU8VmMxkJ/lRHCHMTWy
1OP2QZXTOkE6zaLbrPCB8Woi0rtT0mm2xfDqe7jcWRX1LhcZb2Ko9sFm+X7QUlUK4hSkiWqq/VAk
0QbRKGdw+tmxmLbJ0wfxuijDNBlUDrtyzEj4d+8iu4AOyX9EB6kkV8kSr1geFFnmqlTKF6Rrcd1z
ZMGEtYE1oTNX8+3zrq9Oi/nAvC9tS4bya2Gwf0mLnpWvUd72MFlFLqE4PWMrtNMT9Hs51sf9iBXD
FM5xkyTb/pYxD8wxR+b5iCY6kTNiQO845li/Wu5UzwU85+KiKHLIfWWt8hqANSyZIgcjEhZnLvba
KCPthfY4hISQt713W9RozZJUQMjMDMa2WP4Hw9wqP0tNMf5wjIRD+N7HMejr9napyrst0dECmaBR
zOPL0fjuXa3pVQ2o7eHUexLZ7DSNZu6GXjgawSX7RDaZy54UDUU7tfADUVAMW1I4xENf2GV1wyqI
ULkPqvC7uHqFrdJTlm2pAlIHg6vNbqibNRXt6lS4HgoJ9ZeptKZi4pkqwDPadbAvr8XNBnE/9Nmn
Mi1rcT/BhKfznqO7hAqAovhIIzcKlCAdDc7BENKHfLKWxmpUTFhflm2zYkMIzu5JZCLrQk+FTSQ2
VUCyoEVsmBCtQDT8M7mxm7b9zkC9I81bMweq5rVTKVnRHoKpzNPBaPf2/RIc5gkYsMYq5HNDqd2Q
kLe2NUkIKKuTPOBrpFwTq6qUcgE/n1z0mq9LEqg+C1zbN/2+LFs+ewDJjER8gp1jNHEG3/RbPg50
KL5D8iCGXetSUrk0l/bzMUnoIg2aQBPJlwJpsOQlVr/o/35Qmf33L9NjUdYnKfP1fjT2IwHbMjPC
t+f8cj9dbvZV+OFvioeO7p5AJBzCwLwEoi5LmOQIbaE0i9ySUoM0j7qjinE6ORzNzAwvLhfB7fty
+RXE9U3P1hlyQJ5D0+DCA7K0bXtiFLnUQsmsPO7pHZbOxPIVKD7nxTJwIsL42zJrYprawNV1g/sm
STDDvfexiUX0xE9moVpfFCykOm+thskHm3rJBwqZ1cWEDt56wJdzFrig0Vb6GT7AHUZ6YKnDxNWA
cCVAo7GVkiCE951oYmFbvlaGxhVULNcj2hpJ6VqRzRw/ycVDs6dmFOs2FxGaYdR4ey0N5tE4hBiv
yAXxYtYJWyLyHcGH9i1TO2tjVteTdjxVeiflym5su7b93R6Ki+3mbccRJlpCaW4fdp1KoqTThEFm
QB6dmpjFMADQgIxqZVJ39mK+DhtL/Vh1/hAmtu/zqDBTEpg9B6ZTWdJkpO26+XVoUXmRmvDFSuLk
gnbUDabAy7Sw5RkFYnY3F007IRauPj/0UJOMPkpWEWSVtOc5ZXLtVpohlWHXH6m7PLySiu44bfql
Uuk5k7vi4A9Hgng4ibBgXOyKVYvOzUEMDhoQwgyCJrPs38jlLveFTtRJvyWEOeq7Az7n4aBJwNnv
4R5S3blArobXP1OdnUVfskKxAH+akeXa4Op/O7bnklxZoOXy429uDl7WB8DilbvtxneXtN2yAnnZ
TmeOLIDiBbHJ6OIkCPfnUsDj5efyTaCfVrv4Iwi5h/KttHyvLqClyVhcrDPQbOCidXYdMvdxxTNG
mAV3SJqVNcrvyCjflypHUZAuMw/1xCFhiIVJvs3h4Wah7cw13hMLBhYKwslYE2GqkHN5/fBmTfla
5ohk2/S9MpyxcS6Q7dcCv7wOwVGuvsL1uz3izpPlxWgoCzTxM42us2YfAqRA6nmbKbJaBlx+3EMa
X152KFI/hGn8pbvSawnvQxPacx/hpRjzd/nTr6jJ3dIllXVypvTs357TPH6fKLXeBwN76WIzlHtN
FoSDuaYRa3KI/cYriVsUjjf8bpY9Mu8O1ELYwhudCPfDu9W+y7SdSBzCpBkc+n0lVvi+6ks9hgoC
C0imKs2jOuX0B8/eZ7Sgx4uUr91npsF5Yc6uwek6+DEzhEFkkHijssTIrqMFA30WfQ8LV1ghjaCW
YC+FUSjH8A0EO+fGvDrxFPZt2hBLnUbyvyhZFK7d8UkDyGbECDAcw4ZiMEVSL3gJE8xnCKHNgQKi
oLPv16sfkj8lHhkmFGV2pS2ROUVRy2sTqtpqQmJBPaRAglH3RF5nx1Z/b2hjHsK9kJFOsxQolohi
KbbN6CsvpWjsyklTldjJNDxM9ESluy3YFxJg/6ctVC3VBZSn9SjCCeiRCeZytdA3ITnV5DLEoHqU
35boA1wBceQHq2G/k5tcx9ERCVpvZkc/5xz/1kz1iqaOxoOBOVxri64RgeRcvcWIZpKk1aKYL+hN
BNdXG//y5Xo8jattFEf8mt94T/HCjNm9BpxSCrFBe0u1SSfw4mlf6nCswyDrpujdf4F0o4pDAB70
Qs9d/l7ID48faxoHiv97cyEKDUDY8f0lkokR714hzSolil66nLYcsAZsQCnuBhrem1f7Xb6H1J5y
A4xX7MfbNVdsrCnrKw4bFZixOTML8ZzpwoilZPzz6czlRihEHZ57VlyJlphkWcBMtjQQViuFX54P
dpPDzRpEkkg3McIEPS7dq94nHPlRd8uEFDV3AvB+1ajk+63fSoBY7ZDS1wmV2ofHjxXE1bDtLovQ
zI+OjIVfVj7uLq8boz3BGSAdqEY+WGpjlOvP78ZCUTIgisP1c1pd7F/4Qpu4vgVa5PaKWJCn5/Tp
lup8tIyfrCmI/Cg/suu3UrAP6oOQ1+All/UayO0QywUNb8gPDBw2SXi4jnum632T5bo6I5QqemYf
CIyCawRtX2gd63NZv9FflDR1KmPUxud4B6ej1Ae+N6N2BP+xsT69RaM8SGSlrfbYtTJgZb2v/tLR
Z5bIZY4BWrkTkUhbS5mxw2oUUyM+65VE20j9YOUPtNWRyyfxGLnr6fba+K9LkGApi/IMFJk1ylMn
qPrO00xaZSKi6ykz8egvKaGPxnl+V8VtPv8sAmTDCRdUw4Nck5TGpYAqnQBLe4H6EmR2nYqoM/gj
P2wd+RUT1uwNQIKf3NvhTDxzXnjBTceA5QIUSPtH/6lD0RBaDfdjIEwz3VoDaVPq9XnnMBbQ6OhL
ijWQ4pYrnYuPJSHjNMzfI3UEfkRp90d2zINjihY4XrS679ra5q7nIciZoJREjj8kw4HWgK7CaCZL
9zToUGHMGFFFg3HYVhGDh1GOTduf2UYhZRe9Nng2DHJq9Jlm3Wz4ov+O7iNWkswS+pzfcvZ006EA
/W/2WX3MIGv903OkK60PErN6e/1astj7DLK/HGpMvOOSOykX6kaxDJV7l3uPUmnXTHDPgtv9aBpK
RVFP6hOaDbKZGvIecorGhJKgyZn4/dvzIQWtzxOWqO58bnwXLwhlUuGTf0th9p+CkJT9yufUwZEp
KDHOnRJ7J391tFRAJQrnjBX5sjAGJj5j9ZgJc3935qEpvPKXRakTfXMYnGitNmPtSRlAL/5uBPv/
pLWmiQ5fOyt4AMg3jw3yX7+49rlhLlxDsWJSVfEJmF9/2HoqhVBL9MAe1BIun2wousvCmQmbTMGw
b0oS0EL/LEuD7Stsn2k+IrJ8PYdgHD1oVhaBiEuZ68QGq72c3n27NZWp9ptrXmz+RL1OT6Epl3t8
bLUIMAei5FofYK9lLXPVLdlQ3cyOCOhUTs1sIKG+kR9OvBlEoxL4RWPm//K4ZzHN/ddYs8boNZEw
0BvF+ckiRg1VJHW+Nve9TW/ubuRNnTUFG8VqLZEGEED7e2KdkpZsr5Y8yVTNjhWVgGjrxMvOLQi0
9ly3gl9Qq5bV2mq5RjECje22ym+2DGRt6+Waj3vQaI3ryM+re77cPAnYqgVjUdRitiqxloYlxhhl
S1QIdV8IVpDuWswbj36n6FO6uUAjJ1K83zWpIF6/LsUMDZdrjsMBnkjmXO4wjmDHYHv2C3a58+tM
OPzI742wO4EY/DTX0xnlyWRErEFcCrfDlZBh0udD//svazzjFhp0imMUv6jx6NjcktneLmWE9IFU
XqLsyrkG4/kst7FN7K/AaGxDTH+jV3TPnLr4g+MME5q2zYFajSIlkOe91pO1VHPRfbA1agANoPfa
azFliyeoTeVSX3he4JultsMJydOdDCYvucI8juQWAfiko3PnB5Akd3M+X5UvQ2Z0P9NWnnBdM9j1
sAVtIK0HxhZEAlcDvqcJkm3cbF33ievjukQfX+EyEEzWRc1qP/7UJ+3G9mjGrbgBdlgeVQsfwBPJ
LVhfGtEy0T0ulSbDjeyWsBRqt64VIaARoj0CJG0Krqhf1i98KXAIXZQNHt11vHy7bgXALGdf6+Dy
OqJob/ppOXSsHYlY0jsSx5RNJUM5DGZCpLxC8HdxH78UPhM5xkW5UCjghvg45pQdylCeHKRdJckQ
BSX4Z9AdFhTX6PTxlsYkmGWZyG9E8SpjNtOwPtK0nnfy0EQgfGmnRN1DGoPJz9iJGmgqWy+yWzyu
EYTPNNFTLC/Rl7IptCxGytd/ChuxDnFFGfFjs0gUWDCOwS6Nd8MedDPdNq+1wYgVKnykL+f37gwG
ryDDI9E82+3+aZ2iMWxwYr8MLFZWzwTLHwP7w3y6kVY7rn+gAm1YcFG89RP9IJslNLHbVzdpxspb
WqGXCzqM3YBHu4NuFBDx/W+dxTSxZft7K15LekymmeBOrXp6bSVjg+P1U0C/NTUF5N+dfOveIha5
SSw3bCvFIp+h85axRG8SPOfMABfhwjWCGUZ20n1sbumY3Gm9fmo15PhF0geumoKiJKdloReelqIG
UmheVV8SfJn5UIpdzdKRRo+qOO4rcLU9vW8iQH6MUoMXu6nFoeVOBB9SpfTWzbtpfnOrcvLFsGkh
EIHilOxB/MBqaX6C0USy9qVOGlai1fecgV07rHDbB5HStA6IrEkbNj0TCfvL7x6DpDBLDBKGucwG
XudE5oOUe0gXjPCTFdO3Lut/Hyy6WqX422HlOxL5G0FptPAvZ4XS+8VXl+VI5dUWosUMK3mmdCAL
oNvNkYgJcHUjlBCD/XPQz1t6G8Zn4MjNx7zE9QnV58EG1p+bCvlD0sVJ5hwrBcp4JzDGmQUbzTHZ
sDdFGugP0iBZFElSQKiElK2yci3MvqCfHMwTg2GDYAhP83VlFHF3nlin/v6GQD1WQz5ZxpOgKzck
JI3fU34OvAXdWwI6gnznr5EvnjpxgmZD/WhJqkqoeCc1KHMF29zlO2wIoUEZ+mrvA0SHScwCAHUr
a07ZdayWpnWXHtoQItMFi+QkN0byNt86gJjfqRCugqTOQbOmS7YS1iHYXWP+ORmJFXuk0p3qy1XL
2MwnqwD5UZe8ycZptpgkl84zn8qkiRUF+boq50LoAGTdmDDGeZWtO1TKVN1x8KP/tmrroCZUXTHB
SypmVLxX6B9UDdHOapUDxfBxho2oHkrJVmuDQYtFrBs2Wa+r/xHYMEW3tQF0TBLQI/xuSiTvWGJ2
hekrsak0rW/6Xk/xyQ7EUwBZoC24WBpyDlcy26jXWVlNAWQHHw9jgTEcrPUU3lgY+VUf2zze5puB
1oSLUGpjqYPIexZsglGovZT6Mesy9+pR5loCDy20a+21ANUlEqHvTebkesDpRNJFSrUm/pPXmZ/H
GceYZcS1YirjWOycr//sZjDcz/GQUbbh6++HZBvLIBCOD6Co30HsstTOwrotY9YQ5PcMNHx1pUIT
d0L+kOEegvKm1CJgybdTdlcg1Yn7VtOdYkV11C1rT3SpB9Pifzly8/Z9cGhc25KG0qf4Kwu+sbQz
8a7KcZyfG69ODueULDTr4W5hqpSEEjpoGIM5MXXtBVZ+aERCrnm+tInDNXQZANc0CUOCtjYY0ZWP
FI/INpnXUwrBexoMVy//F1j9V2VfC9eDM6kRJItwqP97W+UwE6gD8YLzc/uCO928GsW62H852sK4
5umsvGejmGf7+Q4ppDVGJAo4jSsVue+XayQdpUyG3GfOuQWxL0AYTkQtmZNZdj7ZPR0sbwACaYxB
wwv47IJUPw8r43mkMT854JTj6Vyed6+1GzBYaxGNUcZqnSGTHfWbnA7sEE3MRY+IGLmJZPOHlHej
zyc915kXpO/m8w/bYP6gGjgnaF1d6zmEpLcBUB7FM+xzn8lxxi9LoAwZEYQuReEIYKKeKMufFgR5
ie45AIL7uL35DGurECwBpSFCaReIiHqBhNW0s2k5y7rF47ePa1NngpH8xWDZUFGb4Z9o+aeYZkGx
FsmKZWgznFhk9NWrtxU5jbu7ODSGo82aW+ox8GU76fVec5Ce80GyizarWu29acX0gwFAhFsU+mzI
i9f7DUyZzew3xnWnqpUMBkUYpsIx734ohboGD5rk2CQdY2IbMmyTRZdyN5SkpYd/kmtz2ksMKMeb
ZjIZ1lwsiq5arS9UQpiVvxZoLHEJ1acF45dJKmZb/30ytWdbU00oRfd1uPbjN/9kVzibRKOB5oYi
2iUS1dhMxmm1/pKI4KMi7zpvqVmycDc26cCoFfwiU8ezi0Fv6DKIb8ks1YlM20pJkHe82wzU+0jw
GjeUlxe5vruoBYYghl+1mJ8y3n+sAjAeWzH1JDXcOnb5DQFsWn6wSgG9wKYEsflNBlKkcPeGfp91
7+7APUe+M3hTyKbFK9lszgybJlYKHq7lOphoatoE1otmrNymR8Dw7EnaEJaynnRMXG4h0TPoA4Fu
Vo5U23bmW3hTU//lfg2gbjiRdzPxiHMB/M8GpPct2bKRiObrLUOW9Ni2z5+i8KAhKrt6hKsSwZ2t
XFQ/rz6ttlu7lNeM8bVnXpJHo5o4Vh+ndcFl8RvoKJ9CAx1E4PycSMgmxVyH9+u7tLe+6jZofEAZ
0zdabzbp3OjJ7EH+leZMQLddcI3EhsmZ83HBXEDjkMocAD67IqsotCDyiMOXl3ASEZThFBMpqb9l
igKTrtDDi779hGgV84s3SVh2aG4PR+azu5pny7DD7L9gS401Qm3BuEYiK+6Rfuu1+IuNrX1zMhkG
Ns9Q+Abxr+Fy7PwXtyjHwPSIDjDE6hB08oPtfDvsjNl2Q6pkaxqAwCJetmuz3ecoTOOA+bIEpx5/
7ooaOmQNd5Ar+OepC7+IfEz5x/T8ZjvZIy2JMLQl6fMSL1oiFqBixY+2sC0OoZkMg9dmTNmtXvAZ
Z+/5hgO+30nK9kjKyucuyPPOLvD/cPw6WP1tELUVYVXbgrVF1v1KdIlzdzuAszFonLKJikua6Ruf
95/yVL8tLb1rX/t2mHr+tf7I/+1lwJuF+YZBc14+f0Q+wQNCDsf/JxemhndiXjpoNmEOjS+mbbm3
J5Rx77vbWSWY/Zg0creLtq3MmFq+hEd2NqZvMohSR8FVpBCi/BMY70fLqAV8ObiSmkuNkbUiSH2+
LNJFRkIeQ/XW5i6MCKcr4BdyeXYvezEecKkOaoxQ55y+riavVds8gotdgR49PTb2oFmfAmaoh8Z8
PGYrlB8/54s6gcBLwHUhEc9TT49yzLJOoYsbkBveqaYhQTHEkRO8oDj7TOFEv7NgzAoOcGNuJUvG
rU6h7w2VV+d5GlUziq3q16F/HLpIWkAg6eHFSx2xsC0vU1NxZWY1MKeFRaDL610ir7ThTQm13fSW
9eLNTvekNaDNYyHGQZ0+GLsUXujtHRO22t8LFUsn1CY8R5hMI3Uy6/lHesmLeZSD/6i1GZ05lKT0
5wFF4+/EoaS7x0Tqysq8a2WrnooJzFnufnngWGCcG0F6rgXhGWt+J/SJ3eMVopiqT6hBJ0T13tuf
dRFS+Yd19bwtjK5v1SkS2UkNsVmt8liNmBS6VLvTYKbx/rPmR0Fe+xekgS/GWUm1YMFzxOKe2WFB
Zxkdo3LsEHQQNFIC04dMhJCs5hGWZ6ptQ+d6UJI7plGthR12kZcSUHzmEDZ994jX+9glqJqyP+G8
ATHm1tCY8JR3WwWkduEZj9PzGzVKo+Dsr27BgLQbizmO0fs1TOi5FEDYOgroNtJFxMa62K3nu69p
+ctuI96tvavP9GWVrcYtYe1+iJ42CY6gVvjZjE1hxL48fzvYMBQyS8jckcDfd3fVH0SPtW/8UH7S
3TGe4HG/JdlEuWO7hm6CQh1PvHu6VxUpQ6wk/EoPJr69Dd/hmX+YbGpms2+V9sULihlFRW59OiTb
t03hVX33ZjxYPCC3pDGdvF7dvhrkYTw5DwyOJdACPsge0bmYH1P5UNPxNcT1BVOSYYyLUy6Ryub8
ZEcYYsXLMBKpZ9w31SuOMqY7rVhv0bd4jXnV+/CCBPwbP4CQu1ID3NO1NaWKG3bHlpWzofuo1rlV
FZgBqwX1rx4599xD4Ch1HQ3cDbczsBNKNR58lnAL9mrIZd18yjI44Rg9luWA7WkDtQjOTe2ah7xb
tjrYO2YxuqTkguboN0/Cmtsb+QkJRLNz+bcIqxA6UY9YjneuSC7T7adaiBM5WHYY274g5rgo2LCh
C0+pXHYZ6EWya2hOUPAeHOWoFoDOUWC0RQYSHPx9sPnSD/tTnMAOVEF6QRCnhkYkQ2GkfReqwvis
aCUEkrhC0zs2fnTbS5qUrRLWa0VwbjvltUCqvMwsHO0ujsDITb9Bc2gawsYG5AgwmOj13fEm8mRy
zgDOF4eKFKNmGa6n0eJD1/3UcC/BzdRp9TD5rHd2buZXMi6+j/y739C9li9mhnneiP1RRduz+dk7
4kf5N8opNbAShg2DjNlDyyPgwD0v7WsllUGzmnd+UIn5xYxz/uYwzhXGWoQJIe/9JCqGZHfl01L3
NJKupJVGFE7cC7sL2MaLtW0ty5pqTwYXiDadOoWxwpcRabUO50ud4IzwLzc7gI+LebdqPtW5wnRd
cX0F9kz84Es+Mf9vg0GSa5ZGzDBb9xNpIW3sf1RLeFoCmADzrltUHsJIOjE7p8YZ8YKe/b/PAjZc
f+SK4mcufhyGeFJVds292056X9EfzrLj0zhW9jbfZk5iCzXZ/d0Km5HMAEKhznYErOSHA63Ccdjo
Wb1THwxmayvaK7hHfEk7ortQp+ha1mY0xWN1g5QIOT6hO8DaEsCrNAkVIQN29nkTFWHSr16CF/oF
EE6Uhyo2gyI53V0o8moQ2W2Cm+FpQXZtoKUsHzI449VPvHb3jULCdYHZ0584E/jBDt/bklMsNpI1
VjXqv6YSEJtXeoftzgMhJy/7GexOoh+33rhGyCms6ux/Thtarjs/iRRE7wFdTwjoGKpD05ulsgOc
glHptHJ60sKI7OMuxkJP3K9pSaNPC9052LmN/3FJyv3FGIqXRuDwyMfmYCY7ySp8kc3cSlXAkhuk
KHzM5GVLDdQvBX+h7fFRG9AgsJyyiykjQ5Kv+MpFgQd+CEsCTRRvnAsOI7WoNlpngtGeL16R1ot9
gYDkS4p+XrgXYd72d4IRj4cAOEbc1uEvUZQNlmmg6oiTgtDY5TsXivyxUdJzpbBWJV5VAuewNDtH
M5DacJBBB9eT3kBe02xiixqxM2B8CZ0xkE9k14os1HsoorUpnb/7j6SW1SGm3dp+HAArOFiFKzhy
Q4v4iIqGhWNXVtCABc1iJHAZ/9FwxF1CmNx703IIN5lNmATMhDixYBLC5te8l2qWqmbVPBTEer1q
1emz/9B++uw/DzPtI7hJB/iVbCREfX0tPjwk8L9Kwsg18WLaoreHtyfSYjiqO6c0qlDdae9EQiSD
q0WXubu4PAag3AN1Eg3nBwPqzhQxMLk9WIJLVWeGqsnhUmsgmbXoVPMQdKaYKjgNk+4QF5ZCW5ma
pZGquuwnOzECM+PMAydN3bvgy8pprXbCAZnwwsDnEG1D+hDy8q0yoKuCO2EKrt+fl2MShuyX3a4Y
jctgjOGMddaeTyIMiR9b39OTDivqGVzS9cdCKiUhZfeHkJwu1uSMc4nk3vH2pRLcnlyWYFyEMvKy
0zGDYFtcVlgVt4vLGjdZ7oZ/+OSd8F2C5lxglnAJ6p/W/EMwxacBXWKTmWm61BXmSPmIe4GMyipW
Xolr3DyROIf6LhXL6Qn6Z74LZ03a/rMIVFF4Tcq0LhBgmD/JdpORG8snou1O6xPY3q2KiXbBfYbm
bFeJk94QQujJu8GuMOM1RF82pf4l/mXSHB+nrs68hKts6MI46UIBUfTrA173pvkde4rBOFR2zsZl
X8evQnlmAekZCtNkAchcrdVjI7PuPdzgBs7uP0vDqteLFZiJcqdZmLC4wAQ7THceueHjjV+0U/FS
qALtrYeRLcpCgyMbV16JdLvbO4gRP3G18enrV9phMPT56JsUMMzkDfgIKFCOI7aOsJ4DsiEFa/t3
0mQMLTuaC4btBWL2I14NFXkQMnCJmM5P6wB1GJcVjTOHalijYE5ORa4Lm7NHLoCnNT8xZbG1M1xx
Cd8zWk+VNBVxAkiKaoC10OHQgPXjOZOuJXbogub3VdO7C9HLMFO7mAN8bQPvbagb6rENJWkK4L3w
ERd0j4fOBNY/zMJW0lXBRQeyYYeSiV3JTHFo2rmNuz8PYegr/JiRlH9fkpc7inpUAAmPBN9/Ape/
0PEhqeG7MyZwFG9tAr+XxvgZcMd/kG6nitpkp1L5Qa3yzbV2BVENnm4+d0Y/XVpmbEeE/FQTE4Al
HuQeTIKByL4+3lTnF5xxrPr9kCD+bEpJ291nJX3yuXYwIcYtArzQxquk7b1mIvkiLYvfyFIPShuI
coicWetgVadDZlL66PUHWj7++o9STjPtR521GAg/a/xey7u/q7kgwtfw666gTI7tmzU1glPey3Vp
fO1xYeBR4mwiNRPOLka5gL5wbb5pOYTeysFh3fVYCp95aXMv7sKfUctqhL1Q78OPcHm6e24ve38d
ASYBYYVf2xa37EMpwOl5hwb7/Rkzdhy2iU9RxURvXqy0nBZ5hjs3ijTrbzYTdKjLTwk6JOlZlx51
j6ATHMCphpeVwKwtcEN6WtRIvliE+uxNWuRzF00wHWRw1uc0olZLjlmuhIEA0o1eHxkq/2k1rAaN
wH24xltihdBQZAjQnM21I5BL3MuKkPCuX9QGMV+udc1OoGVIEz3HJmxqYirxWGjuKCHNRunBPxg/
xulltv3h8wwUJGZU6fhWLB6DSYuP05FCj2mFeQz0D59awKOCFtD85pSNYnSqYH5UB/Ytxbe2A2F5
TTrPueWZa4+/bjXJP+31vcxMxFRAR7tr12erxRVWb+PAkaBUQEnb1e442SLgZq9KiFGgFu/JBDVy
nKsnlEmWpMRiwb/aZcj4FQrYjO0QigXIcn1E7LLRy/cdx1vsAIvKmoGMI+/OapFUl6Q5csnIJ+WQ
+/R4xDYnRTk2rBsBDei9zV6dEDdESvBp/0lwV0ZRCmbAb1rMt/Fhd3IOE1mHVSeMS7EhiAa+s1Qn
aO/RGfI6KqgS4o0EVOsxaqU/upzgUC4A+H3NNQm3U4thtdVJ6HQSfste0xccOowh6KtR0bzavqDu
YstCMHmrrnqmtwWF4fJLbNc7H0jA/IYv6vdyi4pGMSQqKueX2TYd4/Q6jrEK2G0OsfMlH6HZqAfk
xbnrBH/qoP3Ifj/gN6tkumbu81DwypUguohu8rY9KSMnX01FxGzR8b2z0jrgE5AAh2lbt0HRslLi
urfF9nMYpdedd21TZ7va7K2fonaYScJS1ucjziACQBUcj+iUAjZM0Y4A544isgyDx+fcrOMT3OYW
EtcaLXpTK4WMEMFeZc/9K3v6rwwHCDhJecvvZt+Be7Te6081hEFJukSLN0/ki5Fw60HsfKy9YEnp
YfLcNWH3Lb7g2c8IloYeUGCKR/IQICMgrrDxNJzpASqoj6i0GU57uwj5YVH7d/X96fgPZCY4d3fI
IgnJIX3dP0WjK3GIm0lL+tMdtJgyJCdBA6rpMY8tmsQJcY7bB5saZihpW/LJcXdnOsFv40cw7Yyu
YNi2ywPG9Apw1BloPsTotRM/eCBw8XZERCbuCks1BYqbTjWGdvfDhA3gt1zANchTq22cWoyLU5Cu
1O2RrRjo45gIKV7fmywSLxaVMogM7dxjn0Z4P1FEygKUk37tvftbPe3x9cKuF1qPHn6Keh5P2I5K
9fRx+sTjULjgxkuVLYe/2xSIiRbhp4MDkH2PdwIsGXdurAdSDyyA5nQSG7Doo8ZM9i7Mt8QjAmFC
7m2rEvmaf0rXbGnqmm6A2Nl6NjtmQHwmBsDF+V4AjBsc9vr96Bk5HQkAtbsUuG1kDw2fbbA7dpBa
ZD7XoHsZhK7TkDRar/OQREmeX45R07qFiIBQS0POXS0jlfyTWiYBbinYcjWslwUKJejmizFImmSV
v4B6GOCkC+hlKIld2t09Rq/JFw1HTuH+KA5dLC+nShkv4TfvQuGsEK4Lzya4lHDkRZW5IWAUKZRB
Np+hj1UYsXMkSz0h+BOUZRxXj+72eBX2Y5dtE/Z9IykYqcbbWleClPbFQWG+i7zjRbAU1QWMR/Z0
mDR5RcLQgYFgB63+a3urhr/Eem19Ih5iMu3JDDG8zypUkKUU3UX63maitETtOr1w5maHsm+2Lg2H
0sKg9C+RJI/0/UceNcs93s04PLwGyWKkk09S8YD9ybVF5N1SmbVAy4FVubBHquplqnEOdLvvgRc1
ZYi/eXY9UAu2g/M5UlhnPA+tr6ErMys0eDEPISpgfVKHJkVMyHGratQdUeDBqKnRTDDy6oV2KXWP
Mxnn7y085/ON4XZqJbi8WouoZ/hs5Vqdxevst60pWDGWay0GQjSNarRrxGijq1zTZqwlWUS+KA5Z
lqb67FtbFfvdu3TK+9jQwunrE0BOUyVW09LI2/pIJAD3znNxOXhg0FDYnOzO6q+v/FDj5q/Ivz33
WHDsOVUVIcoXD3ssW9Op/fLcHWzYxso8T+W8K4N/aE32KABxweUpPRjm/N6z3cgDL8ckry2u/T7n
J+ugculRfrIw91K6ui5JJMRPZCKxvJNOnnSuJXB91wxIRK3OygxK5qDKNV4Oq8oBs+tLQlfQzg91
ZdDXT8NN8fZCwikUECHymSQenK7uYASqZ3dNEgyeXJzpvritlvyIt+NiOAJqDHU0Iai9+Pouv7Rm
pyagczqvaGzoNTXfXvk5H9NPeHBQJBmg2dVNJQgk3fD8cYLZBiBZDjYXAgzY9OBawbO6SxXFGiIV
IuNOVA+g2z7SR+W0bhUFifxd0LAV2FqjzRevfUG9Nk49XbkJt7XHabuKveypw5nUoyoPiPu3u1Lu
HTQDnzfutpkK6VDAiMa1JpJdb3CR7opNL+E5UtXMLfK+Cl1l/1NxD0Tu5ECjYIvY68XDqVxoCdVk
Hxp04xqtBlEB8x0n9RP9gGPr4r6thD7hcY0aDwNBm4o6O36mPqwkDI01rrlpmnupp3a9ZIsXHhSI
hbmnzztgYSfTAMfvncfTJYxxD8Tme7Zh526OE8xBP6altKHgTEB0wHZPbIV+tqFk/DCe0zRvgTv0
Tl+BWHLKMjJTHck/d7ACjWK6sdm9PoTDu4iehmSGkFx5XGQPSjTYw64F8zPZ+koaXwGgijpWzRmz
qZnVyX9lV+rHUG25zOtmlcd1XqB4rgrSRJt/2WusTwSqjLCDo1kcYGn6b7Zj+0cWJFV+5+GI+5pW
GOb3MU6H0OTirTz3IH/MM8dZJ+D6gTcaoz76hjISG4nrjETa3hm7iVcSMd5FBcu3WvN0yTEsLTl3
JNKcAZKvRRg3V3DEp3NjYNRwDG8YFTXALa1Sr+0JyFVCd62UBfDy5EuQEoD56mdcrnMRenukwp+E
4Y+P+7uncdyHMIQRpAGvLd/DB4qiZTkmAxTJVula490/Uk7S6pKKyltgb7Eoftx6Z7UWvCp6fP0y
dMmQUuG37H5N0iXcNV+w4TmL76jSm8Wu+LT2n9yoxuPqbLP5EvPQSivCEG974iqtUQ5iUZnGM/JI
AqlLTk4jXNpoXgfJ1/MhtYSWty9Tl9hV9RTStJMJThO19tRKJTAqmui465SpSt45gJOTeGTHbibT
HuhxLiw4rLtB6aW5G+KUudGGT+D598MiwrHofhBEUgaGwhDJv5cehF5tpc1Fs5888YXSU8TdS+R8
tyKeEKeGcqMlnUX2AXKEDrmBcjEOX6ozSEIv/5VzdqqqooEBf6W11oKf3sraTn1ZEZ2ImGrH5Hb3
2bAb22i4XTH1umreH9viXBOfGHKhJ6RbkkhVgG5qmPT3d1YAv6svBDNhqp8hrXPEhWuTdz6xoHL3
EjCg6ZQiLQC9VR00e96jUv0n6lx5KtFoNIbMD3LYn+ezM6JVbKOXU5SAaKPCR3Ke9vVQ48VEY/iH
3Mng3d8dRYBssMF50Dx4WFEXEQ1vYa04sU4mJPHU3mBIBxXOboqqgUidRBuwcCsFAI6klPAUll22
FIE1YoXeGf503wOuwZl1uAeKrVIFYwEB526yCVFCh9OUlmypiSLrPv2PWCIOR3/4D9bTooOFghQb
VQ0vACVs/GHhaxQjq7WwI91DSfOBMKYZQSgZ7V92C1dPQB+WXRJCOgIoXOQKOBywoLYzKeK3vOqi
UJG3ydSx8kMcxGb9lKEhfyyhmijMyPtYR8835RWjWVItAN7sVwqV6K7s70VyWSKjnzHnZ56w+md6
45jTOPbVXXCRQq90nYzVOHz1MCjkeW/uw/Sfbj+3V4L+JSB/hXRXpnkjeYMWlNG+iw88hjUFIg8I
p1iDUFCFdycYoZvpuhvYnFNxuCWQ/3CbD0gtNHZeVtWxCRWCKm1wrVIt0CQqaoUJ7BGsqyH+DwwF
HC1ql0YAdfdYAWLYqyXwUvNTquBi3remjM9ljrZ/blj4AC9igkQoZlwgJB0bkLdJ0/pttoLhJmn8
SscFlwkVyHCFMIFESR9Nrn16rNVz09JoCZex+Zr/OTGtqwYZGAVZ61J+A+Eq8JQLbbbPMnEbuD71
oCJFem2V3HSCkSGAzreOMx0grhq8T8MIGqWRtZ0dB3x9QHv75um7EiANox7pGKSoBEkZxUGSy2Gj
SPMOAminBghoEJeQXQ6BdzUxansoxLE9Zo2gQ+on6Y+BYpdWsKdJ2/visbQNoAc5xFLaXVPv1M1C
eIuF8ZUtd8UPXDyFzmvL99+bsFhLqvWj3S4LApEyNtl70+Sml0OVleLoXD/k/hkc3XH3u/UAfyT3
N7hNpWyA14A7mksWKUAjuT42NBIL45deZTUjwD9UoYZ3XnPPzrQ4bKmCPD2yrmLaii7VhHT0Slxd
x8MOxL3y5XkaX9NnY82L3YVwfV9yBm2nlm3+BzhejG2tM9HxOu0KIPaoFdsWh+Pku6cbuuA5pYlD
vIHEmlNSBNSggetFSuAVdhyLrwPYiJ+tufRViJ2KrNrSuvUdPiH8iaayTpRkFAynVjtufTLUQVsu
2+Ledal4gyivjvzABAQUNzKd4TkL+VURclXig/LtaFtpcFZsF+tHT03LPAcRHunvVAZNJxO44P2e
Z2AOlU2sSxzNVrMP6D/vsfB0EBBsI1b15T54Y8uX1XjRtBWCY2JNfqbwHnWg7m/kZuO4R6JZHptQ
B6ucv9LUxH1qkmZWj+RwlKDScjHGveGhAJtPa/wloSZHmZzK59FAC3jL+EDkTCmz/jxicKxhPNz2
EopYwLBiaZOlNzSy8z6Sqmn7OlWb0NT+w1pU7ZYnTK/6YoOg0h2Tf0qH3wCCA6xJc5bET36VFQw4
3nH6vU4cDi6CWbd/XsNPzTD8/tBujp6d9c9sEVOz55OoMsAmFuxcsZB0up8eVt3OX/RWCKVCRVzM
HSlj5IF672BxgZhy7LNHXO4bEPO+VQFQr8FhoSfJzQaA0KiCveqjQ4m3p6cpzhLFER/ULakQuML7
WqcynMtii+8Lu5tqvZZVNTBRYPW9Ws62h04K/OLEgzqHmDLw0SsJbm4A5NHaanP6YPh4ysCT7TIo
W3RFfEQBzkI1wKRxUuCx7ApVn1nEu5vcpFfmSAMgKnja7Y9uQ/1hrnxZGMOLWBEdOvFPvUHoP/GH
fceZrTFM9KCxue3oZflj6yBkve733RRLRqcYNZdm+8tXPdN2gqn5u2A58QOrud/MCE38GnDnc/2r
e58ZnOGDY3Y7DhdadD+BUtZUnPpowsjQQR+H0w9JVJ/q/+NP0MoQCYWCft/QpuY+zmvdwgkfphmq
r+jsz4t7SLkSuaS24gBJ9zVWdfTe7QCnkJjVU1NIm5T4g2koXOCIivBgjRx3/JDwlV1ohdIkIJud
hLrjET6/mTS7gBouOI1yTk8jFJ5ggFqW4SjZaZvytl/jBiFK75h8LO6WUvfVZn3nz3848UVsBC5N
JHqzZDHrlX5Cgm+UrtFww62dPYp8JTSX4rY5OOF1qPUKis1iwngs6h7iWDABwKNpRSu/BGs0qhXM
6cPrvf91hc6rA0rq+a8/+knbCGYCfn1Xb/K/2KuZ79N4LG35+PzbIOjBjFOY1XjhzekdR5sgJA0H
/I29nKXWdij+IQa3IzIEaBu6Z4Kiteyy+gizcgRrN5iWWqo/rBgBrvs9Bzr9gm807Ct7cOMu736k
og+MsHU1lx0fzkS7vZfmTH8cNGe7gT2ua8YnV7E3DR2AfSV18IKjhenXXy+032TTk2o4+IN6hJKt
GoC2T6IsmOIJmGI97dWFzFdnb1sdY/kFrApqoSmMJ3zN40i+uM44gtJXHASPlFSFaQSpqMWhKUle
fzC0zhNSyNkuq2lWeYZ70hj/71obsr4LkyMr3K62uMDWKws9xzglxqkykgtFJLxVleOC+nJP4PiY
mMVkS0ldE9HVbLlWRDUgUKoJyY5ylcW5jHrfRZPCxAGodnw/lgXgu6nciUYpMyUJspx/TTbfonaN
Od1XDH9YuRgVlys9IV6F4NJoYZTtzoCynuYRMa/MRGYnjI9qi0ZqeARx6Y0XLNIS3yaXZ3khAMOl
2K6pFPQGeTG3DN1qDzInvE9JN4LlyXOfw4p1Ch8Wj3J4c/mX6PGWUZfXRrx35XzwrDQGZMVydyJT
tEEbL7VLJX2jnLRr5u80F+Jb4wtx1S617DC7DJDZCyft9MSkwLrpLYe4Pbd8b2s49P2q19ysMAmn
d72tZegrfz/NsC5YQM/cuON4/re9kqZ8HWH2EN8uFwVdnmHvJOC9sCdt7ZUdyPsiUK6kPtTXDc6F
ISgHf2wPgtHYeCWlND8DW7R6s404rmSCRKyT+FnZrlhJ87aIFa4kJtXjnAsK1Pybsb3hdQZcgBte
ueHXGukxoCNXKw5QKl0v7M0ROGs6t4xCDjiScYiFBSUlJBR7qlrgAUdq9ExrMhMx0/auejRiBGI1
EOM3Z9ukrzsN40pNCNRa5QkXCda9K14E9PuxJ2CsBGymBiWfkif7XxFc/xinFoQYuZanHC+VdQu5
gnozhalzChMyS6P2JkjGt3LWSs1tzelJkD5XlxB7iFfgUXmw1PmpRuaiugIZE70kZCBV4NylX255
j2kViKv2xTr9wqYNJxy6NwzM+5BKqwdbusp+fRqjsQL7+HkhustkKS5NKinOSRadXuVL9jWYKmUm
XJFwT5JeQnhZhzPZpFUwXDtYpE5Q1NYScOLlVsrEFP2URAJAD8FnW2ZSOAbLRAmWwbF37Xkj+Nrd
5GGxia8PpHEgYsvXZN8bbUrVkT7U/Koue9InHfIMc88kpde1PzIJlsZAbQrnx7M8z+IQ/LlvEVIG
nMsZ7cKF4Te59OcQr4KxkptQs5/TlalAH/fOPn1mNrDVT+aB3IuVqab/cd22+QO45S2CkrmvPher
xHnYY3/SivvUYgPmhuwGC3IpAtTi4qYxRfhdGBc1R6PKaSNOmLTcz7w6wi5z1x5CTDWmBP6XulLb
UOjKR9mkFQOtx3jR2Pd9+OqxwHUAUFUKxQQ1BphCLW51TCVcHIJ4S52Y9Cs+k5AkFyAT3Kq7VLw4
xAfUyoUoFcXRPSmhGgWPseJq8HBoeY17F7vnpMlJBV3nDXDjdIAtQvUIKbjf11ATjNZFWg+OLpCH
4IYZzSS6lwR1LM1XXQosGYevsU6p5X5XLgp0LbvYmWPdD23GwD+AEiDNjp3AYZyA3tC5Y//Fi+KH
3K0BtA+Tpie7CeDSUdU48PJvP59gcsjdrgRQn512vSRSlcgSD+E9HUCNEJdSKU8uu/oUdEtLwmTg
ccBOfPnXHQHG2vpEI6jpjcyX1I7kGalo5tPtMMOaYUrwEu4HIC/wqmaqvvSAZ2vR6MO61lEEe1AC
7SydJk/fIefThynRNti2F6I+Xf6dYFj6yuGHVVO+rnfBK5dxNQzYl34YZnOec4rLZng7qOR6nvlF
CC5pl5J4xBOKXw0sIRxtE8IlCLSxOoNPxOh2pR9Ov3/ZGYFBby+b+Xf/iFElRL+8O8dL9pHd38fW
FHte9o+YFWSzdIO2xf812y5F7ee3688RmjYvbze4rXrxRYpwi0KnRwlpYVgOVWvyS2OALqZdkx7f
Iq+DKN73Uz5+tuvt5NOx0KS/Qy4/FQeT8gxz7SfsiY21wYXCN2wLh3/Ox0ybpf+oSdGGYh2tsEAp
C85PPpYDMsr+Z18X90jr+Q20Glmcpo6ECb/BCSR247mxDUVVZTeziLw5ec6z/SmqY8+dGuoe7hOA
YT93XEA51RMkyn/JOWBnLJ6RBUzz9j6lp5JMC68JjRWsdQzscaBnCs2GfjWXOIvWn1pKokbN798m
nx9/5QEmcNPQI7CtFb9i4VKM1gXlrvUk7oTjzDhX0XbjXRZj/3pIGkmKe8MSNVkRBdjNlkmC3O6f
WwLFT7LTOyySVUPSyoi7p12qHf9ZLEK0qeVBlJqEqiIsFPgm0+czScZycKPxYLQpjhURYgkiGEz+
DG76e97fqjMWp7gS93XOYao5ae3qyhlamgMUquG4JsUTF6V8W1oFh3mPT9r8u80qj1HfzjyOrEn7
N731m9enUw8xs2HKel1tNC3EDliW7CCwmRgGlyS5y9n8Fe6S30g/ietWMF+LmJAhAo6j79Qos/sc
Hh4Dd3UsfeNXzgAJmukUxFLA8HsXbc0mWwcUJWWE0wSRW+gf8YPQa+y1Nh2Od4hFtGAmsG6IRuQF
1rzPsp42k++sTZVLZDddXDWR0lokaxOW6oUmHmbfRpsi5YK56NoDT/E+guwmjd9TTz1/8UdUGT/N
UkfJNk1EtLdOVMWNCx2HLC8NbpB8APBb0pKtaT2f3DJibyL6am55URRhSxFAbLa3xVA19LuYhZ8R
caRSa1I/bGZjHytgimyEUkCu+KmFiynKlT7Z8hubcnWLEqoUPohIiRci6Z+2uqzs7edx3jEaZyMt
HFNpddWTy4Ix1EisImibZEua+3SXFivlbBus26Wdk2m5QNEN3QNVCBGT4eT4aw2EXVuEb2TA8kDA
LBB0M2mvmzGAfezs0ISDy+lAff8e7YmDKJge3JsxQ5n/TjNfWN0w2JSOZZhMeZdnkCeiJY29i8gs
nuTMWPvAyXx78V3GV+iLdNRs8o0UM93iTBvs8SYLBX96MYFqxuZqMApWlpJ1sFNeY0djciTW7Tbx
mENgdsP4NvKKD8X12ghU1Y0gs7AxmoroXe6gYox0SiiOeuBgjpH/SvqUXOgCSeND9oJkMCYJw83l
R/ScgsDmSgkbYWwTwaP1+HWrkGCj3PI+0ebx4saMGtIuKTsR3BtsXamMoTIaP50jXqtMQIyk2FlJ
YLefYf9XK1ARw1bKdbpgoF+yKEmrxX6WAcL9CLu6njwBP3CQzbdB9xzSVsh2VmT4s2rcHp9G0XiG
8PesBmhTwwPmAH3GFga4Hguypwq1sc+tdjKdlYP4ZpBa9XABfkMiWbdqNFZjSJswk4AqxECgMDHu
UXqGzHqYdtXTfH75XzayB201O91VcJYYBwpHVTF+K3N63ZYInuH9RBDnCRqlN0kVmIgwGDnbt5RS
LwbHPhO4+lGMKAfMM8qJCo96ni2lu1ERgKVkVP0PkySC9d2ttj/pmJj45pZyrys2Cp6NZapGdq+i
ec+xLV0Z+Hq6Y7nhWzs2HsuOBsI1lryD2mfHCt7OuR/RusjPMqHeV9KEYlo4XClHoBpBd4O+Wa8W
iBeUNhzqJ/ZS5OQUQaV5u/mruTf7F94nGCwFdxYSzruAoc95OTRaIRm1Ze/KEaPG0YrJ7GdR06IY
N2bi8m+cSvst/CWk6PNlvwwQ93rSgCUXsrzW8aKnZF9dBhdO39fCpguH1IUcTg5wjhNTVFKBTh4c
mOvvt7HdWU/JbtyJd8Lba0/XE6XnkdFj2t662EVVtPzIM1wCJZY7FEQmxcc/WZjVz6qPFKe6Euhm
Sje+/GnJPBOowqO5QwN3cr9WmxCy1uUJY7c9qALFmxlnU21JQXfNhxacAJEjZ9VKnpfkps0Nen6T
WjXOD371yQxpSEb/u5t9pPRtryCrCtsn7HHSwpZzK1kFdwagEjy36wOSDx17gy3satWn5haKSUNk
gooK+N+n5dvEUOkcj+RTCP4EHV2fV+1dOWPbKKVPTCE27OVtHYI34yHJwobxCNA7bo/M06/kjpg7
+zuRMfvt2Zxbh5L/btC3D2jtKJcnFE/tK7/+e+b5xdmyb4nzzzPrGfpow0OS8P3RBGlW/GPA/KdO
OGJogYy0dPCJ/mWsRWpdjbCmvwdghScScENI89TaMoYjo0FHSr+Ap+8+OEXmQJBjWvAs1rUBCbD4
C4lB5NORqWL/tGCVQl7SO7iV2VsIjDuGuRSF2WJJkrcecFZJ2RDQCuCqS1u3iNs8SJq5hd0CzKDp
dZ8BvZe8e7YZ9W0/itTnkpU6QbvubSuSuJB5FC5KBCrwosjpO4JqVkjaGn3J8Te5AJvHaUadfMyR
I/X0a03x/dBG6Ak0FWumhVD/hSOrD0SZtfWpGK3sJB55AdGeOQ6eOYvsG2XDey5b0vO2xnzVc1iO
HO+XRnrZFbhhInRZYqMe7pldQ5va6wzergf0SMkEOPS/wX48kXrsi34I/xBtIXKo0dBQniNeadTb
lpjNIB0DAhRh0zM/UiKsYDitCBKF07WJfSz+TmcXTqo7wF4lr/fjQjxjC/mtcOXHstx5ELDG6F7O
ghd5h+xIs3EXc+xYupbZlLJk1PIR7+EmsYmQexDecoOaRJaNPTcmCDx2sgibsUGB7uxMuBEu3TM4
HbMPh3JbY/suvVNILmYx2GNk8vZdof1WhWZucKnP3G82F72gb23unKmhT8TlwpgkDrszh0djkJP2
MdEryytUAksFae4oj4lwqd9Hh+sWBxMITjaywj1maaAgmhYftWYwqlh8CvdvLZnEPZABy5llcGnQ
wij8/sYh/IGyNA+FETYxVdh4pevG6x5CTtQAfjy61z5BX9ca7LqUNSo9TFEsZNNJjRl3h/TlQnU3
WPD//c1SWDmtqW96ys8C6tHUBrCOdyjTVkwk/reWerm5ZNN+KGSX7ppzI9Vkxo8Q3EmgNVSqWbFg
aePOoaA4YB979SdkBcXDUFyP9OgoDCOzd+ZSMbYAQ0S9eJkMDFZmstODWDQItF0KNYduogfPB4yg
mETMPiSc+qZ2pltGhFEOjCb4RhahZzeMVU6W+jb9NT1iIc2NjC5zmi2Sqn9EUwQSNR/E18l/2ntJ
B1ZM2YMhns8H+NilU+EI9LWjhgHDptScCnwe/kiH2WFfMrBTcLl+sNXQCT/0gjJGWZFRiLuiFzle
qYrDJ5NG5sA+qKYDHY3+TGh0SlbduCr9yx158nJNccQS31WmsPuIr6KzGnHZDj6YU1GGaCU6oAWF
se07tD897Gwi/S+ehrLADre8z5Y3RlXxaBvK1QN1Oen8N4frJX4bnYIZI6nmytyZu6UlSkk+HHF2
TF0148wGH0MpLzXcyDGfJsSle+i7tUzKgGs2sY5CAckJ4zkbPVcVn3d0tn8Lr5rO+LIUYXEM/kL/
e3V8OQ38IYXv3b7/P2kT3C9mYlcKBwYcjQFDHCcaCnQ5HvCzC8K7WgvEq3Xba6L5wcVO+ZQ/sRqh
xJ3zGz4w/83H96ssVGoW5U1AwyliEACzXB5DxGU4XuUWgqLw/yEF/hMUvlm9svUNuZBLaws33435
eIlNiLnS7YV9V2KA0mJqzcSWI7C7A3z93TE9yqLQvnDpLqsDilvdtFWWpr+LTnaFVY3GaqJDPrzE
bCxneibiPM4XetduL4QBwnAN/C3tBJrt/nsvILhBoNVMOYoucR9WIv2uSQsb+umYSpuNc5BMrz3T
HO0GWLqtBpb+uP5Dhlc2lozXzHfpIC5sA812AbUPQcwZmVMC3bPUumNPz86s2s/Fi+7gg3jn9g/Z
WtigRQN69ybMijHLKjRlrvzdvdljFFz9mrnR8mfQD9XPddGth1bHpHzEdAZMsNJwbKJ5OvFHpTDA
Wnfk43IWsyI9AerAF2mdmxDckS80HHqTvhvcGsQldxMaE7F2aOtwjj9ix9yNnVza9LUUb8LoXTVK
k8Iyam2EBYtodgxiNl6qkGfziiU0lqvNf2J8S4ZKF4K1INwS/2tXa2mCmIzWFxIkolhydm3eL7f3
9I5PKuvxKDLwU+mFsUBy6q6Crn4X/heoxbd+/UDeEROEPHHsrIlML6fDdvCHQPYqoA0lAC66EZ69
vvOv5X+Anyv96k/6Ewu9AhwdPxdJlPaw23D0Z7xDe4hWMKz/An5XhBdy/WnBCdkzUnONT/M8d5jc
V8QzodciBq6E31kUGizgRUtp4QBKj5r3zdmz7Pod7/ALHgD1YFYlWJrJG6x0KRMxUJZqrvTmR6VM
l2Td7JnKzdEfiHxN8DduxVVFz7geUND3bmTOhVt8o+F1Ek45E51riLqrWHTHohDEeG4b3sfl02Cn
x0vBKB+OABEHNb2zl+XxnVDgqGK635LNtmn23asR/BIplNjZCNcR4X1fuhJWPoTNWSw0L96OE/uh
YumPhOiISsqWgcipp2OqFaGGDPOjnRtEybvdHjkxwbw+elSI+/lWU7jNPtmZP1sUwDOj5pOEELQG
qHTGoE1bohrczcgesoJVoOm1I3iyYly1W+x7DUrwVgOKRaBru5H+a7nQ4xRAmt/gMUX5r6LE1I8M
5hy4mY0onikx0OVc2Qja+icnMuLc3oTO1cU/PDsGGNPjXnS1kqP3sghrEHDn99XxnjFsL64GXn7d
O+Mp25hd247LV1XdzkQk36QIda4ePvS3UcIdsqMxNILyiGKBjAeDHlzQlbdrlQUzfQl2xcZnfmBD
+AEVhlm2ezYjAsyxlTJLUS7rCx0iSYBlJN2fGc6lgvdvQ7fD8qlo0sQfM7Hkh0mwY/I9Ed6q12n7
ql8Q+HAFXxPzO835ORjywBfdLsIwFC9DasvzYn6fHpayRm/CZJHPLG3g+V5SMVewfrFag1p6cfrZ
BY4W5l9XgNVIZ4fwiHhK1FWbykVN7RgGSyd4jvs0D8pV+8d853l2RMnA8oG8obqOCJplEkeMZkKV
lufqDI/CezuESeNfSEk6BoTRw+g+faF7TGs93vialb1Lf7M36bG+XRPSKiiaXgIuAJ8T6mgmXeOQ
UnU+SdXg3KfywHBnMhdfc5wFR8E4vtpFx1LQ78QoNUsRfwXITAvrc1H67e6ScoRJnOM1ks2FhcQf
iS+THT3zDVBgeBOvqtzeUTt+9wCxg51qQGNcX5YDj1aFUyUM8B9qdW8+B5dXnE70ARmKFbTyRcAc
fYurHmKuNNzo78g1AJfAORnKUz5V54F8Tvpuh+NT2Fo/b2fHrjyodCCO00NpYuwqi1z+nLHx7ScK
ixlO6yQzHBZbJC+FszpjKq75t7EOteIRtL/G0Siua3WF8ZKwSY4Gd4PTozfKvg+n9ZILIVjgDY09
Azf1Be0I0vzwKJC9oMYvV6BqIhASgWsT04hgnTSnNo8yCRcmR5G4xYKg2ecWz0uZ95R97J84bVFQ
w15mDz7Ii7AbZqVjD701DgnHe68fbRRlkRb8QhNtSh7uS8Lku/KYfw4ms4P2EYcBtEY4hhFSI+wR
9OaLKdrB4Rovd5lkDM3TOUV6K8sobvAI8aRHU+Nf+4a1QjkZCT2ARvquzm9RSTmeMnRrtsSsBjRg
H/covKREVHf7WN3FDvfzeuq7bi7mX+ByzuTTYqTJxrwcxV6wDx9H5k4mAheAdzeC6OkhvMD8zeQ4
7OizvggMBvn3hIAi1YZOxu122dkDtGq7VcU1V8T4d2htGQWHivK4FDYGNCO7sFcu8GeuaMIVtYbR
ajLK4GzUkONZPuCrmcS/zt/AyFt7LhJe0BYvNqSIo+3nq1BHNHIUNr6vpxGvLN7y9V9wFUUey1B8
n+JvlJA5i9/dBk30RIt01nq0fkglsJj4O2oPWRPHojVWPL4PiULhqpaKoJJLK5Bvvvx8PdUhAlWb
A1lxFlDEhoujjWOTQFdewVUx1HfECsCoIGBMpnxcXv0nNa1mUxKOig6Ug1Lpg34nNtCMPgzeI4O8
r6OkW90Jr4JqN/iXuKY4UTTmLpBLZpJsGiLOU1NOr3dKxHF1qWo0RaWhx8hQRs9U0I+GgjKwjfrr
jGJ3U0iQ+waulIAm2sGPbbId4e8VETjBIiaC5DBwizndi0ZFCTjTPdMGMCFTUhgCQjMY6DGE+2Py
KJbbbSV6HgfviCO7TrcSawKiMgYWdSNfKVnpmn1jlqlh+PdSQaQIBRO173Lu7ER+ORhfTTinEesx
0sI6HnNg9Gs1MNtKhdhLtYdx6bIEPMs1cGWyogho06cD/RF6hpCi9MHzIBdPxE9z0SapUF/9tS7a
aj+tjz/0UK6dwuRddR5FxR6YVybHVuzXtC26tGkafWT6WeVHhl6HTiRBQj6DoSj5vwQRWP/tqPh3
Sw2OtEKfQrypvHtEn9CDe4Ocz+fJ8hNsbuVDUCXEVkCwaf5R9ESCR7Yu3NwqY2xE+Aby7dmTffvv
aK7khon9STBqbFTt0vGya6vj5+/ssWhvLKZ1t7quz9stDmeRoK9XMJzntfoRt0PxStND74pmX+f2
Vpmq3XAabbLIpSZ+EaQPHnOwlaWEeh69FtSKSG7/u7MZVzezirHIgnsf0Sfo8Or6dOy8CdRaeE+S
0NGPRW8y93IqrWGi4IjcvPqTCt4W+lXbByqTWqxMj+3vle4Tpk5b8t24GD1KbUepI9XxrP8Q48e8
P06D/t879+DQtmEM40Vj2xaO9coWiwMH+drammd8MfyexwX57fiMqq7lSMo/XA0ZatAZ2W/CPVek
VNAAqM1Xfff9dgvwCoRTdhAl554ulIe+gL3mWAfE42hWrGwk9SsI1eQQaT1ZtKEvsyrqjKgvUj0C
wcWzvoPSaHwkhZ4XZla4VnOsAFegPfoavs13m7qREZHPvwXjhgOIMf3Q39IUqkBBWPbP3X9spmb4
qMnbTMC3KL4y+2FERct9OPsoBc955wZrUl1uJipGj9LgKh3L/LYHpo42GY2w+1HjSi76jswH/CMA
jJHm3y41KIFrY4u9IO92pUAThp8QPXYqRPBDAvfyeHi1S0Cv8eJxgw/qBLNAJrwU7wdxz23uFT2j
D6y8R6f2k0zxKVt3o05DP2eEo9ptA0s2tYCzkDIYxqG+rJeDtJgUWIB8RxaTngPLPNlpAdR7SvZs
z/MX0nvsCMM0PuZI88pAZx44+bpAKk7dUI7MjR0xr3CeO6VWqyNmkl9hgd5TRlWh+GNaxsQTsbJg
Fa9/C+OuvivFa3YRQwAwDzdhKXRVsSUfoukNA8i9rGwV58Q8PFeGcVUA4kyUrT0NCeUsIYLOZi0T
K3+qPQDhjqOYnIGBXS2CD3wzTAY0YVtNdPubj60yUMbUtfA5dB9szEZWL/L4JT6U+K8XXRe2Ip2G
zMdDRwm7XHTJdaHyI0b/thgzdDGDAUVqZqdXfahc+Wfb6OG+HmZF0gxSFdkApz6zuT/xL9XsO7Hx
3ipFQSDs+ucz9qyrs177ye7h5AGAe9A8ch1UsidDnlAvG9AMmL7ZVqPPVgAGId1xQaLEknQ3+dxC
WEOUsyXkSeHeDH2H+A171EBqSbFzLBNjWsDPF8bHg+8UuKrC1Ag+lInA1lQG5+RHt4NPabHSW0DP
VrPiffMO5jQ/ecv0rx2xTgl6LhQ9zydZ8xeQt3MdEcoe9BtPvWmdbAVGeVRq+Ar26exLuaOpB7HD
3bQXgRmvK9V0luLr3x5rRaK7GT6pLznQEYH9sCrlRnM7hRgr3+qenoF76fuKVgM+ckE1yFuRCSSN
k9XzjtqLlIbGQouQXD3Gi6LYmdcZIOvh2r5/bL4/BgHAC9nSaX8cwrRYIHVqetUnHqWyOHI88Ls8
+UzttqKtRoK/K/U8A/0eBr1kbf4Wd/GxRPDO4nDVT3GpoVmf/H/iQjy9qr3NnogZG7zfig69igeT
clfI6WG/2glf428iRAgW9j6r+nzr8y/ZqXZNAKAMVuNDKCviidPuVtdvTxUt+R3xk9+9yILYXT/G
Ktto/563WMM5NHS3vC9m4w8hUxkjHJC3FWWUsBCXnh2PTKdanOusYqBmMqrZbr9YMqJ0REIFpv2N
ghOLgrLN9mx/oJSF9LXQL9YgpRj9JEXsBNzDJtlRUiWwGowWmuBv0NW14XniQ+93BuWI9hfzTDan
GpYX8V4yhrcZQaGgL2TK5ynF1AFskbmexsyvZbpPqIEcbJe56iaT76i7rU7X9cMo+ALYGOA0jpUs
bPk96xM+odfueYgnsOCHOfBP3q1ooSJ7HHb2BXMv6uK/cdLS9WeyV1BGx9yJs6FEFF7B6+1COrnq
cBYeFfIGQQJem6hY6jhxJVsM5eZnDYyxF8cgFt305Gu2Uv9Pj2u3KqTtG/V4oIf9CwqWDNh+GGIE
yFfeAuQVNkP/cZW9lAAilx+tHhfDfJQhlkoWkiuMYDKRPEOavUe0CCWu+GjR7LA0pBVsSWlu2qYa
xlepNeV7nqpojexLAGirZ+E2QMRWt1oKB82R5OSOc5MQbLlCHh/7DqcYtsk17SSZcaFVHWUTjcfv
WyoJuaUHHztbWAcnZ5j5SMdBnkLJSuBl5BGneEVf2yOMi82Qf8U4hs4vaUNHJWY8aArXCNWOFj0v
U7+9eACIEH4NJ71Lc1a4A+8ixvanSnBR6dr0OmUA58jM6vN3Lew7lOrIUGVXAM/2+/FVlXYZOfHR
2eXJqizohx6cg3lSQLcNvftYTSZS92Jlq8xYylbbgYRfFFZAVG09ikZ7qNjKVIjEtrhdsVAEwlQk
1HbF5yCzQgYmjsgi15/a41419UpAZcpullsL8dnNn4mfBVY0fWv3tivOMDgMaSA22uTJtKkFvtLu
NMS4cEMA4hn4DQbxvKx3FUyqJt8nSHHRQmGoR4dYVFG8Cdrlu73dKeCIvZwd73I9CaQAOAStDLwt
ViAWjEQfeDpJKSKqsCGQxJuMpPR6mV2a+sIXaIPNaF/7J7F4LbtLyCiX37syAODiIdfc0G7t66Po
voMM1/V5zv+MTXHeuXari5rj+dVyd1AKFH6hZrmYC7lIlZmStOccKw/zmqdnr6Bg1QSrz3V4oKFX
bHW+AGFQLfyoSGgMLHUU56E09l7ocL/oD5fR+TetSE9XjqvobPVc5OTDpDh4mG4yMwZANxSPwSMH
1vfyLoiHyverQ/wLFvplnydX7Pxb+1HcxHfKuO5EcxXGqm0p5dO+m6mZkzOgW+zCcuigIrF6HH00
H/0mYOv7t8ksbZ6h3mtBeqgrI/iobE0ww0BkXT+pXC37b8V11oqeWCrxEykxuxls3GOaiTP7ltjZ
O7DPL7c8RwZ0bsUn/mxhoINOr31q+Ajr/kPRsX5rSerZvKrE2XRS7KtatCvi6dBBVAN/w8fqcTHc
UJxyNVcAYdFY/2HSDlbGVyi4MqTkRwIXylKBJlQZTcg/HvGBmUjG7VVlf4F3cjJly+Edsvx6sjST
knM0i81hhDeP9T91hcg0bwsyD3lbFTFn03Zkx6ZWU2y9UtSmDAWfNo7MIKRdN5KQ4uoGq4mprCrN
zJOQdWAG1JHdbdt5JfFrYAmlS9isOMYnStdK6ELsbW9CJnV6rGDW8g1lLFYGp35gAOUxl58/PI+v
zYXzwx7bUC9NWQFrTGYfWIvBeQ8RTNLA0Pi4iIIBzanjGzss60TdA+Fnd8D20T2zuxs3qSk+1cW7
Rd6UyUNiJrGVMx2wrqZoObHFuPr0DgntjWdWlkydYkmrv7ACLwKVL6ok4PhB7cZvvpdAB3jC9/c/
Y5DafWZYtcU2hGd+eXS2MqH9a6AWX472xTt69U6K+TUjiFYcDviVw2g9O8AX89+vGKd+/UlkBmIr
eGX2vx57QeJEHP2ofjL1GriDjLth4//RufYZdJ0Opet2g6+T0r2yrW8BWPxSFst4JsL05bRkT3SA
1VcqrTh98PYPfsZr14MA61zXDbvezIaqjotsaFCxT50N96DIu3uLuhKlvTrQWGisGNFmYcPO/pFN
VHJkVIAeFHTP5GLlzkPLJbOdzhMPUzLJ8rpH4AG9/0+t0kfasJbwlY3I66+puRknnbD2ENs1xLl/
BNXvM+Dwu18S4hP9BPbzK9O4gmoXVkQmia0cALJICQmLl7j5DBVXcXmpRFz/GgvpL+dj3aX3241r
pIyv8JOppFXE/OmrHyqA/nvE+XyaBrWxcBCjLXF5fSn1UzS2Ke/2y8oCO23pWH3j3bI2+/GSq+DW
taGgj93QXr52IOg4NWdlIIWbkMUB7wQsTpb1XQv0AN8yhFt9k5H/4hZd0jWuJ3P1JS4SLUYH6Zt0
WewlsPg1UtzRmWsrgIUBMjLwDtVrzsM5zbZg/ZtIbRwhyDhG5EI4wsTOTXgWZfY1JRDk8Il+Q6d+
udCfY8+cO3naYhFBGXbqRzNWjhBSTSRKy9ffX2/5IQQqLzAo8m06y+tWaXqxjoPRyUfyAHLSuH5y
HxGs1pkcPFXUWxkRiQA6eA123d67sUWVLqGF233XgSzyBmoPzvNkqSKZacbdXt9YW4MmDeaK1yFf
o8mm/HUtf+VOEH3s1yN4a9nDnEicju0mnfIdKsIXAL1NME0eHorUFdLAefqER87SDuGEV7GrNw5a
4mj4ZQ6kUE/sIqgZBpSVCKZOE2Pe8/hT28zNJ26EANMrOiQVYohE8sordM+Zl/kIJjdb992IgVys
gaGNa3Kzt+kaXpLBN37pZa4jWrzu9akvKS/dqz5BOUH2gYWTDSwT4qo+qoZVdIJ4RyCvIRrNUVNO
4hfZ1WQPa+7GCoKR5/6Tmtapx3DEYK6OqXNaBzVwv8RzDWiHiibW2I9IwHjTSV+EqdNiX6uq7r28
sNe0e5hm5mvLoHIVju4AYcwnNSCrT0fBOJEnKhXYwgMR+vx7DcPbCBKlkgTyvO1YKjc1G5+hqUMK
sXgMbNaGKh3mK0jAcO+HQevZ2jFa8KrPckHhhmnz2+bc0TEwmeVFZcw+tY/BvCU5LnZo7/2L7W9S
h6T5ZmPPFSGM2PyiaprIhIxdI3agb4w16vXrhOEuM2XdszfBS5Sm18awFJJt0c20pC+1q2sP75rt
fjCxtFv/AAVkPgjnlOYDXXJzLRW5xROzkp7yyZpOLFaGRttq11sEmqp54xLO+sm9+3zGy1rurRzA
O9XgjUjKi8Qem/lUhWbiPNqX05oQWvvFDaZOA1OQYJYXbIhSc0Lsvfokt9pfO6NRH/aEJxlFM+Ec
O2Iyvax7/EQR3TT0ZTiWVDzoPRMhccB+30O44c8/oPTHNvtvDFKlpSoeI+F8UqghiwPla7EI9ZwT
QJsWtUQE7OZomzkygb7CvwKvgUECruBPayEoXYQA6voCk253cTXVx54nzs4T+ZhsO7lDMpoQw0UQ
q/Velujv0zU+5ZYMAgczv8TD+jqLGAlnAyF80hWtjlTgoTKZtklLFhPxltoFtOw0sS+DMv6xWpNm
nMg8Nk92zucmv39PJCP97nxXlBZmEZvS90nQAbcM2KXw03N74xA07CVlkYIwNDzXEHCvLb0efgOy
wHxFoEJYYAuc8Wv2mtDzlIuY3H/kJqhEeUcCdGO3DzLN9pIuoT5JegpLrUs4vWUFSsDQdp56e5L7
OkzJO6XqDF7IsXOeSlEfeXAPruOgWDxOZsKcmQXhXmA/UtSkJuXyNcIe/fwLtU45G0zbEKXs8qVZ
H3qRkAaG/yl6EUQAXtQMPXLBS7W7fjh4Jr3te3zAc9nUTKCNzolJgvOys5x7g9bIFIJvkxl6m9Sb
sLnMantNGQtWtlPWeh+MqZAFGo83d8jY/GJVZ1FMoYokroG4Yx8oWYeEsSavVGkFsQTZ7566Q3q1
to4ZQKRVfl7ug0tXzf8VqfJ8eXfJS0WcZfLf2SQ67cVX/IB58Z51NV3T+JmmgTBYresdCrbrKr+R
Tg3YDWMzybKqPPea+jnShcD1aVmPbh+Fzy6z2qx7fKqJiwM/ReHm89J3BfVoVup886AdVHKlP+la
gRylt/8ze7K9aWMK/qJup5SeMsoshUD83Y6qw0xxUkI7EnZXA8ZF2Ys77Od+NMpxuhTJevww5KEH
ZHlLUHXLezU5DfC+4F6w8h2y89cxipABBqzmSCXhUSVBZLeXPX7KkitUcvN6ubv5gN9vrjqkcAiF
neeS/J4dWBk0DTyLEjgKWdwGgPVN+BCq1DpbDonyN+0MmzXKxQzlFfOkrIqha2n88WNeMZWfWhUT
tnoJLN9zti4AjAWf2HmDudTFpNDs8qI/I4FBb4tRkFecaJXBrSK+liy6e/xVOKq0RQLzskIJjadq
qdyE8zTU8OIK1ye+ueoEbYC8o2texos+ja1rNCILSjYeoNPZeCrZlgV2SfWz1/z2qcTGwBfwYoVe
+K70mkC+VXRanDgV7WHLP+O63FPnINhBZqkdN74ojvGiI9OD96CdqlTx4SwpyUhxh90iPEHW20nL
AcEumudINUfCWoFdpAoHSDjwFUTvJ0AQRPFoSZXf+uvYihFZuvmGysfMUTryaRMo7mlR/7S9xzKk
uwkXnEISHPHkf1cLwDc68h2IpakbVa+SmIFEwQb6J6LFScAPoHTFuNgd0ooBSIckAUO48kiYhasE
xi8/rS2SOiozYrP8XWbhE+SHM7ADyjYJnoA333W0IkclnQK3P7MpzYSNJHa7Zv0v051I06/U4Ds5
f003yUI4cDDjScPieptkynX/lTXpBYmOAML3102VEwyglSX3zdeb6RVRbUzonBmMh0Wk2I99SK4e
rdf7bd+KoAtBrURhXdDLQOL7ors4rfTG+2QlP8PC1Sc1+rkD6q0c6sL9pHaT1Zc+ns3HNZBvI528
43WKU8eAeDvuVpZqoD6ArdOUwmYRBDE6xX/uxgllBO102305kRsNZnU1kCtBRi9cTNT801h+Uf2e
0MJoqaSpT3TqpzzRsqwQ7OtAn7lAxTuXCuBws1t2kJn80ba35GkOo9P7oKJg51Dc60JSfatn0izy
RQAyusOn59T6xDWAlwvn6SN+JNmB1DrscY6whSuTNfbiNpLj/my1ee2ixzo0m34jKzt1uMBpTpft
FIQUcBKn782QIiWMsURgukaWYIYXhrpjhpehKXhitZmD3LX4fUKfFJ6ZqEtpuARBx4rzvRMBDkAH
Yd41uQRr0qyCQoLOMjrSKxA0cfyLJpp7pDUU4OXyVknWZXEPBdB5o9Q3LBb2Q7ybXpH0fOx2l79X
mtb00n5oSYUg30INiWQQpNIlhr3qQvIy2AeDLm2kS/vc9Hd9RXulw12NVnjmJnHaaRvWNMRf35XX
HSCX1uaw7cKt04GLuyyGPCvZTeg7h0dlWhQj5bfgMqSOCU/dRfyvlNsQ/P7r/MApRBNANVVG4mr1
7g/+ZPbhygQ2OSq8aMjYYswkY9gEZ3SAhNfO2hXBb1rMf1deVCYE80TTMM26Evi1Kqwu75kaUpa9
aNCD8UtsNFyhy6g+e93KHiz89M3Lp3yZRG/yLu9mip+BszYb1UZo7OSqiy09jSKWrU83KTj5AkbL
vHJs8WPlTAAsFE96Z0KSoCmvjw/FdY2DC/zR8aCmqjK+Sjs9eaaJ26WmfRxT/s+Wf91TWwqrXGLH
Ewv/PJnFPYPqfJjQgOwr79DgnbAqsrqMnh0sCBmWo83IJGxXGIZgdF4Nc5Gw6mgDBOX0ixQPirrX
ugwWZ0H2U2J0bT+Uot/kpgas/azGW4ml3Z/UBps83qoqo41AOnCdv071K+0YyRV6Xo+HqxA7eMn3
voFemzHBy/7nDz4P8dy59heuW0DczJwV4oeHHaOGt9FN4r2p+Z8W/g3diNyrXR7lfCwAlJz+mEXw
2Tc+mQPosdJqiuVfshowNxIPGtPp5fXt9d++9JCPz864YqChrBAjzPBZD2L4Kl1dha/opmIBd4Jh
nLcu+f0xYRCZ8SqX57+FXMEXuX5mr9bblp02s9NGtiAOXKbagPWdCceEFgKrsUYIF/8mPz1jOpua
1qWqkbsDZ3Vtle94NaTsw2FdrMkb4BM3vcy3D1a0eq3xLt8dEVDsdxRrom54CBGlfBRhoMLa4gD6
XJ1XvAKllbQG+l4Au7SU0oOOgMFbp6WOpXI4QV/LYEN4Jtczv9oAXF/YSU7v97hFAHggHsHJoCrm
shh4w9JuF6mWlyV9bRmhjsWAb7WCS8bUONl/xR4h4v25ZRULzY4wV5klwA5CO5TwqPXyXL57oAo6
LKV2Uz0wTBPb3q8iR+L60rdNNAXQGnFNNfCNZvYLemrud+V2q3L92Z6yOEEYwRsCWLxaYF5uOlaD
exvzziVHs3zsHXQqJp/HKR5wbYeIk3EGAy2/Fk44+cSuVVpEYaZFOLVLHcDztgYg+pn99TIHaquf
etYdP1is5TiiWRTesYJEHZ7Fpdja1xibTaUic+ZCNVzjW3obur5tElfwHHwDLmxZ8KPZ+iAb6Pa4
9HTDxs2vOwR79XQUvnX5UP8oV9X6p8WNYGuEDGErnHUt5ttwx48DZWS/EMGyuKMNKqjI2oYiK1TL
geo76Z0k7znPKAFaDBohjFTlsK6FnHkBAiTfKh8WuHJE/MNY75LcvmqySsnrMnyeCzixNXdk2IUw
re2pdR7qGMnaiDz4uwmCvT/RR6hCMg5lUMRPPYvG9tErNN/I0m+bZNpRoqopAfQAMYJ4Rzo/IOjU
mru09aIyt4kNLn7JEWpvHZOvzO56ktFpmH8GTepKByLaFutLMEX6rb5bSzrrasYsruvcR47gPvTG
d1SnQ8yGZvwEsrZ21bMXvd5F7dVENNyzb8kPG6zPKy+psrlbIOdcBgcIZyZW4lahXbcfzUvw2hDQ
cNwUtiIp03XdzARh9ZRpeXxdVMsfr682T0kYyy+/XBP4KLJ5kLuQjUiQB0AKYVAXdbLwcArnePnT
GkLORuf8jJceG3PSft2MMLcpTdOz9JGOe1L3xwZChrQg4I9aAM1MxIbBgOWn8hHktdnpPtOqPFEQ
L7nOArVe3xNItIDRqNmMXt18DW6dhjI3qPe0opXjbIkYwPvsbNgYmSl5++EGuLXaBxK92rMXQTg3
cVlQHWNrx8T5llszI48ZvhwEnamfN4fTPUI7f2Y+xhqdXWWfxIZW4ki/MCcsA083zgQf5JmmcSoB
BatuCAwOCeuqJPLcLmaPwWiuJeDQ8nW3D2LmXwoD4KKiV9Ou0uDEN9ljstXb/V0kEdhNwhF4EO30
JkrBqtxUfvsHkiava07CRxIpxXJYWLdeWTLjiE4Z0VURNMj3QT+Hn8vJ5D07td7Qq/x03ETMOWn/
cGoPADFrBtVoa6PX8ffL2DurSgnQSkgqcRSAEowa8NsQg9JubcerHqEn9zJYSvmXBP604jNC/hOH
JXUK39o09twtqM27sAudHP7tPo5OZ8Pf5f5UH2g+NjsiZLjq1I+QB279If5eeAn1wj/c6IpC0xaw
vyRnBoldhfzHhgDwd/86+vnZ8IsFRIfb5TYVQP3Ol0lA3Pix8iY6QsAjqF1UzW7JOglj6IZxXiKE
+3PneoqsFaV75xKa6j6pZ9M8Av76FsRa8mSJOME2e9WeCO+5ERKSeG6zrRvfc9wMVeOk2CgUmsvL
ZJV9QQNDsBwLmeppTS8pdVAYuzzFzxMzH4J6iKdVfKKZARaojhEgmVbvAuci9IXabcenglpC5xv8
6zgp50wnRADJyuaQm7hO7QFfr/hiVrvG3+pfurSurTMZ6MtRVWTjt6C/y/3rWN7zEbT3DdL71m3y
OQkKGjEST31M/ZzbBvChN3q8UiVOJQIG4qngbSw53F0BXL79XAk2DuRbXjX+W4XHgOiwtA1hWFRM
ROM4jHzfY+f0yxw6eDTpsg8xXwQ4/en2C7EsoAHgmggjL7U/S8ebh0oR9U6iZcgpr2O44HpP3Egl
tQPtoHr8QB6h2xfyUl7w591FOffgQNLHV87thbd+RKdG1l8rnxkVBnmwNhvUH7ab5R+htj5ME//2
wdwE92Q4/OUDHNRQV3K0aZbTbjIcqzA4MlV4m3lvvZymT8ISNQiej92co7fq3WI7AwjKZnY9vKgF
h/got6IQoNn6+5B0p0u5ZwI87VNnBRANLtmKs49boHoIYgFBfHHephHtQPm4xL/IjVSUdZk8v8Ln
t8DPhRFuw2a6gJ8+akwcREbB5kZzX+5otB7D+Knxtdy8nIof7PKDD0TlwizbI0NAfyKORCx0mrpo
BT8z/Y0frcxh+FjavjnK10h+bajYI/b2/B/aGOxTZv2VgPxT9O997jVcbis5mS7Vbk1IzgmbBw4S
qLzQY4LPc4wlFxDJC/HMAoGtPCk1bJIFAUWEo9SW4hcEjvr2Ti2oglNfjtAwPoRExLt9+QKBJnja
VvieFnXd3EHFJqQzUQeOexGKJm3HXYCdVLslCzHRugIQLq9RMXrnXs6SXmSAXGJ8v/yjeIoLJXBw
4lKzhbuOtegJ4jQ5NJGA+FWnEC6h5Oh19e0iiEwIqtEqeCoZb8YQggqetsalyFDDwCe1v9ap/z4K
Va/buIT6Z63m6r8ZfycAAML2NtBOML4v3GEKdxAU6yJ5qbuDx+Ys0sljEr24HZ9qyhrEO9hDroez
2rqV54c06p55TKiGyNPFiYQNmf93jjBExv1WFHwb/y/wyEL5MmaFJFtuGXd7pej6xGeP2XHplwrG
AsXzA2OEGoGTyh0/hV+ErTjOwi/yBoUjP4tP2oMgA3rvaDnTkui1OTlxsrw5/RNP87Wk+oAy1IRJ
gSSrJWskMTlESiRwD2nYoTCvv5tEX1khiZbKwXkqReEJHkDGL0eEi+R6WXPd8iz4sfn77c7BIa6p
Jn/5zu1wQ39KZzx3O+twbVN+yslJk659IHv/qTfn45HX1a0w4fhthdRfD20AFZYTdLv92xVMo+72
DUthEi3+ZcLb/2LinO0hvTp0XeIjKnsjklgY2f79DRMhFWRqaAoOc8Uq3P6BevZAUQsrT1w36Dkn
ExoR930/G0PrLab1S3SZDJm1CR572ebRR7fPZ927gasDfRFbFkH041IKRac7Uwjw+jS37yGZxhtE
7/fGleOHm0n5/7O7cn9dIvADtgp3ussqZ2ulALTZpA+6PFdKRoSKnh/idUVCfqtBF7RCR6knjP+T
lXZOEgYSDo4msgOgKQj2+KvTni+RPxKxPtii9w3zZPEdYdaMkRha/Az7nnPxU/Too+daMGa9hF1B
OUJF3n+vlMRmg0EzIrrqehaZJQD2/fUM+bOLD6Fk+hYWM37utfzq44EkRWZFyfe4DtgWGYZhJB6W
rpdJQMjPQDlOF/gnQbrPSgNrrD+n6LydJSdlUggzuiMyeLx9zkIgqwYd6vIbfFEexW5Lh+AXY8C9
LkSXPZ26cn8ScGJKBZz2xIJ+Am/uiIzDE9+fDx9/yXly92ED/sau4UT9IOHiAQ4OBW3kYxIgM8S2
8dObbo3tT+RxhTrsCQii6wxdxrvDtm5ah+IxXecMPLV+N9g0fFLPQwMsAf9P7JggxeBiLiMIQtIv
oP4Eiji18x6U/y9iTKqr+QKWG7xEozAo+9OyoE+d7TsE6gTKa398bMbDVtidxSmyrGgmgmww9t/X
iCifHq8/RTDYXRJtaXEjqJHdAF7EYv/hpF7u6JbEaU/e5lBk0lA7EVSAru/Ni2dAdaSHrMe5HAsA
rDGdOmH339V1ZQYAcvoW7ZnT9tnIeDWF3sRloTgb8lqpBYufFShb2/VKwCianI2/MWXaYL2vohVS
jM1HjAJDT5aZhH7EiGskY0uOC89XBLyInLa4hO2pgH+1IM4QOP+Tq6jZ2Q/s/Ji48wEidYmNb7zI
9zHbORLFi5IeUWJvRng8XItnsb1RWMwHo8ZDT5MqucmAXnIBAQWow3RunZ2UTBa32wlssRPhNG+X
fPgr37RTi8nVG33XjeSuwSP7cx/FrK3gZaFk8YsrXHdXbVQFbnmhkFeerA1omZ6NqQa0Cc9O562r
6NE54EwBVBiTAR0KtCjn9M8GJWl/ixR/V5jtpuepA+F094mK3e96fBD5eBI5gAae4kkEGSrEBuHy
lT52yuSK+vxD6xRptkEi5IyC1fNLIPKfPPaug4S1zdKLzV8ba+M3zqDlk1yQ33j4Pa39MKCxfCkX
RDEZ/sORSVxtT8cxmNS9hxh7NOCGLwrhgaMzaAfq9cVXsK4iL9wJfbu3NYU2D0fQazcrz6/ddkt1
IsQe8/Cx/MMSiG7aBJ5yR1lU4ZDgD8C80G5XQhsMv552MS2jfA0Wui2XHMKA7+LC5cip5nEZ+oCz
I0y4nhWshRS56qsNIJZvPjuYlha4G0mbJsq7yQebfUtQtgBMKkRn0lIUs/xpOHo1WMsw+Ki4uqTa
hGihD02r56OXyqr7HilCjdm+dPAEh5swt+h2AI0MJuay6ztxHa5+vgY0Ztsh2b8GL65oOX+vJLMd
PVg2kJoSltsVxSCPCie64GqEmGvTxDdHCOzokH534Tm8wvMlx/XykWvUeij4OQNRV+DDurisN21r
ltvNdjdad9xDic2yzCmSn92i5AtdHcKXJRZPh6APG/LjXURSbqyPNmfHpcPZbtVbklEDdpys84+0
/MrCdx17qqeTdcvVTW+GlEoG92LuO6Gw8tKz+xKbQRaQWi4oQBCeEwD1W4yW6a5OQfX/hG5k0xnf
yEm5SUA6+pYqqJ5YnBvHakvcZkEQ3h6kwDhY1CfNtkmMEzRIw///NyoUTGfsMzU5c7RsTXTh7vkV
KWPKABcDXVyAGSZdMgY8dWmf9xd5iQ5dmQvvye7p07neNswdQCXSsKDHaW7qZ/jc8LMaiVfJR3Gu
TDTe7ZxjemrwOQ/w0oHIpKT03F7XWhhl7fgXNK0LCwHzkaUNiKxYxsOKo47+2dC8XV3aLhg3Rg1N
3E1xPkVCkRFgIukMiSUkdU4CGooOIQ5dRosGwWtIQnW1oFBihUadJao1uhW+ZeCPSrkwtuU50q8V
Oln5lUDqWBSV2Nxbbj9YqJhsRpIyFjznuD+ud7cLwU925JGPLsJ5ld1CH+hpGyK791hHrTBsvE5b
uGTmWREptUemcBn2VoH7TAzExzFrLEXoIZGF4ya+Oa0pYTuBVqc5e4xC4ZYQGljKIT2vEQaXBfie
qrBYt8LaRYHwUwSky69QO8MI/v+Yy7VRwiQW8hq4KisNjt3v4rhYBP8KLx25f8f6vebVIU9BcAV4
5M+p/YQdvMKUQYlKOuCVoKuRCkJf4U/uR2kRl0Ig1N4cPl/rEmCxrsX9OfAj3RhQgaHBcxXm2+8U
HpG49veRabp+mGn9v2kN2+dv4TmPeupoMmVE0ol48hYtaIivtEJjRPzxktc1uxKa562tg7iXl3qu
yBZ0uw3vF71uSbx3QeS2zm6Q6WSfsT4CsLiSrpVmx4YWHg0B8993zRTgjssTqNpvN8RSfzgpNEsl
O9c5rQL/cwgvVcLYiz9utX80IFOtTNRnso36d3e9Xew3ICmZEkCSyPYT3kiC1O7P7iX9z1dkuky2
2kJIJAYzykKSES8IdnEgg3RF8xaJr6EHXIGCEXTpLmmStibrELL+VOKU88+yLpMgscxaigElajtH
QuCsTqJnsm2Z1w2wugmdxfStz7GVYVjE/9OypuDOyV+JxYkH3Uf56oY/2aJl3eGztkVHg1VARYck
QDdHYdCHwvIPzIBDRYWPYg4YD9T6Y8tyQGYYe4OWY7UMZOdjZ6808wau0W5BtVevHquHCZafr8UK
DVBfy58xim+aLSV1M2TQyg2ik3q6pAXrQSQCHnck3h6QEIS/lVHKJRsaUZHIZsnmifYTknc59tng
rw0f9Mk2xIxT+OfJ7nIvTr1zRgndcWBbvcEC7NjVy6YHUt3gtX9iyWdCw/o242JkT4n7dVJBrCA8
etHVk08HA1Dytu+wlerNq8WMkYQWmBAViCYivgLDIubaEnoDPjzIgf1TS5nxa7knuN/FO2JC0VE+
X+uqFd1vzBsMHTQIoX+4IjuHE4969kjZbcMqKcFmKdRUTo3FaRVqt7sGIf2mVPKY6RJiGBxPrSeR
SjodQ82sDuK3HeHSwuhjCcTeAvXDn9WfmFbmSmm94vReAsJrqB5Ow1I6ngT2tFHFSpocZWcuoDqg
v8NQ13y8IwQ+5P7RH0AUNcD8ewV01+ghFK+PjxFfS0NdWwqhmhEMkKG7PL1n8qxR76P9L5GkvBdb
BXCQW8JaahDgHxnYJvJP4Zso84QrTNAWkeEbXPZk1vHOgn20+xueTJccM8Yn7subgTMdg9VE6c7+
KrZPUi7/Sxr9Q5RMEgaB0t7EkF2L1bajRKWSWdVqCE6gcbVjvBbl7rrsJaCue7jP5bOY17fqac5e
rKwgOZFNTVHxtk7E8MJFf9MIzMW5jx+e+BC3Uny1wmzqnl8DceHnXYgU+80JsiRPfwnipcuPrcxK
F9VR3AaXTx/91GPfvQ6wAdIt4/etYFqO3az6RkrMFw0Hs3FkYly4kBD6+v6IpLPalklytKfdLgky
k4gVNBvO5YzkurdRm92os+Ka+VXFYv/aU2J4fRJRAKP/wxULoDm7WIFZKyq03qFzYuS6TVjFyRwP
brHJYudOGdvluFrsDU0koEcLm/XTuCsrhfGfQ1mQUo3wn7V10nDsAZzrv0xH5qSNjByi4cAtEJ4p
oWrReVFpJ6Wz5WKPjMih3U486Q9HLs9A0U+AljqpGwHOP3m9DLspNsENqVnjOmq+jclzekW8Hvn9
9ro0KGNrdUObf1pVKWBvtQFmniad7h6zEVYHi0s5XjLq+1y+LwRLG8Gm+M1gbKPpMzndnTlP8FNn
nX7D26AkquK6uHwujbyMZRC8ht+HT1ynuyIt8/jN4kh6OctazkEJQu+5yiGNVqg+1tMwmED20iB+
Q6cfzDbhVgxnReidfiNTX68lay7m2Q9qRE8jqceYIwAsEgMbyrFt6CbEz3ew0Y5P9KNJo8Q/Hhqc
We5/YI0Q0uIwgnrWtbpcpirf+H31/S+gyahHqBEabb5OseZGm2Odqh08PDoanWPykdPJlsvp1ReD
W44gVEZ/53PAPl8I+B68yTSmULmhF9NmNnWiRGkhTAsUfYH0s5okimF97oUqBN6QVjnanFPBifmB
PIj0wayzS+9B+4geekOGze91m0j1hTfILc31hk4MS4cHl1rEHR41xT2sN9GiZkCo1kq7kPoQvyks
5zklWKB+OQokiWVyMk+XyTtuOE3qSL8uewGuGUMKGyf4mT2qW70u1ZJuw1CxWKdJXGT9vuqHsNDM
ZvzR34m4MXcdy1yPic1lFer+vJmcImj7/ZOID/M6pkTd79BFN+DK94jmIKx4IqD1lI9zStpgEGSw
d8US9IYLDL3mku8x4rNo9gBqDRHDMCFL6Gds3NoNBM7pL6+9bb0z0/NP/L3vsNNpK51l9Cy6uGbO
d8HL6i3Ro/sk/wBD+3khAFZmvM1bFgBQPi5l1YWaXFVfzInexNFRPMHqfegV3pHxxkGrhaN2b0mS
BZGoMzOa2TY6UXnjy50a4kMyQdG2G73vmPlrdBh88T/o41B6A3v8r3rt3FNZp1gYvDw/qnIUSOEY
umKvLl6YvMvfyOWc9NzNgAFjpuJqVJ7ABqG92fMHzyyZpTrcrGCWZpHKphJkPi1BW7+jm2pYDx9/
C3mexz4nVrX80OulPM/QM9rx14FGzGQXOwsW2NRKnyb1OrKBTDSR+q0n820bcT4/BjpwMEuIPyAb
61uWSmSx20og9M0kFyRC3uzFn1IdCb7i3xGwHrCwJqCVBX8y6xoyd2mPk5uel9dZfOzVFLBw16SE
v2N47e1jVlqM3pvqGA742H5tG/eQqx/W3oURNyVWVzvnd8tsEhIRUGsDoR6UpvPVcw3ict0UFKWO
M8FsvmFHQ861m/GHaxkPpBitqtGbSd/VqkAIf2okPxtlQd7a21lxdRNSPvAXfVftOewiU+HNOvBY
E6p/zNsTeNLoRWVsVbUoovxWj3L4EkBIzwjFC98sbOI7cgVJF1xE08lap0M/8nw8X9lAeyqJHxKP
+izANYEoMWLhgeoqIWrqMbHqM7HPsLXrx3NXFYohMKVZ3Neo6gpbxG4dPVSi6dms/6j2Gtm5u3cE
uxxeaj2Xkk9QOok3ar82zbhxohN9XrftRlarirL1k6dEmqFRol/FZ6bX//l3berOE0B9ha61Ej0n
JtsBq4rf3HGasrhjY8vpPup0uWVXePfWJb3MQG9i+iWjjDYTHV0cGLkX6W7boSRx+ny3N7mNpEt5
CILsfnar8/DfeMg7gQMT/SB3g3aqXLgyY0y4aEbYgRJced1fM8vZ9xZkCduB0l04JBY8zo6J03j1
ByVNQv7rv5UKHIXIRvraFsIBlImYyFHW7bA5C5QUs5BTvn4XpYfrQ78eg+eLYw2wJsLoYGbatSp6
Tlp614kukiU39J8eq5+cgquetssFMYqhS1jBkzzA0inQmnJpd+SJlX8zsvNBDm5XAtQs7jt5TVLq
PSkGQ26Qy8FJgILpMYq2nke/fFNAQDsUHvBzFsxckElVa64Hlt864eC4yqhkf949x+oEH3ksHV6M
LEnirDhxlnga+hN3LP/4Enlo0tMuZ0haL9XAblwYteWiNMoGi1L0PUUV4n8VttKyACmQkubmvUR/
MY77vJNR1rvARVjFgkoCVlOKMbLCGuwsWe0NW0vFWSzFsE51Wvmzb1D+AZBrE5iUjFd4a2KQB/JT
SP0mnICxpnz6o4oqD6TmqIoD3db8Uk421jyYmkRhkqNZFKkWaMr7pEcBU9fqJbW0bqU6aNXwiQWt
tMSNY0KpIFbajYORLiE1TTZLV6H5cZGe4lJ9wi6kt2WNPMa7erUspJXxU8ZkgfkR8Iay6eMW1hsZ
bUp/qxK7hM1oJNieHQQfqwLkLlVf+G8a+SMKcmnowSqx2hvIDlK479fWO/xd4gDPg6NgfBPTCeVM
yB+3zPfP6IKG0q9zSR38X1toHb7v5FqZiE3MUXTO8UMhSeRsylWsovsImhckDwnzy5py4IgXLwdT
HC78rxUAppaJesUEpy54ChFVX0+ev42cdMUzDim9987n+XJhL2l5LB0EX1IKfAywNeXvAdRpUiF/
KSFNvD9HPSK9IMj9NNgU6lQe25O0Hg64D/4pJJ+VqdWnqcdr/dkyKM7DtjWbcQjNo2ZhrsYLw/Ni
lX2NE6UNovg9PS8vL+bCT0ebR0qNdBLT5JaugZs20+iESm0EaF8PQ+aie5/ZiWXdbIWimvBqHX2u
IKoqHtxN8oT37P+1EnyS2QJJwibuthJlOXfk4OkvuvQQnlgtSAd1sJeJV4KPPtxNTpSVIX1CvwY9
dtAGfgDTBNbLoujIREDb5DA6WQakPZJ8aFqzoV+Q3IKFzBwv7e9ZruJnKFN/aUQgfrWJ4WRUirTZ
2kuDqTyC90LtD6X5lc/hZUb/nME/m9odx+MsZ9kfUDqJccVi4ybr9pCipUid7VOUaMC4c3vyWnQd
HXfaFvCDaYVlVXzpQlXsvs0CLCbG0cQvCltaZAjoQHfMMAedH2KJ8FTBveONEI6C65O3yNzn8Z2C
b0pMZxBf262ykob89R2sxUl9Y5Ycj+34hriFmg4N4wGCPdZ8xSQ3Hg3RC00EbDDZpcVdhZlk6x/K
4c4MoOCkUEpyi26bCv3f8zAO5YLhNl57uCmcSzAMukI+nzEd+1tPlvXuV37IDIdRj+s3IPf0B/A2
hSWoAO6dhCks+GOgzDwJaebaNqUSroCUgrRHZtsUmFEIG4F77XAzkI6RZWoQOXnYPyLLVIKL97Xy
BT5KQOPnI0uXuTm0uwArs31kfg/DVPWO34SbcOWTUDRd5YRTyGl6Z2eqnk6oOgMHTeWyl6cphD7/
2ZNm6Ur31tnR894QgGVSdpq8yUWfWI7NpqNkNpEZejhlxhinKu0hFJb0d6gZFKe5TFaVq1PqD2x2
v/wwdOFwmLDjcO8xvCbnSxSAuD96gFL07eM6PDejir5Uoi57qXF3y+nkPPFp5X+cGLMh5mgHsVKy
9ux8MRs7lZhyqWtiLe/gILAutAqM2kNnE2Xp2We6MP2AcLFjw9AEuXPlkNYKvzP5MHFe4CvbnWOD
h3ikK53yTHkp9hHLs5qCvAUkzF9aRQAymMi/S7JMvySh25Z5leAR+mzzTNCwX4ETg7FPkPi0GLIG
Pyq47A/JD4/5O7kOq6n53bIAVMz/aX0L+NXBgg4E9ie0ZAYT+4dGUF4XUXwQxETQmc/DcZ3/zSsl
nJ7YAYf20LwoPIUrC65GXYYqOXf6d9djlakGvUcP8yMEZvEN11rF2/kCkh3+4FcKLPCKONL3G+15
L0YY2GSO38I7RVBBQQTatY3y4wfRANZrK9930xDtnVwM2w0ZQ7Q4qkow24jEGXsiikRVAs11BqhQ
1xoKNKOVhBxAwDhT/HZavYNYWmFif5SkPZkLlvaDEvT0uUkPWRnkq2i6p0rbZZEcXQXy4bWusGrg
TBqFbS7/I3KeWSJ02yw7t1yd1SzRTaIhM4Xv1IKKFpjOSdzKKUBl8USMbHse+vNsRdv5dM5STO+2
LboyertdhccCVi/1jBKU6pGW+2vsEeAzJ+AT5DdYevyUydrjICyd8DxhM7DxgZhl44jfvdW1hhYq
eXUX9WjYafJ7YybrXGUnu7jn/F4qgYD+JBhrPhr3UDxiPc77y9K1g7yEwHt07ANbkBND+yOjSg57
D1phWhMHWdF4U3Oh6b9olw4DGLGeF98VbFJDlqZsN/bSrMbpeoqLDaR/t9Eqp1C3pELSpcfXbkv/
Gzixc92cwC+r6WUrtYNPYqTHtCPC7BAoulZoPYvAWpTMfrrYyH4r28KTGVqF1rCPnHJYOuL3enhG
+9uwjHPv3gPW18dwHvlG96KgaELsL/3ytLOcY3lUKoJbYkyFHzPYzPRNNrQZD+B/EJIwcyWXsA1V
bSg+ebzE0Yg4NVIHJVB7FIcIeBGwcU7/bBv3ZGdgu9AQ8Xn3RVEn0W0U1/6ytwJIRUMI7KalJULK
gkRLq6TERe4+7MjpiXforhmF4S6zV8NNbX8ffcR06iiv5c9SMeNEa75Xxe+IcrdpW+Nnljy4xzWW
x6HLVtqNGfFvIbahobL202lM8CMfQ1mAeIWd9mDfcN8MxmSBOgGyOAu20idLxlZADsXb0D7qo+Hu
aueXvFVBEHvG/eUwvlBKiueCRHqgpiGWGTXPW1sDkhE3yGEvYovSnM3US6TShOCZ7S0ZJ51nXOz0
xziKys120YVoJxb/BJ2FhRW+M7lC8kmWsV45razBnnWtDtIuVvtd5RNKGBvO1BaUwOUwvprQVkiO
azE265bo10rXNvM+Zg7p1tu2tpeCnHNGDzi1gkSQOAdvJgWFzc7e0u8F7ef40NPC6D0fiOv9dlGL
9TB/p0NsJtX5ugfXgXarQcJopoMc4uHh8MlGCyJKFpEw2oSPt0OAHmEaHY1eCDDxgORtQYcC2Cug
kd3qSMMerLX6RVljP1yk5daS+c4Aam5dexX1oFeVmGuZqDfV8vBAAN3XV91/B7Y/76aSOVI7oftS
5DPuj8OYpOzIs8Q9+MLdGuihrPswwuCjXvv4A5LBF3xYbVtv981XHHSc17xpUjLIcB2DRSYjzGjT
2cQXVqPKTK7d0EuhcMeec2dw/D0xuTw8ba1UoaQWf9/u6H9c2IeNBST7fs8SxrwwVHPNFhXNsc8I
ydNAAnCW8zA5h5OCOYUp+K3pz10HEquVzr1qXarb68l7qVFzTotpUa/aN/wX5T2z8m3g4V7FHbX5
armrGX1hnP526SbsDGgkEbVt2NAbeR8YmjhYo7XZNNqLnO6A4abE1+1qSrFMWCA7gjT7vKjTeNj8
F/j5aVceVCGB8KlG8eKuO23Wbn3qSJcALaoa89AdeVjb6x/W+VCQKjMKocjbiE2gqJ826XOdHH7H
HBTT3HH77lI3AvL9sr9gpMbsE+GDJhVvz2089I5wvEy1UJRnuKp53++xKpiQ/+0EuL1QJwR8o2Y0
kTMiwbuowqMcTNpDFL6jtzXX58RddZrc0/Ne8W8IEZm+vYe9A/SRzlqghF7UXJyla/j2g9jBpBh6
Tee3tFNpmRXacb22+7nNC5ft0D3bIBS+fZjONsRKP1AjXtqAUzJnoVa1g6z+ITNedwMhcwF69sZT
3iSJX4IlWtXWpieFX+GXQKNljFXGjhtsAIXmw4PPs2gRYh0PNgDA8rR2JByegCmPG4tbUVPWXVEx
scR+fELh/iLxMdKBm7/NqqLX44t6Nw5oe302/OI3dzbnuXUruCzdS7c1UIKWB+T7mVVyfnb75yU7
+GlafvDv+hTkHWkLr/sG0iwn51GlpBnV56hbjx15IQdH132ckK50klWqLISN8wO0x1RFLKG08kBw
DzpcCx2532AxrI0OBddegDwSWOscR2WDumKIBXUElWKmXVBYxMZnsgTexMm2oefDFKZrHCBnZTzK
A0G0Lbc2DJcB1tuldcS4lCYENy6J4zWIiHQZwy7KqyV+fFXic/KsMs1QHYbjMt8zfRzJXgHR3DUf
9irsSlqJ/us5FXsuX4sSe31oE9+pWk1+aUOK8nEfo0bn6k40AuBFP908ZE43Jx2y2KW5cF2LZ1GL
RaUs7OFyPsy2DLUi+LLRZ52FH36tvVGLaE/Qcr7RMTfgEt0F21PlZo/Ad0QUBBmcRdIDQzb2SMlc
IRFLDG6oD6R67MDhgvlhwKXqKX+mmuOaKQRrbWMLYoOF5v19v5MwPc540vV4+Tbv7t8wxJQr1w7u
BrnttyZ4TaWCCdoXRJiKkX/+DOU+3kErH5ilkvECjf56yTQoGnEWIgT/aTsYqpm4kdvZnrlRW4m+
2HyN0TGVlR65aQuGV2U8T56TY0u0G1quSD2R2qnDvUEaKqQHZE0bQ+Ty1L7gPyx1E0HlUZ2nPwZl
fZhBeXUdTCt1Jvqx0BDQsfSu2Hn7qd67BUtEdHWRw3QTXsJ4x6Xg+DtGGl7awmkH5Epsv5nFqWDg
aMHYvdHyUKcAVv7SxhproY9in3S3L84lPVIkLilzoqSjnePJYFVJvcIdw5h/2KFFntTrvMiUdE75
Cp3afff6WbK5q3U6dKs0B1A4/GGgyqtRzzEJJ0m4fRk316CUr+fwwEenzMWVm4jAl9fui+PYK8Ay
e01c59+FGCgq82QgcZoBLcXPVQfUEGxgrPEvm7zCr4O/0ZvJq0a2VLFagBaaDMHkHZ496C0HTEE4
NM6kYCNQ7xtyd5z0lDhzAtexl/00BE9YulqGv/kz7Jcmb2E5lLYhR8u84Nwxx3X9EnaZq7nUXsrz
/vbJZsERobU9f5pkDpar+VN/OTI/nU1/PJqccXOA35t4XqlZZMUVDrjzUzXJg4Jf3soyKLnfYYYS
bUC1zeJoCYVktiUQDSpojECwOsjTnozHVQbzBFCrv+RqSJlrkoa2zEhqfjTnI3NMSFFIUT8xnu8R
c0SK6ykbhF3eNpZ+6nxUQmVAINKDYwXzX1a1qKeFV+8RwP1rwmTCCfS6aj98wKlmKI987U9cbvCZ
qSCk2vQkzVOrJptTCsGjIbpoaL54XdMBTc335Qf2bITFJtXtEMkrCA8nAC2ZcPqsQ5L9yGQhvCy0
9JDMlSBIkBdUQy5Rsyad/FxBRLHiwsPm+49PxKyksvSFfDyb6AMQbR2+IZnvZjerOfsN86z9n7h9
IFwfsHjOPjFYYLrpj1bZsyl50uihT8GMMk6Ma67Mo6u76yflFnCPc6u95W+06spzd5zl08TTkdt0
+UuK2B5wIEhxqs5g0Fsdhm7/RHm12l68UW3FvbP+0EqzxOUjQmigBPPwf5RoZ0k4R4QwkyOb2Gop
zSPj7YrjxFu0iNoyuDM/L+TNq4qXwiJOZqdqOlEFyObUHH+ajGJiqkf4vCVIrid4BKLFS3EiDe/q
hL3tg/XVGka+V1xi8uKFCRX0f2KxhHGIMI0dvKqq1LLqFFdY/Bcc0e/POvdrycZySDXcAtCsTwBZ
0ElhX52Av7P9jvSDnWhr2rHSh2UHDJiMqky6QE/oK1rqsSM7fVxyi/HFRJCwcE6OwkizyK3Si9aX
ncYrcDvfEYyX90ADfTBXuDD3SWS5LKIxZXYHIwyKo2wVPEb+6346v3NsOZ4Bkcpd+WhNKDmb0UTy
ITVXpQ9jEyHbbecwlMqH+JaDJ7tO3gjmjznvGpcGCThI4nbYF5o2OT/12CzZwgwpu3CnEl2Cj48F
8zQ9CeNRhh6JCMGkIjYhMjaT5OmnUC7tUpHRMKj8LoniuOdx0u9wmWoR4CAEvsUKXrfHU8Dko389
tTjFj/ZfznLqjVeiicJki6ggXYttkdMWIpyA76Htimjg4SAUkvZZItZvesevJrH9diUMBbStAK4Z
/lK0RQWiLNRxDgMamB7kdiqCeovz6o9NGoeIVuQo67zhqlCIuE2SA1A0ORsucEbpmIgSMp/V7jrg
71cg0Pn8g4UtcRnfk+qKSi7dP44Lgg0HtzK45j6hdiB4TyWK3CenvBQQ4ptyLMNZHrl/vcy/ZwJq
kuULX5kr1ij6xdoil8jKYwmMwRNMyrEZ3nGqKy3Jg/k587jQIf4ZGJaHnAo4AJsvQVyFJLBsG/UY
4Xfm3vwXZLGQLVGXv5uRaJw1A2FQ9lrHn0GLWgutPY/DnRIkmVyAOosfZ/yt9HJKZ5WnUaNFRtGE
bhHmLZYYMyg+iHwlmodLlmJJ0L2Ls/lQaHU4sAgxCZUxzyKqybPoi97QHg+dnbuZ0lLjLOogNIGG
ydfhxuMBexaB5tW9dDfm9hlxkytJuIpvJgk5NGhcoqNF4m96kMj1wSBG1wRC1MirTDSVsYqwXjvG
MydaTaXN5THfMPqOQv6nguDs4crCT8uYnBvB31wxY5mvsc853ZE0zmDhyDx5BKaeJL1GbYGJ21nA
TyLnbvGMfnhYkIwGXjeShV6oD00SmAXaRBclwonn5+25loAjkUC2VQ4vMJ4pYkbtnt1fYPbcMsXQ
zS5YfMvNU8TM0eV1KVOy+otgORRwgC6ei9sknhCXJmJiOYRP52WS1crvRClQAk/2iAQyi/w5DqA/
D6ZJ/PMQ+gieUzzZjRgIeGGgTLag0mdEgpng2oKi4m17JCPmMc9WWWevNn2gdLr8snq5iXZYYQ6k
1AOEa7ySOYzPoyffLzeT2sDBlJ5H1L8Zacj5PhnLJRvy9sHe0MdrmfTcEQfNr/vNpUPzTf1gOcgB
u15REvDetcOgwQwkYt/NIvSE31HlCRhzEtjauP65mLCc8RliSPEWeuHcs28tx312ltuYOZXF0XEv
xaWCfvmfLFurUwIPTiXljjVKFtdxIKH/RvgCZdMKmg9aB0ywa80GzWCVaoPEA59Bb5kL9NzHVQzV
RK2Pq8kEDnLiLEZBBvIlPtTSy1gXBIovIVfW5dyA2h7gKnq8XqwEp4Tm7GkfdBjHPlTRg2nJ3DNN
SNJ3JFLJjZncc6CwF2/P/c79z8Qh2VfDpW/sQuv62ybaKia6hapQk8MBFl0YHh+uC4gVjzm2Yd7O
8qd5+ZkaLjQFwlTISh5kfIOh87VrSE0ZdWT4rteHGTN7CNLYApluhE9Q8Np3JZejCSmNBrYoQeSF
p1e53DtOeoCKQ5/1K1E2eAlI0tORJIceo7yUfwe7BeK6/JmmI9P7id0HguYKrfbvMFF+eaZlGYDj
d8ZCT3RXqYKLavjwJ6R5wCFDAVL7feltoeuMi5jnG+UXLBO+j/76NLVggmfSU5TeD9w7SDc5/LEH
3UDOYsQF3WLtqT6nfMOgvJzmvLcmIH+PHok3V2kHYlODoimiAHmU26Ba7rhx0zlfzMB1PuHecwZn
x8N+cUK0Ozdzf5XIqkyU6w+qp7PL9WaTMD9ck/8nMI47HDNZWgzUBeYQrA2jZgccHcAqbHDvOoMg
8Z/dscoyABuCk4GFX3rRyvzH51TRHRnvhZI/5TlFwrLoA/TJfSMeRI+nl2fH4iUIWf75U4nr8ekX
qirNOs5DCKIQbZRHPaeVb4IayH7mTId5+iS6JRK5i45R0URrE8+fW7YL7XC4PrVTeM525XHhCRPz
LUtC4z/1gAfK7QmyMsMR1T/2lIy+FpjGsuwuPnC+0SxSJ7ueAGcE6T6fPs5btNyqq8n1ois/3LS8
oJpXcEJGAFKi9g7ipjFKncS+381tbRXcRnaBdElMQ49OuMK8cK2v2qT7dUGiRBJn9Ng7jGkDWufP
z4kUIit/g6POh+8v4dk8gJyc6aq0kUiBn+WNJI+/0Mkjc3sX931M0QjbfGtLH4CuBcttuzQCemXp
3TdDk/bVzYgPSB+tnOgHHgmjKcjMevc12hrN61Z4CDuDe1HxWXPGs+Z+Zj2lZYhuXXcD8tE5eAm9
DUvO9uTZyf/OshEk29ONEB98glI9AtKWucFCodPWFvzDOGpA8M0rbqe2VdoTmW2j+pCV3GCP0TjG
YqULJgv8mzsvHczsxanEJncXrfyNcQG8VOeSpT64AeOI3i1AAS577i8/2DO7kecyMOO+MdggTzw5
pq3MZxPTc8meDmBzrkhDilJKh4OM4ik26+9ZbSQeXRoz/JcQG6qgg7NH+X+gBVCSiV56AIzwlpET
/sdl95tXBppWuhahecgfPb+yrZZqxjFQctTU/ZqdsPpYHUPnKJ3a+SH45ebVXiZxL3L1A81ePhMV
MsyC38TbDrvyP4AKhMkiVr9psgLp6arfiGQzE+miKpk1cefly2CyBnne7P7g1u2uaT1ICjmvkz64
tyITR7l+9YXZi7LhCrlv/NG0ugq9adb1mBFdPVzLTpblmD02GZH+JJ+CL4peJQeI9uv7nnNfH1qy
S0MSH89BGNY4XqdIup6YOiyzgxAI7hvNllB0omAAsEuvBoJOt11y94k2a10pPXUzFnAEzXVDCMWX
PMc1EuZVYZR30WIhd2HvRlLKNDbOUEUAFlKgizrDnjDTNjWl9s/kXFhMCClikHVpR07cjfiT2hMU
9GpNbvo2ET7wYFxEeyRM2e+t5H8K40c6pRRF4uB6Unatdlynd6uO4u5l3xcrqnocBT/NMekd1IsA
B69K/JP2bbiWjDPCKm35uIY71/hxEvsRP5Y9GwHQlipljwSJCp5/zp5ToBC60yl8LK2eiHS8U8ZZ
2SoGY5HgeaZjhY+1rP344BvKwBGrpLZxUC5SKCp/gJxhK5RMLurFO0PJwZPB4tlFwSKc8MvRbl1F
x3Ez8GOqfxQ4Sl/hqsNngQy8Fc3MtO8EniRNv2pY9IKP+Z2fjcg3DPK5A/Q1GkbEAJh6hM7ToSA3
r/H9qB+QB7BU+9jaPZ0MI8MHvl7LjGrezW8pcg2gWfXrrcekTKxeWzwWfcQJmsOzkyDrnyWfBRVO
myzo7IgLAILeh32VwCvn4PAUXwqiyeTjCjiY+VIpF4Yl0WErXYsY4C/x0kfGKzkGR36hTNgW8vRd
mObDKfNR4GbM4Xp//z347teLP4FFW2RB4M6LS/tN4OWsD/YZfhM6nrDC2cN5rVejn7flEnJ6gc+Q
V4dGWKN2GU4gYWZC5DIFfrTRaGtV6ZNVV/JNa2mg36UIsd2SyvVqvBztEaIHDkcP0+aa7FyPUU4h
qRGSNbUgzaiWnmv3qAKKOkhxPVOeA3FVVMc0QbWYzekLtyeHB5CLGYO6UZG2S2Y+/PBwy7JunqC7
nYkqJ3D8m1yfbo87zOZgXGagvAgyVxbCGIU4YBC94I53u+NsrQLmt0ZnU+i/WvLAElmSU1omFKn0
NhZ7YrMkJiUpuIEZzdEp7k7ek5IDOncdQBdePsRA1ax5ZOFqT1/9v+VJI+OaNUTskplc6BFPAPO2
QFdX6C89gvMNaOw1I46+AlE8CZa5VB7ShYbG9GCyEP2Snet7N9EvAZEY9LtAjPBFQ0PDiskaQl2h
Gf7YiSk7836Jh4d2mX9uBYiPKjz6uUujpYWu/XQoR/FpVPQAF8BDZeL8sTgrA1gd58XXUqrMVspx
+rtwkJPgn9mTrhUyTEqzXUhRwB7bUeipxNzAAhpGjfgTQi9fRX8hSyKuJk+Fkx9DZL5t0OTfakeX
rGJg+vNowzwfj7nyJO7BX5iUOwDj/XB4qT+aI4jAzV6e59Z7tYeo74sTcfNtVpPIKywx1sJl+SBs
lTWQDbkw/6Iq+m+YO655MjAO8ZNCuagX/UR/y8/GY+WZWcbCUcT3JQzkwzju91MiJJ1FdF1qz4pM
JTGahGxbnvLRjhR1pE9/OdsDmH8RPzRvZhj83l08UtuJli4E5CANWkfap8CAO1m4jWRDURd5C9c1
EZ8fCv83orXmu4tiYtCNInJKrdNT2P7aT+NoVGrlNibbd7GpeAY2OlpkInI8fsHwwMZl/zSleL1b
dgNHMapLiEMyEDvqiYV4aRwQrvyCLGI3Hwj87vQDSOKEfg4sFJuFtlYZKfs9PhcJeZo0MKk4oGOU
YMcs21BdFU9f1Ma/KE09iFqOR9axbEFPN/EkGJX7w98j2B6n9Z1HzXf2wwogQMnSYlwtDC7Em1RR
HlkeAZjYBvk8Lm1fVVouACx4lA5jpsKin5c+jLnCKtc7uDoZVFvUjlQZ1bYddfGCw5xuHFq7nPGh
yekw3pixJ40NsBE3r5wPIPAhjpmWkkO3YcORZ1TVhZk4cYQAJh4EeSATdOP6kNIXSMyEPnthkOZ/
X897g6QoCm5DZI9/BdGnuryfNjxzbABi6/SXHTz2pTejGOigG1pfinM8EPQYjf06z2lPwD1MvQbq
dg1bayM6YQDcu+OdLSWl5YNxMMmaDqOjhE30xz+CejxpWLJ93IiDUAVbTxhdx55htNx1hSYYoPiF
XR9pPzmTHvRKT0tarpAkM4hN78bdVBS4PufPNzpRSxwf5bPvBr+b2R+PmOLJdwkfKKc4u13kDF1U
BdYpislUlR7w7xk2nmfYnzVASXaSzY4wytAOxrWnWrgbaaapNlV0P3MQapZxs90ca+Q7PRnfc9Mj
KITMq37REhYO01AdPRUxIftaH9sFOR/jXxWeYJy65nyVhlTlqPopx1PVj7DGIGosTHqHd8ByE4YQ
IZRYPv3IYclZg+ES3WZadbfMDjwqia2chfQsNbP8hNYAJdYQgvs4DqSWgPwzggNoODXL5+f/0jUZ
B3fMEVmS/eu7/wxCG7ksNxl+NKzMrKe+afprC61Z6MC+Wp/99HIa8LZgVpWbzaXt+HktUPUJ7Z8f
2YeA9Zn1caFxs6gQFJGIyrwQAdQBC6ymv0HIGGIfU6Ms8OtEfS8FfUa/rq4Pxj5maWsH5YVM+7Aw
alffBmskCQWenBFbPVWWqQZlZk7FYjBmjvZdZUvZE05nO5Zp/f+txPsBfRsNWCT1OjF8CDmNVBAb
kUsXxr553gJacQjM1+CMuEHXM6v1mF6h7QXu4ZgJzDKDwwyjsTcKsegqFuLnGGsJDvzSvQ4N6hec
JvkdUxVS21leP9mXjjMiSVn0H2F+eIyishxHogDGJZK0Aeqgtr2soc2PO/YkJrdLRDN3HCAYGEjB
thBIPc1EvWjhYpIvPxhtOolyP3hIQzOeplvX1ZN1Buf/2aFpfYGHquZqbE6G9bW0NIF9NJT4FHt2
PQli3KAo9YG1O0xJw2BmbbqO/XuQIRXgW+X6d/+UMptS6oOG/nd+ykcqgRP1+JFJEPT+4DwZx/nA
7QKE+8h5kgvnDugYFBupKJewL0Ffy6V3mkHUQUsiguve18QkpURCkm1ZrsgfzVX4um1z0Hj9u73u
9LNo7PMzUzZhKBh85+3XmCpdtdtu1fIAfN6b6ZdqWsFUV0fnPTE7J/cCxKuVP/5poFIpxFetv21/
gM8wryup+XEEB1tEicp5nlTuEk3hSbrbEcRiMtpmrowAsoqP7mCo4vhlwUXcb53mE0kspncEek0T
+2IfKOd0p4gxPOnVSWOt917A4ZAlqk45GF4cTONTdXgNmvz3r6ySuYcV5hfdiBWdZ6/UI88VyOaI
Y94zdIMzGHfX3E8hOaYtZpyK6tTpSCYY4aCfThEdhZZ07xqU0/ZGjjZ6sGCMReGCRrWG6my7vveP
Ka6JSO4S+ZE6fshRk0hQmDk4fCRLsp0L9re8yAf1Cd/vUL+1LRz6Plautd07igJfUbkHjxr+h5LS
FnnRbyhMEHRGL8DdvRooIO8PxlA72KleK2jCf1D1+Tq+HheCfw/06SZvQA5tLCmO7t5PYxg2f/64
Lf6vkgpNA2Fvv0pMkX7AVa/H9wMdTWpvMyb1vIkp9aHklt9fr9XAvZ0UN5cJnVMdcCfTEsGroYE6
dzdOmnclrR+MCOGtk9FgrmsX8+Lt3MOeojj2n7bJAFsfvSiYbquroyCheWWew1HR/17Hjdmx73tQ
iCcn1sqqmL2bqBIe26Sre0JpylQMfNJe4As4w0sX+2uK6CIkLaZekstWS5pd/mORIZvmvLnZbhdD
RRgZG7E+idxqIG0rmYZyNkIHA7bdFG3Tob+22E6UYCKx+x5fLCt/26uALySlZI3VX4LkYhA35Yoh
V+8eHP3YXguq1ZumQMcoPwzzNlihYi+fJdCWSuWCRzcUmMx5f9YIHc/enj/OW9ZbMVDyo42HgKMo
FlIDyuMitNzosfXYIrkj11JGBOsIpK1GPoCHTge/pT5OFECcfbnsaIJgy5VyEWY7KBhaiqO9evOI
wmycinvFcUh0sAX8X3hWz8cnKdIVlImr3hfOw3zn89rprworl3E6nonnUM08kWk6wW406pm0pU0/
94Ms/FcwI4GvsaTXiVPaDfo2brtP1g+ObgSDqxXO7IlGv1D6ypwwloqB8bbyrWXgY7S0NA4fW4nr
R6Rts07LrNwpcCIaOUei8oJnYpihuo/1GuYctbZPD4CwSXWT3Irv31y6heXvwI0JucwBti4llSfr
HR984QaGCacjjzmGb2zLB634br8MJYKGiPkRuTfiQ4CRjb/kTGhCcs9FgUYATcNj2DLvu0LLXGJX
6WNYPQoBfvNMRf8q7SbmJV5ZHZE2ylF6Ooph1xz4eKU3tJVDxe1H6f1mcNOx+4ziaq7rjI1FAJwZ
zICTzi1Y+wQ4WCR12Tp4HiA1KYc+ikzYdtOroDDVfatLWyPn//0IKiP2ABnYxAy54v7blQjezXqN
2zQSphA+EENh8OE3YEcOqYearCYMRNMpqm2piORSN5cH/+kZ2QJw+3VfOxsGrtWhmw2BryxPl40x
j/3drvK66om4J9MiSGd+8ID9moLD7fim1idINsx5IBq2fXI9r9QsKkHGAHgdtZgdj2i2A6+FZWAD
C4YOA29LBTjBGGXwH0R5/+bNfuimiGHoGNU0yg+pkatISYtNCzh41GmhN9lOMrN3LjZURG7DIfnE
WWcFAOGzr2hwcpDGW2i+9UwHkRgu0Tq/LmAX9qZuVc7inBjxT3suGCDsprCNFXJrnGgL79LXgKA7
+x1sZkTrtc62Ag2RzYvupBgDjvOqLIc+t8Lp6dBB14tVAW89Ss3fQ95jkxutDC4usu6kCODEgTYW
bYrSpJZxXyB+0bAF7C5AXploJg8+dCmWDzX17VqdEir4SQ9LjKmPOvska6H2QLSRwHy2qiV8sxfb
AzkEb4VroDeYPLGphgLHxEPp5WT9tVRAp8GDpEPSfJ/fqzs7X3cQlFzazHNhFawFNl0NRLHRbQBx
HSltQjfXM6HNXd3QnItQCwC4iDK/iWGa81/H4oG68NVp6hMVJm//hkiOzVKo7/Qtm+utTITM9i6l
PqBHaQM7G65nhHillOUlunCEHLcmWJEBLww58ynCRXYDjbgp88k41Lzi08f24hEjI4/00FKxzN9z
0IkLOThnF7+7Sxa3sKhca+p4FTbSNyy0b+NSkGPXKv1WngRKHKnZ8GgIg5HAgUtlNNsBbozUye8b
hetEZ/Shsf+yIVzj5fAmtDyEamC2iNeBDF0sbHUTqp65C2aYyvMqCut8pcR3UegmWK7FWgrvMV26
7+wY1cAxKoTaSuSnPpVDUStaBuQkbyMtPkWmtj/lLInbuir1Hor84MY7W7eJQfVMhHWfY4WzVQ32
BBTU1Ob1FF+xfaOsyl+rysLpL4FOmL8LMQjmmQRJuUq8fMwVjNOwwv3kXRIe3d6j/KRMlxHXaISe
WkqGOXoiQKSeUlQL0YujtANQ7SAuX2rPsf8gIYmgsQs6oqke3+VqDpdPfURVgXTfoxEUbf/a59Ic
j3izyFsJga2IQMAZUF23Pc0pPwyiHEjId1W+o7pDpe3v/yjNDhwv0VuLiWMcDmn6glEA0nm1yQ+h
pAhbi4gQ0OVu9NSxs3KMI7adGI2QxSykQUdKgbCWLLF3UJKpsQLL9po1qgr5QKArmT7m4Be/+JWh
i4uqx085HcKukDbHYwbNA884i+Ho4HHiBuLxOpmJaXxKzHPfVonXs8z/e6UQrSsuVTzMi+/e5CB7
SOh/bfvj8sAlhbpFt1cTp9TShk7NZbwLreeQne1MLsCTwwhuBdJA2wjKxo1gdyBClb9R4GMZJwzI
ThZdNx/xkkt5YqkTHOXyUzheoa8bMAAgtP/e+KOFCIrtY9bi1hHL6zsTjVYNW/jFrrUaJV6sZVjD
e1iDvnOkMKvJn1MWOWWaudCAJOlKG04TZ9UYizGPIgWGwgNfB7yqWi6k54sdCavfgloCq0pe8NIz
vjmgpVPZQZpJdCJiOAs1MMMmOiHoZY0R0pkNLeWF6rkUYgGAHFWNMsG4UXeA9ZD9oakolGTnCgr6
/rBGKwRFP7zsY2wEyxaK96JOBhEx6k/VUOgM9EZaw2s4Wxn4tTGjRPrOtoIUeZ8KO3UufU44ua3S
NDQhbI75JRCXjcjFdMdM5cmZeeUSjYcc/mmWExWttkWF16C5/wrCyaDVHsRKrXBivg2fBi+Fv4KE
vPWuELHQjUPenWrSgN63MsvyVUR3y7cOqOJAcca3p9v/J5bLjsuzR3fhThpNolDOqQad7/EuyOye
89PpqSOOG+cYCHmvwI3zEK8EEwljRlb4lJ+mIMDY+vjVYGNZSF+EmAOQvRzchONkH2pWBC9HP4kc
kcR02eqVBqKa7KyZEnBAjRapwYFeNGDm+RjbGrU21IC8zFUvDFDlSB7sN6SeAkj8XbLAaelXOM15
2giNKXtgQkOAg3GUxtNe10sHKW+UWj9cN5qvs4UGEvsvY7gszbhEFpIvC2CMbkEAGL/mqgaUnwIS
8g1qnTu/v/9rMCIIO0EbyfjpeOOsNvCQ2gCt2vt2moV9rca0/c0r/7HQxHvyBEx/8K6CKkASdEM4
thlv6Ix0KvDrgdZlbsTgDxanRP/R7RzA8FmarjV8AAEpFGcJBqWXX+/2LQknnsmD0zoov655p1xJ
7OMXdnyo/Jy8/glnA8oa2I1PKUtmGOPNRLVFKHGolOUnZXr2S1amxjiY1DM5HKpZvuMktGHtOwfa
bFVqm2zzo0t+Y47gG+Kx0dkq/Csk/whGtHfHqquq43/i2QYTSb9TsFDwp+h3wpHpu3jen2MzYc3o
3iKASlLzp/bi0OaBPSpC6O8SRf2xsXIu3PLEumJWNO+oCzeXugHAJr6hwgeyLlC1mK4mi+X1vbet
0GVx9bwGcUZEnQYc2L0AnryV6f8hCg7aWxnePikOyPpm2WAjeLj5w4E5TodBA9dUVLmYhNSx4+P/
R36A5WKLCIJUuieXW5swQqb5BYnOKUV1xF0j9kt3KlL/hyrdu7iKwJi37K59IiAxKdfTOHvmpzyX
CKnmaeubOVvE932KOo7ipu99srcI7QvxzA3DeOiNU5hO4ySSzlAJg54N5FK8wBoXjHoiu0ok78J5
H5by2jECWldalHimqRbok8cV7BfLoUVyGb8wu5Ackl0siYtUSzLb6QOgehq1HPyWQiyyxuv04BOC
2loYYyu8IZqmWmbKeMz5ohCeLerVlhSxSeKXRN3mejFAs2ukGGvpWaay5ibicuIWtIXk1k15EHvz
wWT11zccTD2mPElMratCHIiIURNSArcpl2VG/JWr4djKAu6RkmCTlyK+wTVPepFXw+pqAwPRKm6V
qJG4G7yQmuqprqca3UoPU0zj7enJMGk84BAObR4fuUpQ2+VGQIBnFhQt/zbj91FznQlQp+CTchdf
yNnsIaOLUyCtnlaRtzoRdN6MA+35d0ACBnR5dSyvq9pNrtB3NNjHhRmauGGr0xyHLqAHIVJoncT0
F4eKOIKKVqMuq8sNB/jbSKhrl4dMLhCCnwY3sfJ6Afqc3W0XaMcepb0sQKOLBHIiGp5bnawN1Ta7
If8o8q8ix8z7JNHuUmJ7rzCPb8XQc9d6M2BTe3DyoGQ7/9XKggpLVqmd6ZfnVZo0CdKRPr6f+hYe
7n846xbgjF4NPCZQwYRa0ufVespL9pY4sMkhi2o83t/OOr8sABlccJ6094TfkpgJLkfrIJIkPQdK
p7sx/S20OvzKtnWX3i7GBS/pIPAYVeQ5N/l0AhTc36TKVXr1d1BYCqJjtTXuYP21U/OyKQykA6jB
N/UKsXJDk3czQu3kcZz4tcd1b5EwC8iDDFSXLVKTwITSU7Ats8tWUvrWfYwto3CzUAch9DQ0Ag+Z
VMJWcORw8FYQwn7G2dUavA1bDY7EdKyoMD3piAZkkIJ3eHrfAydXKzxaGS5Pcl7RSZs763jyKDf8
FGoVYELr1mz7/g6FIIRmgJCzg+QlQdGh5VRjANEUERnJnP2YmzNxnE1kkXqN8F4cPgZ7s/VDdU4r
mmbJ2j/1NJo2WJzC0nLs3l7IAAh0E4GYiPBlS2bx1XQzepe1Z+08MQdTGDbi+YAMYPWe926fdM9u
8Ckb6Hlxbsb0MfR+B/RXSFPjwyrIEsBYmhmFzqW3negt+smGoIgY/0ivnz0PirFOcAysQB0REUzJ
btOqSQ+5wQx9/biP0UOZretIK7QrAwzdAJcvpHDb57BEu3/2iYBuR5Z77XLVq3Q/+e+sn1B2A2C/
w8y/PlPBREPvAS1N5b4qelYTnrrITx0MHB+SRPb0z6Sh3QtItHXKTNILA6PrrCn17WNZLVNmQ2qo
p/KNKbCTPlZr/VhdX0LxSxRR0q5ur0FrHJuLH0zc0U60kd2t85HiQ4lF4W9HBGTJ6jExOW3vszfS
OND6UTly9EwSMCUdB5hD+F8GNRl067esgqf9ygUmRuqrQNwEzCe4auHMBBPwpDMTXWGWNR2BdVVN
rPo4SJqBxx2d19Hh1tK3Zk6/8RDXg8YBY8TG7tKF4vka6xGERSwlkahAF4RHRNHTyKTCt2q0BWm3
Z/H2RZyuIxzFuTcY1kl3gT6z52204om1OicFv1njLKEfnF5GI1rvAhhulIW3JVFBZs+B5c78WzWq
l2mycadw8WKj5JpM25h62TA4sPb+Ub/hubac63wO5ICGjjowbJD+MQLGYyGSQHRpsniD4Qf5X0/Y
i6Slt/hHJH3M7ObZeAV7rQYU4toajBIMuN1O/Pji8FRawiycOKmq95cEawLEFgh2lcukleQSXLih
NPmm5UugdkFpO1pZ9uLX20F/LVNrwsOIptseYZYFNEXwhA5khqRky3zPV/ZftHv7JkOYAF4q/PuB
TTMegSc4PHXZOCugSz0fTNtGInTJ7QxwNYNQBZqhXT4z26LDdScsy5T1OM1ajMJNoB8Dk3c++Npw
KNJogmkYTJli/HyfW+tQnv49zHry7q3kt2E9U54gQkGVhj9LXd3D02DeCZrOvgoXZ40xdskloXdT
VHtvVEjgkgnf1CseLrmP2cibllCUWHi/ls47eav5mBaCBES2kB1O98qPeJvzIyMjSYU8F7VyAvbI
z0NlWw4MRLPi8Kuf+tn9MDCK6VEB7dmUyNyqaCy+OgyT8ISRqCPJsFVqt7HdBobRFHddQegYZrmj
xyg3tfoqf7JEZbXqGIJesCV2UNopFuZQdHBaagnlyWSFKUk5xwQkZttfLaDQo2cBKvsE/7II/sl+
VLuNgYsnsYWtoWLitzF3NPGgedkiDJMyOE5PLWruRutDCYH9Wc9rdWLjqQzDYxNCgnym8zxHTq3e
yGrItkfoTQGfZkGIu1aiVx0ug5E8XPZ30vfFNADjNfp9XsvK8iXO1p2Nf8fZnfIE1uaGBiPafwy2
TFY3tXTjM32LHsD2+e8MrTM/MCgT99CllyLN4o6jyh/ds0sXe6G1o+A7VuWISZs4xzySb/Dbnk8X
qeiKwakep+9vZf6GeaezPZpVAdYeoxSauWgkFQEtvreTPNx0C90+Y36tXyzy9Y69P1wSYJw5YeoB
7NcXCAgvYuZT9IKni4ox/XryiQSUzyc60uKLIF57IQpLr/73Ib1bZAa8c/8tBom72+19a2kub/55
ryRQ1Gtiv0MXxagO7Plj72hPq3hVIt74dbvnc+jHgDE3HpWBJvJN0iVHWK3ELVDSuUF0WcedDzQ5
aY99LjC2GQPuj5GuvQk7aHWtnhODn9V9oq5j5lH5GwsE2EnyXmoxdgJIET9V1j56O+C/7O3hYRc7
DVRFPFqWyNNr0Ad44Aatkhco3+H0zn/m3SIc8a0+scpu2xM8P0Znugp0HOfoMbAFA2RjnB9SZNdg
6sBfZwaX3gIlCWAVG+2/q2rpV7RCGT/CfO4fT6YUWfh+ZjoAXc6Tq01JhGFEy76d+vF/j2KWKHr+
F0GTONWlX4XEkoFhSbgxCnmD+0XgTaP2vkYL69fLN4yXbTRn4BfVFic1EGsQJVBQg6Zc8lW71FVd
b7WnIun2HdvBFmXDJEi23NRuQkwunGoq4Q8MYFgttpqFn4vrOFuvNALuJb969nSCZiLiiyK2+KsF
0mMIzXcVVk5IwdF27rmD+rfdI1c2olDEl2jQMR1W90P/n3Byb6AAMK+xn20L8hgtV1lx+ujenePn
Mfw9SjGIjVHMcnQORMRDIChwLTheVjTGardT1GxuqrY1+wMGMs5Xo/I45YLqJ3IHMv+2DcTxG1Wg
9PM6dCo0mhZ2gdrfEX5KAbucpX/mhT9OWVBXaEg/GgDmrd9RQKThg5thQwiIV/6+9WJrgQM8OVSS
3jR7tlLgNiEjgI2kTJ1UDC9IYqNKR1L/4+W8jjh3ecKB31gy16RP11iOF0vElss2Drmd5glSbVhH
o5W27Ot8MKzKsg4v5LGgjSD9vstcVipiYk4fwxZJkg3b2k2Wc2wozAhMSAghA+HKAU6yrdPSmMoK
Wvhb5m0DHTN3iMBor4jjUHC3Rs3t25Pczrrq4XMV+xMBabwYouEeoa7IeSa/R0Y8UCk9GCdqBxhI
QFLiMd49RsVTlsigfbWL/3VPnlGGm9cmiByiaCm7vDC7dSX34WdHOsRIiHxsN3r691KbNTdR1xSV
0HKqPhuybNxA1zCV1bErI6QLFCEWWuq48tLUjMFi7iTfzbgAsERJh3VoqnhvUxwvyIls8OvvlyTh
q9nD/G1d7+hdTYWM/M62EFjfAdboa4CuIsplSbX3oU+KeiBxCkd3p09Tz4el3DHzUcPaJGpah5BQ
hrV5mlYbnNLdpalXUVs2t8H6RaGPEVY1EygGUiSQhWoVIJhNUCjaFE3yyDn+ws1bZxGkaHcB1nDl
/Y/2JQAGebHmEh9wTUbA0v6hlZw7Hy1sP5QDhlOF+1OHCTP/bBT1+gNzsjYongamA666L+3It7X+
TydSQ5JqpDN36Xtd6jX3K6b7r7P4pQJfeKkL+qhSKrgj9Oaas7l+m46b3k0j5R3BlUbAKnisp17+
RSiVk1m/5QOAA+qFBEjtoteQkSzVpQKji+gNH8Kt0zSTV+uUOktoUb0j6h/nbvLHsYApFpewDEFG
Blawkme9vn0TYTg3SPhaYk5Osp4zy9vsaXgJwhtYjbyth8UuRY7OB4VJvTVOFHhWn5j8KSLscuyt
Zte6UDchgd3IsihNo4IsbrNTJwXbAcTDHNcqAWbGqP14xvoOjAfTD/VAequqh4h7d7brQIKiu/CT
M+c/+OHWRL4Mr8jXyPD1G48m/8UwiZYDtm63an+FhtdY7OBAgOv9jnTAWVfYuBxl6/NvbV+UHb8s
4gcmye3Zz1YdYP5nLS87u0lIIYRI+lDAIId5dP5bDqsPL8Y3TIHwOQwmZA2mtEDzesSdWD/0jfE9
TfFzCUESPlDlT2cvZ2EMbOm7txoDYwpMvs0utNcr874+54kwUidnGLmUp/3fJQ/Lu1WvclyPN0Xj
yPJx6nljypheCoYewrS+C/knDUuzQgq7GgOTKKaB1d2S1LtCIWp+OWYbC5F0xgYXPISCNAdEPcuP
R0Q8xnVzSyl1otzKgR8xavChOccn1RmGy4I66mI8ac+YNyATKJsQ+aDupG4TPmYntZnuS1fhc9wK
hwU8sltmmMj+IRADLeoWbQ3K1xJr25GSW3ZlFI5ebcdyk/iXBFvU9A71aLiBXhSOgVWjW0jtRj19
y+hc4KIMYeXRfJ6gHh8CUsCgVhEEm05OSvJWvvoPEruAuZ7/ZMzUV94X/z0gQnrdY/2K6ItT5LwK
Vn6n14c4YFTCQ2m5XSI0L0bXIX0jmqoaWjuIdsm/wpYhmqWVNY2KRGVO51nDbgcsiXVU06yvat0W
xZed9gXBUP493O3LKmMo6wG/ZB13QtPfmOjn59tWY8HEHTnSfKtNPvjtjXg4Lf0rdwlBkarH+e6+
CW+gIkLDE4NJoqQSyQOvqBoHn2nsCic2ZgfsYkQRYlFf4SM5KVBmz3WMbbgDNXlpMLdQ3RRSAwUL
WAVVx1dApGO2x7LWmMno2/67UBQJuQ0DZnys9ZtTsswX5rPaersTYoQ8r7G4aYRBCn59B6Y5lZWN
xN5uFNL9mr3oWQnm+DB6oELVAEBJA5ZuWtP1chuGmXAE6zhYXFNk8Tz7ZxkZIzvEsPlNPPKfuXVU
psjmCnRSUmfzjQeoQE3gwTHQDTc3dwLrz9JkoHD1/T65JUpKhRfmm8Y4ZubNfNBjKlioD2zD3TQq
b4kW1kBRnwyutJl2snaTFGXhmgsExfMA8EyEhUJfLaq6Z7r8GlRoRVUJ46tTQxOXtVxmkbR7ApOy
uZhhJsXiMCAtK9TWYo77Jj+zfJAGa0ZG/UsFn39VoC1Tg+H1Du6OI7xf0U3HJsO/Ov3GaddE65tz
axtG8trRuFQTvTlPBm4c/ngJqmUxb2yeWvuHWevOktMxlQVgq/fIQCjqkhPVLPvj6L9OxeocwMeo
kI+8+Vqyn0nHBBqJ4kol1+0hdSZPBt3LuwgjWB5j1HVAiB3hR1p0rjs/eO42C7MYTO7amEC/R9Ou
8T0L/vcmSMbA+R9VWLnD4wwgHbryzPMhGcvdFK2Rqgtj50OkmnOfuGxOQ5pkcx0cEt77rmJpaQf9
tRAeGKkjH7POYsF8XQAZ6WIE6PTzxBe0CbVpRQZnnCL1y39ze0kGJsziQS0Us/UNcMDxT53ERqS4
whF2hUm3DjJJY81j4beSIk1dMWmwkxUQ2nOixn9KEMdwN04DSyFqVfKTJPJh36WvuQJI0+0HxSyU
lSVqUvJKKTaOsZZQ542QoXKRBrOKD/Ov/9g0FSDP5zwIcfF2HvT7aJHeX/StyOkh7t3Vv2zbOTO2
DYtGk9x+pgXaZABI6+KII39QSkr3/0KOVdZSVQf5O7gaAawzZ3sU4LxnrVkC1SOJj24smf0qeQXs
Y/I6r2L6GkGNejQSDzXZqpMb9oz9+C7RwhJxU+3D2qJujWDypoJYaOfWp/GrO988Us3UQWyGgSf3
l/X2tPpcdCG1rncrpph5X1gCknXW2G0eodG3gu4qM7GFeSNFthSKA4lTG5EIcUBbp3TZX/NJjRgZ
Lm34Kdq/9qBQUpcer6yO6E5bghddIpz4aEKJTRANx3NA3+X5JPCHAGiYM6nf363fbo8QWnUTJUez
O7hiUNNOPpNsImIuG9Kl4hFdOXeo2LmYuvLKeEct7/OppnFsYRMM3H0CAriXwRdGn2XZUFq7IsZD
0n9zVxNtbnG929zkknZID5kRbsmMXQ0UyNWy4rdx0q7ehVK+6FGEdycpiJTW8CgFrr/7P0VkIxws
aV/5oHHoaoN3yQEEx260MD/gxqdaxza+kOSlxatUgurHLAcSE+kJnx8b4kZilFe3MuCzJz1un/mL
OVECm5hxOQder/fYPxtR+drRHbtrIuS3F/swusGsJRHrvE5Gz8Ye9AoJi6f+zCNKpzGaduJObGJi
zrGXAJrvg5Wp279fzeJVmuus5TJWEMCvjGmym4HoO/uIPj7m6lv8akr61qIeEnRCP5/z8fXviYYT
SRa3i0LKNJNgwkgwwjES34PBMY1KrVHVmeW1ff5dxYNnKs2haWIL60sU/kcQNeZ05PiZSwwhRiY0
NEGM+bka0/Zzi4Vl6GQymTiPZXxAHfqZG9H+Gq/NCxCxUMZ5WLto1Saup7Y4NlHlK5DiA3UkG8eI
wMqzUxHnXpmQUKOwfH/1qBe9QGLaxNRGUQTe2w8FS7/qr8XUm30wuUmcsp0Q/+PkAgmtyHqan+Zb
AHxJ2kgNi9B2yr1SRDAZqhqo9r7yDAC6bkPBeSMdFaEcI1+KKZDJga+g9MG26TAXgDGFg3idvx/4
3cb+8yYwjyDIbl8CByZ6WJ2PCyNgahPUL9Ho/VdZXL4Re0ZSvteJ1oilLvL2Nw0HC2BLSS+hBXhY
QxBEduH6vJgtgTcvlY6gVaH8xa0ZQPseQ1wbEdkc+bHdJET1lM8miuynVww2z170Xjek00TYFc2F
xMytDFYvhHVn+ScXM4v+WudaEU2Kfp1Pck10sw9jalo9SNXagFF+HeMc2Z0XHvn2Rl3WfYr24cDq
6rflO7dsdmNaoTusvmR38lDpBN4i1j9fGa+/JOxrbqWONklrNTvaEdn0ZuZ3O53vEA5AnSjKxvTT
EJsNdxX7rZ/LOIDgPLKdlS75ds5YwQ76GEKuWyozS178NOkxTQwA8bldwTVELV7xEqGMTaaLBpj4
s8Sp5LtuZRZrEpLJy4OQfd1TsQ9mHgytbtM5moDuD3Q2Jb/XYAH/5DtCb36otRMseRQ+D0QV2vfW
rWXhJIC2n1N5luO5YsMAvhMi0DCVTJQvg7skJx19sYJk1MxTD+ga0jkck8GOh68pjb6HK2DLgX+R
FviYljVtbu4untmQ70tjCY4IXSydfpKpRIoAGawp0g/CBjDeXkp1n+kYR2Guc/BsIghTZOJ1AcJH
mHB2FfepbQThZSVlVm2EDBoLr+t11HNThp/M1xZ9KKs+fbhI57rbYhC8AFt3ZqS6WLDr/Sd8n+Q0
X4PpSzxeQKLaSws/IwGDnIJCO/8NAoQTXEgXvzYmUnIabbzvjhcqEhUrEJ5jVF2RzADyliKuDe6z
vLC2dayUvj/BsGeZTYl3+Q2AwR74nNtukUCUYFF9n9MpwgW0EGP3oqFISiqxo3nTyrvxVuilUJ+M
HdKZfHqKIB/mEoPdk8UqSv6hKxlJFP6U0ROm4do6ItP+d3yEqLi6YMTPFKZXAMFG9KmmqzbvLwQe
Ri5H8/yxkyflFbqDzwRUCz4KI++wcG6D0PI9zrHkMVLmm/EGbLh4FTJfysYSv9QtOOyIq28T+aYx
2jqoC74qBuMyiaxi9mFoIc1ehKPVwDhzWcSsXTlrU4AIGMoK0K3EMQeF9DcONRF8AlnQrxRgkJr7
Fm636vjiAlva3oNFJg6cwCkVUuTP/wNGlqAcM/IW06l16BiuPhgURV4zG4vHf4xrFmtJu7Pe/T++
gVuLChYTWSUFn03GHt7FxsjHURpiYsHcISnsywfO1LwC9PtMBYVhmhvUENU6SjitK1mtS+qurIFj
Ov/YipmVr1Nueha6NsWmwsT5q0e+u7JwX+Ms6dDNxSZ1HeKwS7ICXQuxTfxtZDXxztnwGlQBDI7T
sG9ILKkgt9bxd6KUml7vquQ0meGTZicvEfyqAA+cAcnhWrlkz41BK7kMd3hoc1QhFSxtVPXiE20C
9PECf6Dxzw9+WKTmnhyqDDH6xmvtVii2k925o0YmK7Ijfc3UaoaICd7YVDEPemPeTJxHjVL5ZW2L
y9YwYuMTTlFIqgqoxRHDaN0Xu6+hRBg6n8j+6S+687kMEI7RUm/mNaD1rU8QgboTpfP/MMA2lgK1
YMXdCWYkwkulNa7I2LFIoOSlyjASaENcg16GaxEAV2KMartdw2Fuj5cT4dKNUlqA0/NxM+MWl2J0
cqgA3/eO33+3eu4EnJ6BVdFibxcevM1u7C7FUSrDG6XteGFyhyqUKNiKU9I5EiAGb/O5sWt3V9I6
5e1m++rK6uJbMsbIIlpyVpV3AUys+WpdnjB7dsVMhSYWpS3NyenanuiEKAOaJSGP4W7thyIp7JV3
arm+PsMTY1SKmdeqEDxzxsR1zAgR7++YDIxWPXBxsqopaNjCYEg5FtCqzrDz5FgrvKTMdxpzl90x
VRIPpbD9yw1xJEuPQwiWQ1ZLvyk6SHsKUuNJExF0mu2V1Vqjqpt676X8TaILb9PeJhjRHO2Ofst0
ULh9GcazOuaHPgxN2KkDVdAkvIamODiz0EoxFwNZyfd6KCDoraKvo8SBGGmP1o1lJa7yjNK/Nkm2
nFLt+eUwqwDcIiOh5H3g3HKZIsFbP/HjfNsSeFiDmpdM4zwSlv8fXpCMQ/wdsksu0eX/Pja+K5Oj
m/irzNI91cOj+i6LLHvtxFrOGd7ZoEuAxv5593vW5yKyzkeDYIgTcgI83ZLqfTy99CndRDaojA2y
Qw2wh+rZmvzzLVshUSG5S0mFJQ46CDexMlfMbyx6aOQRlPitRj2d8735QJ0wX5nmd8rpWjf2tIz2
0JgOOdvnJtZ+VVc875eaD9xw3i63Jqvzt3OTeKsovMjus6U6Zv9MXeuo/5oJGXc3zLto2/ERqtps
ZRY0/r5UNbcOJ2uEK2Eu47qD/9n6uzEv5RBqKeptCRkZz1gldF6Q+xsge80ZTGa5MqOY2cnrNAtq
W8eSaNlFDL+omwguwJhvbQ+w5c+uXP5VUwGb81w+AjLCI60651TBzvG77UJZaFzdV3IqyqmJF65I
jnOU0rIrnbtK0bsStAxSorZ29kgjoIFzEheYtqSb1FZpAT3oEW4xPfs+b5MIwM20nKFugdUP7IC/
hm/kdXClIM5AAo7g8GTIHVQ8Y8TlXX64vf56ZkR+2RmhXLjyi0cnaL9jgF28vzuOrRGe4op0oZdF
MEAg/z5oovPd+/RsLuEYvMutfCAYtzNiBI5f3lsQ0hfRiDSA8fX/Ez+hKd9ZiCXNpbknrIFPSI8h
XvlwdgWTwnM0gs/lc0BbmPEEflvzcQQyEC2CUmHIEatHIPBS2XOE1ooQmjldA7OiIClXtEofuQ3Q
60rJIxHLF3latKNK27SUuNBH6gtVR+Rdzw8KV7qSqmTCkNgRqrw/Nket22aAscbYjOmhTzmoMvvS
yEQiQLqflRUC9JF0NvJXM0AiV7+yS94XFdC/MeDnCO+CrzM6ttiJVaPNTzaRQwvd6th+CwzL2VvH
S093AwdLfCHm5hXv/wQjhv5CJ/qCyV8nwYalVaI62LAvUFO3hekCQM7T2bqUyOj2Xf4tsVZpjpBc
ODNqa7QI45ePGpEpv2kCvBEeQ7re9aQQm6uTMqId3Xn7SgD4Qm7xDtjk39+ZMH9FTC1XPhfILLCk
WRzQ9M9w+dWgUHixAmwiYG984F85pn1j/3gc3By6blMJntpLVDukkMpzZTP7ytFA16IVnJS5uwsP
FEUFGRvsNiQeneqyQKkdCij8Aw9XNuMtQCNtz1fsvQ7uH1O1NG9gm2fXnPf42Ow2vTuxFe4jls/e
Wwvammmq8DQ47pKYjgCy90r5b4M9HkR+DJ1TSi1/ioeqwgNEza+ofIDu2tF5bOWPyWIf90j5pKsa
AUfCCXaQ+kOech3mcBPC6v8+r8HyOxvYD3A48wLB1TsSHhOCclQFBsoKjBqsisjpr8Jg8bsM7/Fd
EGdnI7Y80pvWY030lFbVlAwecjVXNKVfaDEHSOq+MSANbQZ2Y7zDfk1joZBIk0aGDp21J86rNsuP
eR67rYXIKuJmgJ5x7eiR4Lw3SP3knGSg/wqdvOhgSxOtU3BoiQkqY2gg6wRPUYB+B/bCxiMH5UV9
an+FKuyjL6P9cxT+zP8BCEnm5YaXUJS+WO7gb3S+9/XyyQxOL2k/mHRxIPJTOjpKtu0u/DQtwEBt
Hs4LuJBqaJfn95tI1krBGTkpLJGFWgIfgD8CERvSRmpPf9x53AnaHuftUg5fawN/BzdsG1P3ty/V
2ksDpreWcjPIuKl9V0Nld9puADTr7PrnCu+cBij9TW5L6ryOohV7SuehIW8ywhWmGK03FLkvyrFl
uyNPuXkJrPkrV+rBe8gOW0unTFs8q4bcyoF/20oUx8/dDTQOCMeCKXuYGMmBIME2y7ThggSSTD6g
0y9nxrK0DbniUFsr46uzfVgLc2xML0zXOSHnBh8m+Kh8b5vM7AXSOzVd5HAcI5eI2aXLJq+JgYIQ
crCUquOEX/XWkbX/WjDa6kwjPydBqqCSARiTK0ndh00TSK6P5iMzPgIGOafii/hgRifPt4/NwYVC
Asl9Kdlq5ZClntgUcUpdD/RIDhxTsEhHHAHomx6tltVz4SLsYK5sMKLdDhebvpgJ2FRJi/i9i+n0
lUYtKgNAka/VG065jj0J9g5CbYzoB8e+Wj4CYU0ChxG4jNiYYEVuZGWm4dkz+bNZZMCDIEdc+Qub
4UqN9L2IQJ1BbIqvIFxGTGTB3rTFPUWuO5rmPK4JilhERMgPEG8yWPLl+ZU4xYQixDcfaku1jdgO
dNfBGx7aYgFuNxmc5dHfU4bgFjrF9c+CCVJ1DOSiF/eE+71zC1G+UpsDeattij/u30cHhAI1lhjO
NEfLXh9mbWgCyRP92+58NJGl4DG2UZEjZQ6QFRFc53hqhXEN8g+v9tc2mTv82U2ft0kKYWJvO6tK
tQTv/G3/iGlQxV6N/sEMAA6GPtmvBgy/DqA7BakEzK2h2SQIzpc+m8QGBrfFdAuhtvxntAs3eovo
UAMw7Y8JMsNn1UPQVIeU4cVNGCEEAUavkE4XXteSX22LpOg3bSs9xMLf4HC4/XomtKxp5ehksAhn
weK74JsMLfgWamGBLaM/3J9SvHEnG0gDy9oNYUY03Lw/F1PR22kZpbMHNb3EMmHQhJx0XaR53jVC
1+V1wpREfszh9GC4ABQxk7crmC4EjNqzbThhe7IJSOzJs2KwkvYtLcg8uub+swjhfC1h4EtJ/I4V
q86qwh393pY19vb1dFqfUAAUa4UWoivBOmEkn2IKmUI46VW6oMl+C7leyO+bneG5m7TlEa2veSC5
ujcb3rWNiyOxSc2Mu8BplQtxu5B9V/h2krHivlsMSrDSTR7rwNs3uaYvL2zJR6tIUX14ywshx6wb
cLpvaINPQRCXoSaRNuRYa0O810y7ngGJD7dnrKC30EzMAWLHMJRaJyvzeJjUsHmTO/MEVzHmDPuo
k2tzkAjRiBLZ3W94JajHKeIHhR0KmLpNn9+/kEb6GBdCVBhDg3kmzrA6IZQv4c5FJEsXOuyurFEv
JUIX2zvBXkrVrF3EjZ60w3yEu2OzsqDOwZ8ILtXKT0IflwHOxBgYs4IK3jthSN4RGozCvnI6WUPY
rQSzARvCHfvvzjtP5L6t5IODpm7WVMFEQMkhMxGoux6J3JOOQfu0n0bODreeIkVeuP5L56Wq0P1G
oNPgl4IMoc/XJk3PgMkfzeCCKKyNtXu6ZH/wL744TDCUNldF4qh83lO1mP5tFzms4qV0CdiIDqlS
UwE1+dRN5F9RIcUx4sfFo1c/tEL8P9pFxYdPREhW8qigFekMyGTiVDjnLasw5aflTfzVxq5nSfB+
39SrswrBgCvMLuUQWOsywXFN3tEm0jQYu48GMwxXzdVkIF3lMbcEpZsNYsykq8rwIoKlsfv0P6Bg
R3a+VtLT1kyK9iU65iRZ8coZLHItu/l7NOXSf5r7VeIKTCwOKxtQaQhdpsolmuyIFrfZF8jjrLEm
i1NG1tmTBfVphsMEPeE+WNHiXxdqdTiFrMEFodAokQNZYi//lkH0TpJClhTqpbuJOTpDjcoqz3Hr
wjY3apfdtbz861Qba7Jhap8Nkm+j1WU51P4KxTxZ4npSeSYPBmhOBRgoWj4CP+ZRMjA4NieuQ/7K
q/Ab3/4rmw6a2k0jebkTjR68QxfTmjej6jl6NdiAG0bAona6mc8IsHqkMh4vh76zPbYIGtnNPFpX
KPlXmxPMyHBrw1WVt+vtYlkEsA4CTA686Hccv+cJEeO1BprCbzPxDTfVyrSy3Let6Npq9H8i4mKS
RfJHiz8MVDMCz4CrehUm0ySZQo3iJVCRuzu7GuMZzKHr2C4iUb4Vef0oGxRXIxwpPTd0IssWWSCX
JGs9G/YUph4ieuUD4DNqQDZztQ6y7KwVuDtf76vLNS0cUV4rwRzgU1yyhXjcX6UhRpS+iL2uJinE
rvuLNWJqujupuVpWzLqwE6pIrliHLMEPOL2iMNaF5Tp5NLI/1Gc+YR9d7UC5fegDcqxRzYLYhDuy
L6pwYrCuj8UUjbl3NAJXTRcANwzo/FDyOQf7OPoKaayVcHVv9stvcFnIQbdjNlXCD69GsQszTz85
XHAP4qaoqxt5UxWoYG1TBI5zx90zyiSIbgcYXe6SPBEHgafR/IKSZh/ZbmxU7kBPRddf85RwdjfV
R548pP+l/Jb0HXtnPnePIzS8UGPkPo0BHY+rPUqLWKip2EN4HlQucV5+Eoe9R3WG8ew2Y/U7tzl/
4jwirth90s6/dJ+K9H30L4NFRJlTuYRtms2nckDJj4lSkhsp2AGalfejctBoKEGe/igJTrmebGir
H3QQNiY0tolkrUUu8/bvcPqkSgBMTiPZa/fkOV0TbIC1UYpq0W9oOWr1CtTA4abPeqvejTXoRi3I
0VxX9m9FZqkEnGbLb4wChcBJ/LsWRWMwI8QyuXKaAOoGBDnM2ZDBC0QDGb5q87qpdyPUPoKzKYPV
YCvb4rQCc4eTagj6eO3m+UxZIymgf8TkLdGHEKT5LOq0iqNUG0wt04WkdAk4TX2WBkEjz1M8cNI+
AneXuM0vvCvH8hCcM9yriYcnRiw+AIWWgqqt8Y4t14u+QV1dFfWi6NzKsXB2WHNI8lzLhGZNCCb2
rNhjZc29yh4QlmPudS/yB6BOtOgWJFVk6sRuxJmQ78+vegrHp1QHIDxT35NySSRVYpx63W32ie/Q
zCXFvY+84konfSzg/boZBE/JwQQ1aztyhNKSJteMF/rBOoBA7SVMU6BDQTxarcilNppFPTWRjiaO
n3yt1V8MgoqyVXNfLMaU3Z3/zCIzDvyHlt6fRjS+kyMbr9A7egJY/mMdYauZ/MEFj3+x8AnG76dm
76BYFFQb/GyJQUNPYMIcY7+R3FhaMh6pSzvBrnhzRyI8vd8Bw8KSYmtjX6fb0oyhoJpxhcndH3oI
x5vrGQooxqcuFtCvbaJQI/W1skufw7n4BKQIYFaTz5oomh6OFYFXMQO6fxulGu88WPT3p++dvuiL
ChbhaWk5S0rHuzQ0V9lj4kJhZNGpwXS4HbkQwwTbgj/94dZhAO1dNOgxwJ6VxajFuwwuZLS64jxT
54aJ+IURGkUgj7pDkwjWDJKAz9SXn8eqO/0O2AO1Awh//ZAPXb+PpqA0EsgInjoimkaJJAuC1SeZ
lbFwHuQsmV2x2JFi21OaMwLaGZXPeT2+A9gp0LZR+KwCj06ALRjvmB7BDeLA2PcLHhuhsH0/5mw5
78rh43K0lD0NLBDRBxh2QEV1vu/Uje5p1hjX7pL6EZ0Y+s4gqQYJRizBmUlHsgLm9aXwwIL+xg9m
vyxi4s6snW+vBGGtl+voQckRoIm4nqiHpI1vL4CdE4AkTzMV9zLUTFiZWe0qlVLlKEH7U+0ivs+D
SoIYp+RjYRzQnGnOw8ou23mK4ugLzL7mlkTGg06Py/TRXz3NHZrO2AOlsBGWlQdiJDDfSylorMd1
J+WBXx+7bLk07DOztrd7qJrg8o+R3VtL4ZdJKU7ynJQOcB03Fdfjldd737JswxCqi/eRrfDlpewf
dgInsA7hr+cLOuX9U/U2erKj60y93TEf6hlbQI7UmMxEk4GnNSPbX+/pkXujxLttM6+KeV9tJc3J
kZAqwWGtQcDOmvIcAvuAR0ENtRiBJiaEbdg7hknoKm/LewZtrGYiLPmBHnXPHhwGMdzBM0CsQ1UU
V19yNZprsjQiMYqvkX64JbnOKEb6fL4T1gWlsVuhnwoptWoM9h45pd8yRnp9SYrtZCDyzvRRo51+
otLqUrV8jdj2pakzoD1wkDGyEtwt33zoOhyYmkpvTOiO3aZ4hMDz25Vg5kmJb8zVBKYS8tlluzUq
cid28P1J9mGmSxFL7IltbvSku/SFD8Z2axiPXH9jyCrr//EukTrfmL+CV8HwC2CkOtM2Onky76P1
JAdLvm9nbqnHtNuHr2lvbLxpBWeBNZTnhL1vX3/Ltwp/DRt+a4tC5zN43gb28VJY7HEuPNnbdzbb
jpQhPOSZu/PjNMQftTlwGlXk7hrVYcgeMfbjMWthxU4ehHmUg+14dPh5FQVKgxBUXTSxKZjbfYlY
RKvSDPZY7D0slhCsD/jIL+f/JuhGzu9D9oFsv0t39EKslEfJ1ENtpERV18joY0T+nvxEqnyvFdgD
pPytv/uyxpA78n3c9B227Eo6akB4K6S219MPSnpnviYBT7uh1IWio5QxlTzkNX25+toHl+RSWulg
CGCCvY40pjodfHLkZZxtKwn8MQiTL7+lHEc9suCXSQTcTPftfIjTGWjwHO40aXiZ6XE3su2dNUXC
ybyTJb3gvucO8jSDkRL2Qi6H8qoLvs/6a8mV397hrN+QX0jzjgg3XHNDKIc4BwXW/HgUvOKSWxC4
qE/A1Jf265wRwJNbUjPutiCWO93BGCsJ7w+Iu4cMPMc2bQHvvOMRIUgAIedPM6r5ki4casYgZ8rJ
29sedo7tRLKZsSSDGZKxFa5KsM1MyuOkP8Jqm5tBCHm/FmJtypwxI2n/AuocRg0mWYhVS88iM7pZ
IY9u/KXgObhQZ3Fwdl0zqup/FUpDw+Z47ON2WVShyuZOfuEYF4Hzf1obSyidYfBgeaerBOoJwt2/
E7YWPktpQW6OGADyf4slJ6AGG7F9LBdGW63HH/k7YEv3cOBZ6nsEz3KiY9gxfUD1xGnyFcJUMmqQ
rDiwJVS5GuVnUvZLyObAUIiPSE0dqiqVOuSUOJ+k5GQCkDjAC7gPDyU/pkm2WOpltBlMnwOgmyS/
kxJLj8B12qwFx0ad3Wb9CchRv3m4ywR8/FD5iDc4fCPF/FfVDR1tsBdaIkjr3X2pYXJj6aWedX1h
S/LMU1Z/37GvdPPAnMwodG8RaArvOU6BlYJSjWZuoLcy4txPQKbJ7kKmByAWZstcqjViszNjYAJ2
4PY46+LgmgORzLSt87C6HsJF28E+KNClEiWHovtLUhldjZG+s19UBg9/MosQPK8tYWdbuQiouzEE
WlObMVH+2WI62HPiTaZQmWaTlaxVv6aEYzwGZrPHsv6paG7tuN1IwgGJP6lYs20mdwMIvlf5njNA
oM2CS2PXIzUz3ntxL95USqucE14xKvOQoS3YqZ5uQK+2MQdcYAsnR/unDErURmtCWfyECY11tdyH
6d0hXp5VICUUTa2FgtnHFg6+2/wBuGnNkZPv6ZE3Hi1XtgmlevCZ9pRnTZDDYV97oxZgB+BPAtBg
vtil1kIYH0bsMTcNak5mUIRgCtMDQaHywiPVdjPoI8EugOjM+Po/KfjI12abnylwZ6I3ZYiht+hJ
9JKUpo+ikXox5BPVt74jtyGNAu6clNhg+k/nRej5nYL7cFqEDFxOM+4woK6ftCdcvhghWJV5p4IS
QLtd/Xr2hVMJJKjHchGJ5G0XzxLiJ2HeZxaFKhf6GonimrpTlpM7H+jiYHZE4FggOlW3GLng2Iit
5XwOJJKlc2uZrRl6QYWx9h4Fkox1vrFDC4abzJYosngA8tJcGshAGy6rqnxvhW9MEVVSYH4BhuXy
WkFCNivvD2ZTm50pXf/1wbjq6dl2uiQFBntUSng6tw98x8nRJNFudlBbgvMhEzAc3yzXD4iNe12j
x0T13js6DLZDWrrlMcqZHXqwAzHkuDZlgX3Pp6NcGa7fNcf1ZN/vcMQN4AsC5A2Pg+s331f/3JnG
UIwC9bmFn5JTgWp9aNHxof/1nZBj/8i/ykL6f9CQquDWm/hFudgpfOhg5r847s1tDiNh0BRUheUQ
D5hkhQOp3udbPyT56GXObWTKeBkL7wLaJ08ffk+SS4i//DxfSzScZ4zk6QHSvnewrFj8Ng2l4H6q
WAs7D4f6Hs1+7zMfmtcT5eM/mkYmAiCFxq8Q2AXTuQ/2wVrtZeSClBtWaw+wjZw1T1Sn9SDt2i+5
IakgDw+QWZU9UvXxkORZdOebSi6c4OSY7exxNeqMLrpeP9EAFnz03z8uPshnToFTyFcovcnKdtn7
43luzkBtkCj2GSpNtivZueso5t9OCo8gD9iJmWQOkAXm1VifB8en5H93YVDRUk/Mh6m4WcU3+9vZ
LCLc9fBT4bgWkKqY7FqcBgFbsCewKAlvfCbkNEnhIGO7m0LbfQ42D4MMdsjOwdyGxrDaPtDDu/go
Yeu/9IQUQ46iYzih1KRqNMNbEA/KrtQTYZyHr7ZzpwBXqOH/+GGr8jmB55gKgoNw2wVIoZk9rYKE
GuXBzardYNhx6BxkZtHYPKYkcSjmXXF8peQ9WoW/B0GE9rNkjGNUqhCgko1XvQ50pVNCjwJDIhdI
ulyu1xWfqI4Q713FtzAFhnaE9ZPVZKHNVW7L/T7Lq1B9t8J8QqSfO/bILXZ4fTnZhKxe0/cSfWIA
Ilf7cf1SydT2foz8jbTNVkLaBz3iZCVADVBDWdaoyFTdH92HyFq3rLethmubkwhKnjP/xC3EZVc/
gWs8VsX8mS6HH05hR+nmmC+ozbH7LAzGHwAOUzwiHLbu097irQLPd2v0GvfvmGNQHSNP3SNuBmo1
FCsFXzufvXldBnrXpaAikwSn8uWnYH2YLYUtEGfnCDfJM/4zXtxFH9rj3e+BJCW7ZzCzA5gwDWC7
0DQOvdFHEaJrjQutzBENkqMRoMDhvrgd8H94JkuwZkR1kPxLY2kns6SP6scQgC2c/fuj8wPElcah
FPbuIvZJnU2HonxJxlRksXcY1L45rDbfAO4NlImfxf5pSuUUvA7RJPGl1e26/GuNqIe9lw6Oh9Sq
Vi+OaEui/XCjqCOuR6IE0e03xKnrTGywhtAKzdrcXyiA6CM3DGdcWr0BNKeN0yv+ZFWVPgTbhgls
OadsVnxluRpDsk9SvaH3KQ+8zwXGi9jzBUJfvVNLCqtVqUGUZ68OXNj/IEN9fy3ftQXvQnsPPYWe
evcR5spI7wk+hBSwWqhRMyg7LJoHIiwvJmieocBrmZr1lk6Id9KzoyX8h+4KoIYaDxM8Z41TtsRS
y7hengxUasVJLtRwJc3YBDb/QDeA78YLzS6B0zYjPwkhXLX1WceOfKmaMfPhKwpMLGgYaXJTdsct
FAWwvMQMQlRagHHLbkP7/RVuHvi3S/EJcSPsLwonPOj9kdY5twSaER/MGyD64cVK4Hpegmp3vB9E
NPAg+4X5NLXpuKyqZttw6kp93W1qfh43Eza2ZEXhvPCubiEYjYaW0M6B2BcN1RmsJAsvyLBXM+5a
X1M+4H4dNPvRNQNICk2GAavyPhloC1jrbG+uSvZkxU602nIA1/7t2THTTBlhHkFI1glaoMNBbbpI
qGHtZ4ky3gXIrGT/b80ajfkBwrNLFRHidznQELz8lttobEuKTvMxB7p/OXHmVqWURHvYxbHlEFda
KoLUUbz0s2WP6NSufUusKv0UDOywBGdpc1zl7LUUUM4aFOumpVZFbIn1HBIOayBgBDhgPBRwahAz
8D5qJ0hZQaOsihNCsOYXX6dD1IEqqkA710q/VHlX0FoaOjK6SrEcrITIiPPvAe8fe4eMMFPxykIH
pTxVe2jei06TaQyYizWAGiSUS5jCy7CSyHoqbIZwMXtj2P1f/HL0W1xlO0YCrQ2+jLncYlM18M6w
IdhV/XeYFW6KfVKzIaFtzjvAaeTYS+GroBl/2L19Jk4+kZMpgfWcuZixsy96y+AVkxoi0I9tbWVE
amXnkT2Deh/YPwCl12F7c9zYFzz3lAO3SjnzD7lksU6c9TzjuP8mXuD2Vm+0Hf4r4svQ7rT/FK/K
3F1AITgzzhzzulNWvfrQS6yH+dK6oxBzOkJ4bthKab4Y1zSyFNmQChFmq3TfhcoHYoWJlmyZHI+W
NWi2CfXSrndo3jUG/kvg3a8p/dIblUKPfqms4VI+awgKjgUBXhng4t68XU6rrf0C6M9sBrZVYsVz
1A0+Tw4e6gq0MLMAvkHFaPZjB/1yxZNc7RblSkpJdWNPECZBsgA0MLVAjIwcaaJ0Hy62IvFC3pws
qVNTR8Jmw4t6gu/3F5QttyDF3z4hA/V/FeQ4WGq/1ASn+XcTI9a5ltdRCDyic0Lkverj/Vs22PK6
sKYL9RuiFkcHJQVGD0Pc8+Xi/RNPi40Lw9pBVI5l6z9YmeZoo6Kuk6Qfgq0yCKqvMcvREJ5Te4zF
wI+ON+oMnj5c3fJc3NqPxEribtkv6/hmHWegZTXm5aiSncT9Fj2f3NyNSbJGexLVuBJfn23kzunv
AvzVM8qAIJv70ca+SwiJy3sFC/kdF7LWBIoKTEWf7ZO3IT/aMPdDxUNCDSeuQgBMJF1lznS9/Km6
tafJKmIuzCKL7zPxHZvRzJNIk1PQq7AtnkMzxHhhWLc6wRwCEHAu3XViXfY16TJLnxsPJV6myq0X
MqbKcJ4C0h5uBB6lqwooNfaJsWurdMT63vyyFTrk91putGuqbB5Y1Ht4XmydYYAbqRrRmFlAZxsZ
oLMnru/fAChASZtApatdScp5CFJnX4Hd+RFW+6FSyYAuTGNBeSKp1RCUqKL+yZfYH4H3xW0ZPVdF
Q7bYPncGrG0yVL33Q9CfXzWDqzkYmrgAq35U45a9dan06eJPT0st+QDsThMqRfMmeKpbPzoqWV44
H3p8GKkbU+Al5U3Wbkp2OgCK8RvtQvjmPrfdl3wkl0B9D8Idb5lwdXmrXqgDirJjdsOvmpv2p1JP
LHZrituLyLkllMfH+ozSmedq+zL4vkd58+BwGn1Ullzy4YbLmgQcc9gb9KTvBYAvLCh6wjsBSo4j
yvTCuCH+9YkvkjitYCRz+c1dXOJPM1G0/IXqYRMDF3VaUzFKfvM/GfxNiuAk/J+gy8COQNNVzn4a
pkFkqedzvyi+ClS/vl0J1ieRHh/MMy4NWs2ouOBfLHS5QkNUHHd1l3QUVFQGFhRdkiTFgpKh/E7Z
pQ0KY91UrwTXXQx8lWgMFZl5TpUkJ93jzIqkCAxEKDi9DLWrU9yXYXBfmPZEARDpzk6X40tZOIFB
lNcva3AeSwnup3FJukVWZNKZGwzYJ8Suy3yqIeDVTHNyGW5WpUHbrH+PYNCEcvBjos23qBeoH6im
WEGb7L7p4kDNquOqMHlDbCrultwGh1HEiKUt9eA50DSq+dMWrTx1Q7Ee92zB3CcmFTUkonD3rwW+
X8d1ML4BqGZ+Bb+Kg+byKvewGrCkx4Jhf03sw4Q7tFF8oKfC8c6WJT9yaAST7C0hzmB7278zJXkc
28bt8sfkwshCOF3vJxdeDF96MjcTAg5e9T4/b3/1wkovmuoCnO2EfN7KSzv05dKDYo5EHn7GTVd0
M56dmrF35Eqo1AUaTw0iDr90QQU6mkxmQIjaKM0bEXgBaYqJiX+7pDAiSopRL6f8SiN1TLZbucFH
E81V3kRXpPA+BpU3C8KQLXjeq+P+TEsk3aBbyz01VOBNptYCiGCzLGXlnSZmimqJelGAJnpw5DQ3
1OL4fALPPKuZeA1wBEXxcWpnm2kdhviiJrY6jk8cbqxd74BBl8K4FiZta15E7cgG4LZksJgMb2lG
F3jycbrFHq91swD0nnoZuYnkuupfuh286ItjiRlt1GWJ8T69i08kbJXfjb12VFrMFikJnRBvUc5l
lyrfdjfQN2wAE6WaJmOuSsk1yX1XYLEGu5PQwoFWvCUyFXeMfob8rl4PQ5WC08aJ2cNR6xz9zoVF
oCC+AT4+oGM9TYTelvhD4AWSLVDaBZHtKiGegCv24gtnCMIeSQNFugRtgVnggnyPN4y5irgIcoVT
2RAXv/yJY97pduPmq5YF3kFHQPjdbZ4ERFpR/w0AgqJIGD1uB1gkWO6z+i4x83f8T5A0tfqSwnTC
2nCLOScHHop5SfVdLFJ0u+2RLZYdD1YuguMXBP/m7KwhrkEOeglXwAGEDpogBVCgDOAILZX3Nm/B
PzmrFBy2XGhB/i6mcEFyp37iOiXAUOwn6tbXC5FbsgjS9fbjvjfQojEyL3LaikGsly5J7FZAuIsp
Mr+6X/0ohklJBwyv78wMvJGdcJ0CX3DF9j8cJkQui4E2cVhJ1wvEBGtHeZGmMYjEIVzFL6xT/no9
qE27bXOhxgt/ls1vSNr8dghK/ArC9jMGg1weMhoH4AP6S3VsIlaAjPy72XdZM1jpeF8z+VVIwDJy
lgtC4ignP26sU0bmvImBqcvx8TRDfU+3hhx9q8om7faCKVJHQiY/6+TsxFV3UTXakOkWyw6t3wze
fKAia06kOcWvtWVQZrszIjS7US34YCUvagHBvKmUzQ8D47oiujP7HjcVGcIcGS0T910/M0pvSSAq
nqfRNXRzj1lPhOeQJpm6lyaTcCz6Lqba0rxxjaoTX3Jas4/VS7sklcUAAM1GdAcTiIGpxGDl9o69
iiKUN7TdWtEti0Tn42AVaxl+HR3v7q021Ep0S5CIgBaSUz0qbpWBf19tJhC1cihS39kPAe90dmmS
5aTlFXTdO7b9qjSNboRjraSDfAAy42EYN/AyHjAxm+THz2UJygnFerKk5sdKD/CuN1F8KKhPeS8M
gmBwh+qjKmvcfaNUDOtTlrPkDiQEhSLpjzJpCfpc6mZDHdkK5LdjoAV8mXu3+rVoPBZu6E37WkjD
e0pNJB3HfEP5vwqs8ic4X2KohOKIRqWko7a3hczkvKpZJ9h91Gam9uW39+DuyHa01ZWh7hEIWJvA
nZBX9gQ4325FcAtlXOyDm0RB0INFG6mHihyuLafab1Uc8mTz9mR2aUKZSYDtZfd5z9bZN+CTjqzh
yLG6vpdhxajEz0upfA1fe+03sowawdYzp2+ZyNuj/jsZ4YqsVwuEzHcY16TAOC2G0Wq4tKDGrPpL
dpoANL+oHmg4ka1n4kjxt+xIptNKB5YHRM1cVJW1XdoHyXHxpgHy2v5pM0nfBEB6FsDey9cUBI4G
rJ5GbZBMuU0HcHpZAAC6Vg3uUkXNjVA6ur6fto5Yf1F0m1Pwq2WbyeXsre9RPQOruoKzJgoyMUKI
wsODJrzvD4Wxd3j8r90J+GNkDx/nR6TKex7Oli9VRy6Fb9aXPiy7d5RmWfEqVMllPcaw6MUcElCz
pPz4E94MwcGcTgi0/vQnOXwwofYZTbK+YYPyqZcsXwCa0a0HP4BEh8Qd1dEWw8Hdbn4uATuX4/Jl
x+VJPMJK4Ybp925pr9A7owZcYECPko0vNyrml7LXHV7Mu1E3u5ROOkKREz/zeIqxW0aG6Z9iqNlv
Ja0JK8iIKf/tfTbpvZVVkrpXylv/QAwlr8dVZSMKIVH1wqvk3uvFXcIkZUqg47vr5uAm/+ajYfSm
SRXMoQ0l/eXZmLR6cIaGXHczbDlINFllaqDOSyqRW+mxPDWglR8UKJ2b/sFZCZtEYszluHKsMivQ
o2gQ0/DFJLwEpnMGMm9bSp83kN12Me1Vb7IfHGkJkRgCu92FksoKfG81j1yXd5NxzBFREX6Px2XB
cxFBEVRrDI5Hto6n2LCV0kihMQWB8RpsA+X8bMejecHctnW+xG4jOzqRMpDXA40qzMAW2QNQUsgW
0sorX+foKDrMZoO+qSWz5qfYC9Kakz7Q+EUq6SMD7Nxxuihuu13BldrPdOxHBJNK/zpORyvMjUfW
5iT2uzWk6uCTHgGonSd7oADANtf2o/GBRCUxZL6/x2rU8bFHz2xU5cmrSJasDnNPjr9iqXW3sUta
twb08xGVNiWqDKueicp2/0qYTouQppnW6nu5fAdjHBzT2W+3qQWGMjBUV+az6GEtWfR0lS8u7Voh
A6qCHPWDgcFVg5juIXOILDmhZL01g2N0rZXgbkBcd3iyAlKrjDJaEIHh/B6Gsk+q4klRoNH1wxGz
ShoW8YI83BNwWteV2snqby7raXyFSVA8fJXsWjj3g8NNxr7Y2PTHdd+rUuxuP71hO4c2gu30Dj/t
3LME+X84TxTt4rKhEMRkIEof9JTLcUTd7ZmNWjLh7t51Yq0+WrBLFKLnPq8IPpc4IY8b2xCxra7x
J5a14/W/3kxJ7V0ta5Irjtg4DM8QQrF4iJI5S523KSua3uO6nxqC3o75WfWMLLLKNyZkuY3Xp5b9
tlh8NqHwBDP1Ldo15tCAaKS6Yjami/BjEbbskOKtCFp+ZDGJdRAYUtuDZ/ruS8u7JyoKhN85eG67
yhJ4Osx+xnNzLItJHluom0zhgh8wHd/lpArJABzVlnQLqeoY05npJ+iHZCGayoHNve5c5xkHOZnR
Vk7J8JtNgVZyxZwTjy/OU4UDfatyo2yUW3uJe4bRxq/32DVMvvjM8DgDZgw50deM2XSdb2MbP2nb
c8NxgLw7xBOHw8JkizKktbJNIGO98WhRUpfa1O8x+RzpZC/utOYmcwTZvOfU/JED2uKSZxSR1Ejx
6pJXL07LICQIHt897htdwRYq/wa+V9QF3iIWdhEg/nQoqIJNLDbeDEK1VXHuD5x49r81O3xBCrx0
bzdGpaXuwXU0ewyJwt2wuPt1HuxZH2I9hwQmpx/ivit1C4NKBNYqn08vhOjXDx4a8I16cydVYncz
l3HHY2bufyASO/SmvcvGWMKU1QWU+uKr4oxYjbceuAm3Ex4pjoVM/uqu8Wo9y9h+chqDw3EaIRu5
fCFPN/pZwtEMcCthV7g7rMhmA2b1SdfPouNjl528FrOawH1wY++UdtcBZt7b/AkvhCLHY6M/Gf6X
F5M2SszScfqf83a0RQ8Tmkc2BDofFvFaeexvGkca1bxOqsw0sIfoJF8XBCuIoMNjIkfv267nQ4Rn
ftscvzii5JPy1oWMhQsOzmOCbXw5sFrwguMOJl6TgErUHFOW3dgLkgvhww7cBPXfzAyoMaP0IlrK
qygvxpIiuk3JCPc6tcL5OPeeik739VoL5mM0moGYE6JKMiphjQGz3IZhijy+AZNlTAhXWnZPHFxA
WtXVSn+TqbrjxV+E6wzFnfrd9P4JPjqP7Eut9x6qAhh0b1mX1gygUmVLH5gJXqW2q/FSzP4Y2HgF
8bdpDRthmo37JWcn7r4RhPOwLd+2LLmIu7qqI28BzYbJeQN5tHS4AhCMXsLVWto2jWoVOvlpApM4
UtusZbPkxui0VuSY9LENQAHQVEqwNYc7y3v2FLXJzWEnW/gCEGkb7SlrotsmESYViImkd2Eig8rP
C2bpCpRfUNPqGVEY9HpF/6FwS/pCgkzlfQTgdpgLH6bXfzTMMH5Jvgyu/XJNZbYPem1IcOZ93VXN
CasaAQKKGUOlmUdN46SGMKG6jig85VRW2+x8HgpRfkdPAFynwXjcrHspbbA9YlF+rKI+UhanybJo
kxHx+BLD+Wdr6zx+/v+eDkepszywJTPq7lUvup+QJEtP1DYsfqPjAq22vRqoKeJnzw5I87Wd/m/u
+NscuAVaFEU0vOOw/rHIUYAlETxv9ASEzg+Ci2N6yWP69OQG54UnzTREXNnLwJEqDZaRFe7mvCvX
PlYu7D/mo2JBTFNtMKerqs5AbQoEMP1gVhF0qgeFULx1cULTr4aL1EoXLKUJxo7yCoWEMHTgRHRy
mEPpsPwxq/dpQWOrU+0TlSpmU9OhDjbdi7EqnbnVS+Ya8o04wdvVABEBoFG+RH8nyhZ7D3fK0k0r
PJsw1zI3w9bB9r8N45waviF8rVn0XFqs+bC/rlFC3rE4gIRyd01Sgg2Vp5djgGBIFHypHsP4aFhO
6XNBvllbYtND7ECFA2nwkSWJur3e9ckueArxx6Y4UbUoc/ZNfs4GQwx66yA+lY7Zay8tW0r741MX
bVeZOQCATD9kkB/oUrYUftjQd6TlYkUObQRAvKtFm2xsZhsFQn8GNs0qFDSvo3hGtmdbY4k8ptOa
E6u9Bf/KTGelNvwyPwZE7oLSewqTfcThyeEZFeRrlpHZr7b7MgBE1x1rBRYFj0btg740dNz7uzIT
/g7yZsoe0KTxwXPSX5Z8cOUUl6644UjHtRbfTvwYipiGywWlPabhQofd5FaTr2PUa3iz2h5WFiDx
9XVnF8tWtxXcffcUJrvxpITnu+MoT/70LPAucwsJHE/P/+elgrqW03Sd6Yml0cawusAqpAEscI8H
0yH6Ji0/9N3XK7kKgAlQTcTyYO3pWqgWgOBEr0PiQ6yVEWTYELN0UxxCtMh+La6j6XiCMk8nHtf7
1O5RkRHl1+ddM+hekt8Zy9EnLjIKVx+6XkLzhkY4C8Xpy39SSQ/SURmDRJkGPiPDpyotYCNePNiP
sNBitaT1zm7QU8uhMml4Fxv1J6lBMzy23NhQMcxGie9C51yJyLA3plLN4xI11ew3f1cAgsjjBbp0
LA/KYizJsxZUYTARe4q50wAdEjTqePuqmEWu16VxYxQngQRTKYj3FGivJhkIHG/jj+IYwtHdKZzf
WnHwyKSl3QlHkYHxRCNX5YAgTAkXG8mNjoooE200nC9ubdTVbNej9d93evAGTOpojxq45ntco71e
ne/JQYQytYhYWyBDX31PZEpy5fBlWoRVDtJmI49kL6jtTTTscxcCPsLK3yzsPg0Xf1lpHB5hzJEJ
/V67bkG2JvAmIP9QbeNGLqC4stdPh8/XJJJSNcYfUd2YApplzNXDCX7csgE0ULmIN7MtqryJK8Z+
CngmSx/0ShQAksVAoqzUZAMEET6w/9q/KpMdVnozF8RwNn4JawyLt7Hyt1gVAHXcVEC02kg/lgOt
xZDQWrOcE2+RAgxMihdQTjQMsjVgs/wh/vWxRNcSIOWyCaZ8KSlN3mAH2iU7gwIm52bWlA/G38KC
G8QFBCHuatXC/fEsbFeK7oYMDut6JFJE5xdfzN7/XU65x/Wz3v2DhkIEMRTQugPLxkgSI46NzPOe
gqgNS85FC487n15Qlh6pddnn4zZT3lwMWPGr5jwadjLDIqHS84Yi6EhshuKvkhWNkYCAb+PQK5Qw
lCO9B4HunGhHuD5rmwuFS9c6ogmA8CZ0Rq4YLTUgvE57540VuOQrDN3k+0qS0gGcVBPn9y6kikmB
gmdVnP36Cy/+HLq8NHgNP1kdpcs1/SYdd83BEgkKWyGqAx42cLK1wl8f5hdcm4bvXPAXa4dMHHS+
L7UEPzIVQ+PL8sRUM23jcr2I9sRu5+RlgxUTzPNgh05srcBzzJdVkTjonpR6sprgq4oh1wk49T10
673wKHcdGzAoqnHugZbVmXTpkd7DF+IYdmOxwtpzNpAvkfdjp6B5uOY57FrVCEtjdfr3ztiXRq3e
Zxi2fH28GRrY9f90PCbDsmxKMK/Hdh1Yna2X1BxjwZtvGelI/E6ubIF5PNmkc6qxG/1kdPQM8JVl
Y+a1QxRfdlMEI3pnetyi2JqtWUcVoSJfES2N6PuzkfR46WWkbLLwGmYhJ8KFJ/auLBVkzkNZZ5HS
5uCpBqBQpYzfrdZs3avoR1pJIf03Q7kwMUMvpWB7Hbi5pZmO9pa+96fJmAviq2D5VDburHdImvbV
MAJx6FKbStRoOcZMj5cH67xjIZYyRZYG/Kiz5WGkI0uhwX2cPWeFAjXpEgrPB9LUxwyLG2CrzgTz
z5yMkOXzDQ032u0VRQv0VhVi3LGVlsjfzcU3Hjh7bu+7CcWoX3d5L8xH6aYZQbA2iK9HM4cn+yVS
Z2jkJ8POH30LkiXueG60x9FCa/p6DHtvudWPf/zNkKzfrhwXZCEDFSXfYNO/DZ3eGZUmp9gsjzp4
3wMiPtIlg53oy7Et46cW2wL+hI2WsRcnuqwUhwYlmCuR2bj7JXURTrLLWugdlQdtjCj7ZyjalztF
WpBD3P+c0X58WbFH7pG2SminPnCXjUKTQ4yppu0MLERDBI6DFmTpLknQzf6xIO6ludMTVcqi13St
aAXl3labXKvbiRHsQGydim4BfBv0hHvDiV5EepfTWXRorDENlQIQPDoqRhMJHIDmHkegd+khByoX
9SHhtGla8xv2Sf8GCT7iO2S3huUC2SCQU3fy80T/mbD/iSZDxuRuNak8QAyKN4duvyVWoqfXjv1K
2VONlaSRwiYUMaraxgrp7ovvzS5ZjyydsEKqQsKpUst+IbBhSALxrVBtYHa43lAFCCijSPc69zR4
ieOrE5XRSZ54ec5W6Cwkqgp6kUKWDUaXh4eOw2WgzpcB3HGzHYsLfpIwQZSBpvSbq1R2rRNoRufM
wAMo5sGIdcJ9Y9aRkhUh5xbwhulRRt5OmesBnLUyncUTA9igVccBIzKdISctLxPufotlP5dKqvb7
Ws/QOznWOa9ZFdnxM4k5ALOGoiPWNXo/wmy/m88fpISc3PfVfnWFyDFXtCpoxx7sJUp2B4TpFLUT
QqmF9bjZbGMi8BssWQwHeHPXd27qv+wDTktLPnCSUdd365/j73V7C/0uESg4dHJmZplGQ3zjJYCU
SdUxE3WKbAEIqSZoOe3vtBIAEfkNM4EXNUTUKW43LovLCO49Ep6MpjB4QYswkRHA3/Unushwsiey
4kynWpntExdJhgDbgmhDtb1dOkn4WiiEKP0NvU4D8lBJhMG8suaoJyUKMo4tXo9vVDeC7b+dPKld
KGozzQjSXmOktIGmDJip38tfHVGlngwvkyZUmq/lZ0dqtfybrm+tmvriOoBiBACAgDy9lQro45id
Z3/C3zYzFz8zBxCqyU0qS0194GPO1RmS6tEt2+tcnMRAQSVKIS1CdYYOd50kWNPGzKbpF0gF6urG
u9F1t3L2FO0fKshvRuvPzex8wqFlM/wAs6IpRHicbiKTxX3VAA0WjriEq0/ZNv6AR+YUM0QNNB/6
L7Z6/bEuuUfya9DvxcxPjjCxxsA28OCPXlQ3PBJNp02GaFlPpbq67aKJHW3R4FVJhg7pFdZ+IEFa
vhuGQeNi6VjpAq/eOAs/1JCFvPcqWWJpCxVHAEjFvfy0DsA6TCwULD0Z9FSknMspcEl3Dsmd3iUx
cNCURFJirztyPvd8Gq4ZYaab2W1jmSBoQEm4IpEIzo+xilQQPn6xBB6gy9k26iisVxsQr/GH/mge
rGG8LT3rKmvqWDWyu/2D/JCt44PSD8Y1nXO4Yy6SYwK9QidgLKcVgK4DtddgM+HSDSerd1S8stLt
rpEvvLZIEnr/Q87yGOBJPhdRqtR4SOUkLH80V1vwUH+GxC3YTHKLzkP20Y8oF5SriPoxMcvPBbKS
n3U8ty5l7Pmlg1RXePtsrfu8Gb5yucFuZCxWbN6PnJurvTpcbacPkLfoM9wGrBXRm76C7mvgdKrP
SGW05qjp27LBh288M8Z8hmytbqO8/CyxYmYV9DJ6ssbrj2ZcwEcQOPXNT7xnqZChhMHWlONHalAm
gejl/b4dvx2k/NqK7APkjuCM9MC/JPYnMZtkxEsj8L5q9MIwzQpwvZhjb7RWE0R8yHVCHwRrbdAn
SGnQzigxmp1Ge8jf8QRaaOsxJnzWy2vngqEV5IZqzO7XMP5aY0qAFrbAwQWn3FLorUNtrFnt8ELK
vsVT74z4o/m2ujXgBI28wgZRxHw6ezRxgvZhNK2+BHJU58Qf18iz7HJm+nxmTNf0ypIr57Nvma2z
lo2rmOVqWjh7jeWZd5/YOuwKxI2Bw90Y5NdV8vVe57jqUChsyPFItEa8u1eUk3DQVtLeLZTvKNRB
lLmS96upNZllyz4NmE3exxCccp/qT7K6FwDeNeaMZYJTO0oX+SziltsZtlqe+XuQV4+maHeX76Rj
REWWF7Js0yPRKQSLEpGdTW89rjFQytBzMemhBDenaUxxwgZi0JCJ21HywcOm9cm55eOyAO52qEf0
Nc/QjY5xQ49SacSSRZyhLlG3YEwqejlajFDRmg+JnHUjx3er/CsbPT4hlbboTkhzaZHU+b+9e3Zg
LTZndRtX7RKuQ6AETLU2vkmXftvow7iP+F6i5U8b17AcvuFCgqLmztVJBrlEji0dMH0pFUnshxgE
c2uqVDj4GvZxGOr4DIxTdobisQYo8IDqLxjTRzZvGjPW+pUbiMpj3kLqUng4ALLoS4+hD4qe6Kh0
6gd4qrd2butHrNE3o0N63uZI59ezzcTK434TassZOPK/KlopXSOxgCTDqiBqkrM9FOe9HOY6j3Ar
MpVec94dFgWh+Opi6mJdfhhl1cSoTEB0+BBuFa3+Ye2FvC0enr+I4cLO7U/ECi0M1KPIIB9ItOmM
JjkbbPytd60MWnd4ejMZF7ZLf3WjF9MMW4LIWfmNMQuVFHeZYTyGiM7/O6el3/1ZSICfqezpCMsN
A5Aa/lxJyLyWAFSmaknrvpjZdX9uQH+CPCKc8A8EhwuWmWos97wK+zEz6dSg8sc8TIP3q1ixy2j8
ClDdppzr3dwr+FpNYRaLq9RsFKcIe+QbuXqWKjSfUDaOc79XvE4BRxvcdjv7RHckq32tK20/Bf7p
9C/Sy3QnYvKi9Nyr8ZlCJH/2uPhNWkomFcaka43pk8c8lYNo6e1vrugl3TLhJkb4Bo+QkDvE++5T
s46LrKUTAzkWWILA6+IYGO0xt0DAGoZTmTxieNN3it1YeuYbL1EvMFAOFkfKS8RqI6r3oPDj+sP4
Bb8vZ4Fcp9UXSEauDoaCmcOstZ6+ry6Mao43pnYb4MfzuMEqt2M5R3zssow5YIVZFSvxAOrglqAd
awN0N46Uw48EmpcIlWvePm8e9MfJ5dv7zJyzNaeFzll8lFG7pu804hmcDSlOIJABl0LQ1MeUmwYd
5ihNuy7X034XW338o6hBMNgsmBvHum/DNp12mcTIJl6VoI5RCM9m9bZQjHl7QSrQi+25oJdGNwwP
vbFSLoIB7G3l5ZeGd1lbsDBO5wkXwJgoqCeAcIqpyFOtJFyfoy9b/uiOm1/3NdWrY0oOOGGOhE2G
DpQUsFwev1CI81gSJZxYr2B03RhKq9vRUq+xVLuxqnXJJAuZtZ2q9pXA73QbWOqCSXTWIJPSz/15
0x6lWksOgVlc7FQtppjMpurm6IGPpdAS44P3ikt2wxdWnMm3EKW4K6HNk+AaUDXIfKD4OWoncs2t
9S5kmljSRXioljSNQAGCNN0wiBvDx5vpz/dVldqX4rXdLzJbTJepUZuUuOsi6vyPBFPjAKtPuAjb
oyDaMkYkwGWaXGNbEM3dvm4H2a+XRe3Yt0I7l8CePadxmpXm0ixsbi0YJzA0SvCuLxvAjxhyt6jf
3ZkubfOiOXDEtCCAi5O2T2mOfmsHlWHFcV+sAUNBhuOjKjLU0wyoI+wrCkQ00NvwmJnq4zMHLaj2
qT+HbdHXwD6lFmpHekmCm0yKLI/aBLmG3nlaRrB8qKXTEAahc0DBz1Ykv56n4lU8hZcSiNX1zXWI
XThE+eXktgfTctGfy8bHcvtR103wijnpCksmfJYTk15gIAw5R3EX/ilElJN6cGFd+d3BhONlSbDu
EmoGCSzom9eSlPZS7NwzwawRP7SoYfhXhBu1hlWf2jqBXRKRV7BPRi6bXVO+52HELOIP+ORyYM+d
FLb0eTn5cX3Em58Tx5Y3oKZkfmM8sLaJwJCD94oZvoKhH9PyTX3JQcR362wLBnc5Vvc4hiCByOmC
Sgb7stsU/VH/rJMxf1K7Vy4MmAD0oRf+45+Gn+gUYjHC0r5qNxFtl8xYmeLP1D1KGjWoYo6aNFp7
WSoW1nu1j39DpncGnUmVOzZB0+3hVL90A2i+qvokKisbUooIvhutY1DlaO5GsQflfUef3Wn/8u4x
4/V7rFbkiHW9odiMEGwzKG/VFa50Hgd7mm+dtaw9qnyjXr7qXKD18Qd2eOjYOaIkk8PBX1oKSiCE
ahBfyQ7aR0RlqxzPQ68fWgiLy3NBD14ML20+vX7JJzAQWCbNUoCDFqhWL0PxMtWM1906Ip2ZgGWk
ngnyZHDGlEky62XG3DdpZ3doMBbL4hHFIAVFnaL8fBVydwQDmXSZpuxKjDAepL43UJQXjl/SijD/
tVp3SyZoxMGWHSdTZAqD2OrCCVPdERjTrUa/JXaq26GXL1GjFyqczLc/FknIIQF+8kNYJfxJ1TtZ
KK3YLWF7TMOmQQT4HICZo3V9AfDyFBL8azZTbu4MS7ZAPs/GgbeHh9qnXZcywt3+5IXg+z4WiYGR
9YbfsYoGGLOAIa+/9whDxhNBMwYAahrQLkGZW/L/4l3L66KCH9jMyXxV0+u9FY3eiBlx9phNu52E
2tUUaJejY8tMrM9xtzu2SWPIPq4MnOHXBpsEGXMKurJB9dHricEfQYtO8ksx2eStY9G73Iw+2vC4
DiOUzP+fuvDrqO9U8KGsDmBr8vaWM6OUdcRJYh0GvaRY0oDmfsFUj4nbkTTftFcgRgrBn9A5+kfa
7nQuM3PtHDhRkWESQxCkEE/RMUCvxFhDA1E6YbHE66mOF+btw/ur6J2Upg812O2Wk5qxBkYTpSCm
C09Kgl+ycAoEUcNF+pu3+rfeV4igZAsOwYbMQxAHLZUWfSZfJHjRqO4Ig2+EAxMw5ENxfxXZt9s3
2Rvl9cU8sPB4pMRJi878Fwc/JRXqTjCVGgsoE5s2XU23x/rZJFxtmW4YbsHcP2Rl35xGH0pscoX6
HfH7XdW7favja2+PMI6986RoK23/g7TdgOaayRAY8ioZ0Pm6sr6IZPxj9pSnNmGdGyQiLW8IIWOj
gpIroi919PYXxdg5JtFjiulZ3Qs5W+FPolB+2ItfOKxGVwoahpRk7OwaQLUUfYsZ152ckkbx8xSM
O6Syts0+/XsXUqbZ9zykuPrQwo+DY103BaEXScMldb+Z+cytl1s9Rxwopq90pA9i7nlSJkIA2m8f
07DistN+B4GqzSIb/Mj54WvDvRNzQ1AQmqnbD3MBGEAbZcUyPNV4PywK0qu180SvJf9HDAk/J6NX
HT2OOF4sDVZ5r4HIpB/LKtj4JMlt5JayW++yOoTAejqJwDu7CCsJcScJBfD3a+9r/q/4AKFzUTX8
coWh+JWpc9FUQ+bi3NusBXPqNFaNuKTKTANwdZI3NWen8t93wD0EUzir/p31g8ZY/EKvIInSh1jH
JBkmaSif7+MZ2gLCMy4ku1+osGhaj8SgGfbSlwNNn1yMtjE3MLB/OWgWuLznHsvbmbXq3TRRkaZw
750Ko/BfttU52wkq90aOJxHu+ZktksEilQ3T8Uz5ZJtdbez2RihFD+7WCjs2CKWs/FZy5bMOJZM/
HARk6/vIxRvvw+wtdfblfMGFO5xcYicZ/WJ91qCBCUqgdq2zkfFJ6Np4hPcOrw8mFHBkQL1OmDyD
xgfiwfYgw+uARH0EhlUM5nzvIwIyQ3hmz5dnazucJGERCGsYQP93W9Sy1S98H5dLxGX9Nm61oxnV
HCwR0IIkZeyto+j+ejBBOPQI12AYdgXTC3XjedgHEuLzqSDpZm/jeW1itJlAjl8KB1TOutExXhRs
7QATeTO/HFOMUEefgki+V9GnRdVT2dy/I8BPWYQWe98dvlr5nqFJsifWUHCnELlbiCL1WB2YXYuc
c0+pwHPaehHPkxjqnAlWCjXJV/EmgTN+NW4ZI6WRaYl1dMGE3/RlDMllepOMYqidcUvjcDitloHc
ARN8EdK+J2Q3lQFIVWCtDZD11Syi8V7LijJBkFYBMV7KhXPMTrkgTAJ+FQyJBv3KbGOFjW9qj5bO
BeRZsWlNZVQLBB/quaWbzm+MohN+SPHty7uWylID85CEi+b9aJ3KXtt5HAuncD0sPohBKtAVxpri
JpbtDxhjc7zY2dI1/uho+yT2tOVcM2qDL8b/iynDisfOj/WI5oZJMLZ6AkqZwWjpGn1pnSPqDn0r
fjbHmMR/VpoN0+rPPUGAenyIL2UHbcC/4eS6iIoWX0D+vP4aSGXFegF6bvfdf3vTlEt0OR3jqu3q
gGPwkPMFX5iDtknmkaD4s6Wvdm4zp5tt8XmhiyM4EMnkvQyYZQYIZqpRSwWnDpdIKMbnAYEbKtnN
2aNpvvlygCZBJpO0muUVUmC9tjkSzL9PtENQJMZgD53VKcHayZtxAV1fj5OLMUGO4UEaVTVBH9Ck
fdZY93zXESu97y7wKc1YPXclzfJAr2IB4aZfSyK1A/jiQhhb5X3AaGXI2I/iAmHpSwCtXhskidWI
+RMs0zHKarSQqLA7TLvSMOAWh3Z63XyETrQO5QWa+mTiaDQVpFT0zXaezo5JYmv5QWQSWMgQAFYc
Erp4k4UFej8iJZF/L+UhetUDc0WlhTm4QBdbVlwcWvQkkC6pWydDHJZ7reNSStn/MS7X3Fso6sFi
jUF1+C30ssKxNu69APg530wLWleF0nFSNm4jip5j222/+XMRObJNcA2uKfhnrsfNFe6LchJiw+x7
2VVydv3s4SMrMhBVUnm7JZgZw4zB8Ca9TLOwmh4zaLgDddhLkHq3RGTzVjB/Y2Orhp24rMDCfNah
wTnqcxT8p2smKwOkM5snoW/QHMIeF7mnhV4OTkqxHm0dscgmFwi2NLfXsE1+gGzIfQBNYFa/ABcZ
A2ABwRD5/Dq/lI+RSUVuRSNNqVF6xU+3OnKGMvQJmjL55gwSlMD1DpWc+0903fzaNOOLXBcxaV5z
JR9lCFNCGlrC5uYb782HMxRmIBLmEkiQzHGBWsAP472jus51o6q7K255UjvfoocdHr03D0InTRKN
67Q1LX+fLtYy0OHhWXO5jFXgsg7eyi927IOws9jbMu4kkr1nUvumL8QY3GtU2n1MvcFVMXkAuyVt
yA/RBJgk51IlnGwzCy5JHYDWMoW6J+N/JH76+J5dphNj9fOynrbxYX2Il+JM2uOzGYJ1Y5JtdxHr
qxmkk1F7opAI3ubIuVmLYW1R54FuZML/giw0J4Qq7w7jaHI7fSOltTRfxz+TjBZbSD4+auIl++kb
LC+mCiDlvqs+IwDw6XQXhlhIevNShPosA1SJqSxXeyxbuSpPR/PpraeSEOHUkkATj9K76HiKKxmd
I9JRJ4y4ji8jR6SjjLT2O6noA2lFBXS7x5yZIHKFlhQrS3GiM3shg5KJ/UumFGQoVV5aewBA1hro
4JDyYPRUxSc1J0bH5/TbMOn+0zyfCr6NLmlTw/2t0Ptqz27K2WU5i/WG9an42Y/ELs1NghQLOgFE
e1/Gozq2XGkAyLfyYd+jerqpq2GQqORtB+9QollauKlc7o/gQwd5cyBtMKu5rL/uUaSO9HfBBCne
Qz53uC2r5HrCnrbfHJuFbz9EDCd2LGuJQqaE9VDlaFBjc1Wqdhwvb0G9RrQf0U5/WB1PvKUGQF1U
oBNx48jEZNS1VTr6pEY+KAzfXo5mKV1iUUJcqELLrQJ+e2HWBn+z+P7QX+LAbir9uBRPnlKF2kJH
GcJoEQ4qwTHg0fFA7/falz0y7txgJdlur2WA66NBJwNEkkiYqi1/H3HJyfkmht3pXPojyyV95kue
t5l/wzIJ6eHULGnP4MAcL8GUPKGgbRthXg21A1oLbQrCEeT8peKECaT5bsdWBjG9q77UGkxsajwY
OSexeOebBwXCV7hh7SkHuf8KDkxKkvCituuG7334JpyERLPyv576Hyp13UmZ1udZwoeKQQxV1/lC
1FsHW553BI+RM8nLV1BGl9BH3kWlf3pLMpSHJecCZgMfLgdptJSxTYgVP0mWqXQXJ4kakJ7W8YlW
NBDSzIyo5NTXTWUOtILzJCjGljJW5WI2NbIQegdFaXfBxwPwZ4e2eZjhVnJSEHsV1hmJ6Kc2Zfvb
6AFugjh6t2wYpfvO+pU7Rz3DCDYX80D5iK1+nhpsyJsLl/H1qa8I5Cnhfb4f7nH9faCF/Kjf22mw
21mYVWaD8UPbiAew7k3tZ3ZGaDurEn8Dq9siKRRKo7QQIPDZ+11NYpzqZ3zkMOLTDq+HYFw2a9bp
iR74rdmFuj0scBdzEePX8L/4CV/lV0vogd+zQ5KWRLnWEllO+OKElAvfWC5Ase3wFTPG8/KaFFim
O0/OuXrVuwtdOOuSadVUgxw5zh9VCaAslsujtjdmRnkxHnWb/Injaywxrwcl0WOPjoRbnXs3jNlW
nCZ2W7r5tXVyVxrN81pCpIM7ZNKg7Jh+gI0irM3dqAvSzmK6dvWt53jQBPbcxIF0ufgNGqcvrr49
N/y/yaMYMgzy8w5Ws4fiQN1oYrR9z6mdKYFBiHrMXJga9o5VqsQxQN2HbZSmpLSJSnaVINqIQlUY
HD43wxf5mKen6IlWb3yqjc7yDytc4vS3lLIXJMvyfFvO4o6EN5Mxv4+HBxMuSaTh9fyff62YoA+a
JBD2KpN74eD0qj78TjTtvyMsereS+ZmetzpOV7fZT1MlKfgg76gTTEg9eOrDpNHA7CniPiB7q987
Bf0ONit1OaKqigWlJzUJULfRS+KPBcoW7f7otCx1zjEGuV9TlUcKdRkBMc0QvRc5HGZQBiP5yQAY
sVjk58+xQQ0H8vBCs6NjQzKYa59jqosVyqNcZSRsjZCYvAVFpBSVW2tvoErXHi2/3qbyYmXrOz6k
6x8VYHUx34DVhl012OLwuGyyzlBS67paaJFTLP5PZ8UvjRiLnDV+ZsVxLzRDUPWDILNwt4sBFP6s
TA5ge9IH5KSWGvpBDjwUZXTXqUnR/b5AbiAfxhIM2dF4JQwc8IJIkwc3gfxgApjg41ARDPg/mJfM
kVU+Cgac8puRaRPuVscqgEZWXbK5X+KvjJq26+H4jNdcjSEJH4ukKN4JsgbVtxKRBM7jgbm2Ot9m
pFNY8ss74q7M4Os2jECAZetic95DXPxyHmrM0rQGR10pHblwQ9PYqg+zpuqszMPSNTHqDqWwrUrH
Oy2L4xFF2yNQtukg2BjlfCEeENLCzpgFACCgrTOZ/u7vj7VY7bQVyaH2UX+fPKRxWRdkKB+955v9
BfIWF/FgH47D0eQlScdfkxfzqSEnAVdVPugBokfENgjXYcsr9Ah0tWbJPJTfMo6bt62tPKet4erd
mD2SxdA/j2Tgp+rKIPhbPZf7Ts1fDEV9vLweGyVFy2PUZkcuMIRGBT71kjgNEWGjqirfS6q3kO9S
JsmpbVvKU3E69eXjocVJAeA/ZxIXduNUusnEMnhbtSkX+LxQFSjzDxlID6uJyneZI0y8Y9RQ8DzE
mSCiFHhzqZdSjEGGzADqYm6fqzPv7T/YxVxwZ7wCe162rHTB9dl8uK384Jci+QgFq0M2KSBBpKGu
4JJ6X9BgnWzScwnLdSHwfagjxas5OgejAB5O+JX4tw8ThyvMMrST42UkWQVtE9xU72jqERoJS276
QOku2EftP/Pz/bZpgcjsTD/d1R65/J2+rsCrq1Pn6HW2Tf7FujLg97xv3Hs9kkJTDDVhZL41whUb
s9hYFxHvoRO6Bkz+43lhiuO8OBHQMIrAbj/RotzBSUt3kkpc3Pxgidx/a5U4EtREOXL0q3lbp/VK
vBRv2J+2v3Q4tN76f+7DV+mXOW9p3xXGljwgcVJg+bxQ6U8r7snRwmU6NIM14Kx+3W2Pbm1CRk9X
SrfXZtowtxmAZ9KGJDD26Klf0rd3aJ3ZA9wJ1f8+9xTmhc6wDzmM0SQDPRK22jDVGK8N/BOaSxcF
t+Nug8SH0Cwb0fVoXn6ZEMlQoln/jpJFnsAofmS5IsLbjxrh4hnSQ8PjA7gKRbCad1udxXS6/CJx
5j9bbllHRCICcT8mXgTSn0UNcDtSC3hRXTNaLp/jKNz5cMwfHChcexMNPwesdZRYvzsSeIYcdUm9
1N4E3Ms2M782dmc6sS9bZBd7MM+ky42TPnBAIN1NqgWJxemmN0sJlrb9+/LDriKZh7LCYQLq67oV
GWXmb6EFXnUBA9cK7AXOSFRos6m3Sf79sXnDuqdmWUV/QoSb5R/2uaCRb+sIH9kcX29yB19e/tsH
m13Rd6MRUp0cPKBRRNwMGKb2cenoKyfCxLsO2k39psIG4Rq1j19+xCCKnRLzBWUPugQvcVa9A8IN
slQnw1IjgoXnfUlx1oeDa1qbgDxxTOs5qS6cKe0FJIHjOQM59gsena2Zx8+rzfeGcpcUK16/YiOK
RfN4GqUfp9eaK9hvJ4d1m7c0CyLFGekmq5cEL2xrVPwZnzY7i5OW2dddvApY7Lit8R78K/LOibQu
8831plwiSE38kZ1Z7PynFCq37u304wwiFTf7KuyynMCY9il0qUHqjs9j5d06IREONEhwuC0epzqK
m+Cs9cPR8gKwNFOu9hCA1IGMa7MxNdONl6ufK5WQNKmKBwfsox5NaENPBU/PtEU+4f5epE9BOyKS
fG7Hl/caE7l0G15XR++6CXlBPPVD8wvOBMOjfufVimGdBE0DkQpzFsQ8PjAya/yq8qCrqdpohyKE
PZRsHHIi05y1xo8TUtUNmcoSTMDrFfeGaaZgi8+rbZ0NxzJCRBENkRHEYqEp1t5thG/DFNyd02t9
ky/0NUCZl3+Zfcgpr9NwbBzws9AhrV6pJJ/IQ/2TJZBCR3jNwKT6o5DBVcPDXCY5ktvE/FfjWxkv
nLtpdc5aigBXUpElSkWWH1mUFhg66LXtmrmsBywoMOPVFBjbzmoxFSAtMD4UIpgyx6gHOB63SWlO
dYuOPgSIVZGSKObo4gRIUDojBecdy3TP6YSDvKsB3zlCoMyrdEhnzMl2K4vehv5Aq2mXyMDS3Uva
YcqkfWPOwhu66x83F2f083PjjR0LjG7VOWYdavGaMup30TcG3TiAL1TZA9XCbgFQWK5kwtnjx+II
ienmkkTzLAHBR8RG/iJhmMiUK+VilEoOfEQ2IXbuAii7nRHaVZ1m22hR+Yaryvo5EVyaaEXnTpSV
efKhCW2A/NMhUQvn7vFlYKCswUYpzANrfsDxpiQXNXpgN1xW4SYZBboIL4dQmIO17GwKgA38mTA+
nCQJVGXg2fy+IrMCWdsLDFD8Hqlzsp4IjUJ3hMUxmVdZbbiggWLPalAGIVIwy00C6dHxU/p3sn5d
4AoIZZWTrdDOQKK2VXja5zul4NibhWx7JKmT6GnpmUGK6iJzn+851QYuiFHO3AjT2uVkxRR9dpbr
z2J5ey6VPPXG8bj95WGzqPydq6N3vdyNHVlJfcte3Sns/7X/vX7wUuU6noS+M++ZNiK8/DZ8QA//
e4tQ01Kvy3BtwMH3HEY4ijKvYkOjuNUkCZi8XDz/PvwN8e4IoQLUTivdk3uj1NEb9QlrXbVpJFFJ
Xqt3vDZsNHsGzbmo8/ZjiAHouKSR8NUfDIpcNiz3lATBR5JrFi5d7GZ03901Y2DBP+9jmrv6BaBV
EB+WXKsf0X3F7sl8yPebrGCqGPZLOxqwZxr9T/AQX6pHbcytNuAMxLxyEnj/7uKDT96Zwc4TImCL
r1Q66jqaYCnSlwyop45mZ+4wRI3Sb3nH+GmYphyNoeA+VbB5fEQfeuuB9nG42sColLn+3jnmnoAZ
99Z92p2mPD+9QfWYX9qqvpPXwVeoE8Rbm+VGwcMcQSj+UCIE0N6TiWk+zh7Lj7kxrfJIbw1hz7bK
AW1CtzMipHAXqljthG7VTbo1dpCs+/ES5ucN8PxCSv60eDESFpafT8ucAHyiwW2adbwkQ7ZjzH7O
Cv0sfM6TS4B9HKT033cKLe2ZENwX9rauUBePfuMMcYmpISxYtFC5mJTRLRJWNl08r4s3JB/UreNd
64ven9Lbe5l4BtyFo9wlyL2/7LY/J/W4Mk39UIxRM2SzhJG8tpwmwDawzi57UUbOUKqfYlALYcnB
ne+HLEJnd9CKYLqUQHa2A+uscVqnjXfIqVe+0gjdIcnVligIg+UdtU3wEHAqyY006CcVudnuPMaC
kQNB+piwZrpP6ZgciEOiGZZ5SfvIJRUX5fOpZV95hDSa2t/6xgEcceS4tQosmWqvWGkiiH9qTmIm
gefuF0cfvuMKAYWMQ+hPwcij4l5evzQSItiFHSkcJAdsNlI3TDF+qbB/KNdq2Dn5dlE4LLDbc0S0
G3vR5ySSFuYpOENOdhjYKanJ+RX+SrZzYjshac0ROYqD02E14Bt7aWPDh2zclZyB8GWjhKnfLmYm
O8GM9cxnMVKJVPFXiImA5LlKxzFy0F/IGtMg9jtxQwc//Abq2KufMsUHdY3g3leiyqSu+hk2kBhq
KtAMaASw9U0rnVucU9+A28/7nYOlIojL9RmysxSgoCC9JYjM8tFDCWzKVNabvJfbCit1lHYBZy/9
mpPhV7umlebXYIoXXtpCEmYfO/4OgL/ubSDrspBBnqITnfRwi8euiNxW5in/FY5zb9voWM+Bmw9j
qFynLUtsQd/sMQ0b7JsAhK1hT3R8jqxZ8WxbwbHjaKNcMDV9gFLBCqaBP1tiXQFsgncXDWG3Enpa
l0P2I9FCWSuZhBjt3xFM+1kydBOSW9xRLNTkXR6iTCWcrvTj2q+csaYhzkEvA7PVZwojTR4IThoP
X5JAOUBqYT33lz2v3xl5cnkIfu54KCAnKAPcq5pyMPH0q0Zbn8EM61TXczfQJouI+TQYUYuBZgr1
fPMJ8pvEcatLMvwRX6gnqoH8/thR2DyO31b+A+0kLObCEY/+ihDaj2VdgoOyjV8NaGVwVG94cdKy
F7o4njZuOpvP2cz/H1A7C4hU4OwXESfqq80gmQ8DY8ke99GKuTLMw+EUBAPHLn7wlktrf5+M68DL
3ltUH9Ff/5PkGA9YgvM937QZt9Och9/9Zkw+RzhSDL0sDGAI9xRZVFGaCcJR7klF7ZgNSHp09LU6
Agg48IZoodq98s6RrzwhhWfVLNGapW//1Z84IVOkOyovuaZefZAy7nPkwqf2kzC2KOldcSK+o/J1
h+QDE9pxVEq/+wk2H1yhgglWkAaGDT6QJHQ+bosaGD/hNpEgWHKxVJHzLf4CcWrmHo9pJmf6YhnK
ZDwyumGnAJKMvlSI/Vukw1XUayrOWLsGmf3oInt2O9BUSZqjLDmt4KuOv+a2kkEWcPIGqII9CqH+
7i3MbJGunhDSX1RIKB4jZ/51DOzYXu6+4o0Evp+R+l8cKpF4dN9OWWlHlKDnqd+ikVulJVycE0P6
4u1f7TmVfoZiHod1Np3brGMpn7HfolYJ0FIhQGt5+HKg+poiw+yrmAgTj/LMZ84ArtPhangt2hM/
zocRC9niwxVlEPzkxUPGoh4J4WuqzXh7rws8qnFJfwrddcBQS8f6jS7mRP2oPOhw7CYcctnMQzzU
MjAZII1SmF9mtIj4p777IQF1js+UTFCnDMK3eP4m8b8U/Hd+qMW8xrlSADfGs3eWDlhVkr8ORnD3
F7oLyrBiVz98NXqTEFwWr6fmF8BMZ+hw9BBIn7xhDK/VoMcLQtOX2Pu9yZgY4S4XkYme9bvcYRbE
z0VpKEkB2E3uoUt5IgRW4pVzdzVbOrihPbKG3jhdqdi1jFnkw/IQn5dJebe+gg14SAbsJVN9or3p
ZenVUKAHssO1yyZHbx6yulHtjsQZcFXlxmAI3nIzgvlBr6JSed+8trX4a0EK+xph+aeWiPZm3NK0
aj/y/TOvm0PoBb2YLhU8yYURCN5q4lJ5TdLTp0Z8Z+E4HP5nbNbpOhPjJ1teHau2H6dQU+QmbVm1
5BT4eqT2Tedp8haG9BhyZbTCbPBsD6RJPBbtP+DgEoyfmdkiTsLp1goT7R0XCMEJliO7P13Tp8Vf
z+hC/umg2KIWfJR8x7syNC0rEGJE30ektGSIDE5ug1qFhoEN6W9yBxg9F+3D1Hu48mwBCHpuiGf/
cGMTvmB2AZiKuirPW+TTFYmtzhxE0b/LMaUrEjkqMvj3gUGfbHbEZg8rgBd6iyp931KCPYpyxD1B
tkDu9GX1woSoN998vOkTQS11nSs+gzNNWjrAqkjJzMHuO+tKtmxjBuS6FrnpMGtvvg5mPInFnZVc
KZyqExRbHP912kiLwv/Ri//EAly+Wf+6zXsGmFSTx04JYICLpFwj+/DzRHHuD5MXBPShTUhnA+sR
oYJoy8RReQhV1WkJ3aVdnoDdl30qm+C7XDJ5/xwXDQ5ls1QKWpaAEIu6mm4H8+JraYsRGxV7MAiM
cpKkolzn0FmzFI4V/yeHXCDMrjDXAFUCmezwh4X9CddD66LHheV8kJJBPUvJLP9Marwr571EOQz6
TmSYAg7x3tXuErB/bpc2YoVx5g5bj0j+ZZMoBOMzA9alt5hq3u5zzoTXo+Fuv5LDKTWQWk34raGw
GrwdwEPqcyHTwlhOtN9zpPPJN9/LhJ/LQs6mcQBc4YWJBkpnnLdpIUlb1z70Gntvwl3SzINg6IC/
VIZbP2Zrllc8nQMzbaxoNy1ebAcR0n/WxsZvUGUt9U/aZClZxs+8naN+SUjnLjTh68bEkfu6X44Z
Dj5yBSpcr3m16KHKTvLMHkKdsV5M0LaSSVsMQHETAYpNoJdArL62egUpUjwlOVl1qINhUyJimTZq
LzB8VU4TIfLZvl7Z9sL4rgFlMBwKUn+t16mYrUtshA6V9lLiXH27ZQWsq5JDUPPs8v3hxNwyL4Nf
7/Kghyz4a5l6iP/sPH5Ln/XyjnuDpcdDIf2c8zrkDfXKuWuKXeA+bo+ZousO6zhMSXabgWbjRLNp
k1off3yh7qb/NEj2gRaFZNNMidxY5sWCbv1X9aTnX6Ud6+zDlcqu5L1mH1iyF5KnNzVpyw6UvVUR
695T0XZ4h7vAVkP++tbInEdfDXLOYwAP2koLIQkNZK/F3LxdCqv1qzru3kb3tXMxYCqWpwZeTD6M
JUH9VTQjfJ9U9ijOPY14Ra92PdHjPsLkr3ScwSaLkjPSSrbBA8GzrDOfntOwNRKECzR+nAi/yGVL
bzdt6vo5qwMieUUWAMFNDaiPGRMsACxB6rZ/ImheVv0eseGtfW0nmY7RGf6BgSEy4bQKN/1jvIpM
ud4cB9oBZr5hngn1wG/yk4D9iRl8fsNXe9tLsupZr69802jCnaHjFtFHI9qBJusOQRhQozJ1u981
0bz/YNOeeIFReqJpMBJd7mITIoX8gpJ+psaA/FEvBQWGpnrIuYczsPEgvTsND57bDS3OraUuUUzC
dmlP5JygB5/bnPdi+gWAR9AOh5e9o1DE3hUjJEKh829iYfMgVl40//sZ0Morn43BQqWIVZ8dLap9
6K+P0+fYCxsmPW4ALLqDhqDZW0e4PbVOz92dEbWu8Qd1zVURjB9IZJ0h7IDgz04C78GDvluOjVFE
Fc1Sw75dgimiiIauJ0ygE4YGzI+eeniO3WxNd6Izqze4Oxw2F5koG6W93sKt76PiQtof7CQWQBY3
CzTBy8mBBEcKkc4akQmaFNSTck8HoUUAMjwEsS6T47kNv++l+I+RMfAtkQteJcovlA6zBuSIzjmw
OHhjeY8+40HCi3P4ARXZ8dlUoGwdn32i29H44bup3eqglO5moiWGpf1ysw8o9ogtCsrjoMBJsLcH
sV3bvE5vBIFnA51LH3tFG4x4fp8Kskz7nHbXEfb5EYnz/PD8sQrnG0/9HSl09pJmSmhwc3iWNgTw
P7ljyxCaXTPwDqLSvbmXZF3g+tKjvAqKhf+ZF3CUTlTe3rtQzdB84Acawin/DpVhqMfU8o0SU2FG
GWZkv9RCHUAnUBExn1GRy2HGVlsgWV8HLEMC3ym6nK68HF+BmuKsRSpZg5I0KaiC3NcUNEarMFK+
dOUlHjJuwokgCttR05kPD/RynJFsE4s9QeTZ4j+wv82n573jDK1BE0O3uDOhHgo73+UW2BMwmAUU
GgBNzk8PfafPaJn9ldkZBnkC78S+Klkvw5vWld/5ZAbs6zgXehy+aa/rj8ZMAut37C2OqPhtfC/o
55HOpUyXZvZWmnXRZD0zL9WwovHsDy72SlybZSBj5Ji9xbd8C2psBsK+mXGU16OVqwRTJ7LUvo27
e5xDKP6XAE0zkb8DQ2SNIe08Uon9Go0KEjPhO0dcN7z7GahiPU0fOf7Lb0aNnzPr6FWFc968clEy
/qginWV3InafETHcoA+7OtIoJm87+jNs0fhbjhfUpM+4u4c8h45kl57KG1JLu5jx7yQMobxTGN++
KvKFoDGvIzXU9ryB1WY/WlWxjW3slfg/AxA3T2qTMw/4qTccmVAR+mVG3//N5oQohMYxYJwLA9u5
oji+1bFx+2JOgaLPwJmWG3m9vqmT80gxylQqaXa6sfQQWpxXtNeGwBgmVIxU1N5JbdHTko2xoQcb
by/NcFDpcDoQgi5FGKCdwZFvSowp8FqQCr1AQiJQjOsP2a5TQcwoZTB/sbaFe34z0HJiCSvnMo8B
RjQZ+TDGu36XZixTs8B/lJ58QZ/1Cvg6BXdg2chTAltQcynwHUhWZrCAr5HVuXV0eb+6JZ8qExNh
aqynnc026ka775Hy5hUVn0RkMy1R8qofu56vm9ALved97CeOFzZB/3VumGfMU1UbAOGPLP9Tk3yP
iMDf4852LYilQTEDbj7iaZBWxBXtXDSO8oon83f9yIk08tnWHiangYEOKL17txfiDvsNUJDwjroo
KkF6331cjHHO9YFcmHj5w92XIyFoKNUvgb15T6CbEn3osdfTsbMmKLitj15csVmkt6k2H7s8mSD8
yT+2m9ESM4dJUGrWjtMbwUlqd3ZHjIg4y2ZrWSpZLZ6QCp2R8XubG5pW0RUvnn8zDJ22RuUEHDhJ
QNwC/1OkylG9/6vhW27Ydr1yU7lzlmGJwxn1fYwLsBNVWxjk6t956aS+LLRcTBv/Wry/sgcNpb8N
1rYNq9jAob7SoZsdxCocPnbfjCkNVsCiccdT3PJ0f0S54uAsOutXwWnOK/hdTn+KVcr/E4ObU6yk
ET6hyZ+1LsndMH77rotToPCxZJHdM7s+LKvzRKgiyvj75GfjeZSHqLG4ME0Q0I/C2XguOfeF3Dqd
j17wPPBSEJOsUp0NSS5WX5uFqz9WjliTiHQrDSNtUCJ/yyWrK+L93D7449HhIETJn7d3Y9KcLPvl
mQVniKj8JrIb0esM5qn2S6n9SS5RQhtQYaJx9loZ9DIhV7nCozFjpDchqZeQ38VJzPuZPpOFtYZ6
e0CAVhaEvfqjjN4Z/0RdlsPVb7RC43f+HEIRwacW/QTxtIKIFMD0ZHKTaSp0DRz0JizodGJOv8ek
Xs1sb4/BSN8nK1L8wzbAfGHN9hEWDzA80wv1ArFafB+Uel7yeuZRQIG+S+AYklO0pUIx2TJjTSIV
exInppyvSc3sFgVUtCJwIfup0cxzaN0KF19obrvJka0lcxb6ss+voECfqDN9Ds6CTCoVu9mAX5wC
+oA4MvbpIowGP/JXiLS5NFOLZWQuJ5f7WAtNCXXFh7yJHSKptShrwBQXI4+DRZ2Bb4UjWIZgIXsM
298aoNn1eC+z7/OxcLnhufY0IOjnimjZ4wwgeRCN+099C/CmJHZp4ybT7oudfq2Pj2F9uRUi6oI0
wIK5Ssa06AQQCYy6uJvmHwMa1rnyY1HjMMoaTsPAXDu6eau9TTYmwOjzJO9MsMZKoKf+xebSasLq
Xh0IKLmmouJ7x7Z1YC3CrZp8JgXizpBhHb681DuJCGD7wcE/s3QWrpOHCiyjFnkdjzdnZNz+HE+O
e0dnJpN0q4H7sQGnX6XNd2hcSq1b2dbOKs06dxvKAwRFg3MKTnDMX0HhvPpAvdv+L1i75dl/T2ge
FL6LLv9uJykPzbSIHU2An3UPk3YI9AcztedW18SJzKOv1OKnjn5TBZIE+uUmlKzheG8ouWafrmQ5
0Ej7Klq/StAJaCFtQusXmXOUeGSm8dMdbJZ7py7KoU9oKs2ezbfvrZHFRb3ESHdT5TcMB+WblYML
SRgOBzXzjKdCOcToAzp0julBv34d7F7UWI0hP5VKqs3jy7SVs0MpqjU8OXMmRjitqTV2hFFbtq95
dWP1I2zEJG4/ug3x8q2Yc9gqQtLcvEnFNthYBEim++a4VnNpt8hrn5E8K8HxgRY5OZIyWQTkXFMP
OJb2neqNaED6jP1CseWFFPnZLXCdHTuXF6OEypRwKASdg19p8BbVjs2DhzQgvkwuB0mP23jY2OEy
CvZtxXri3+sKTRdMd/xc6k56TYJcPWcAITl25/Y/rci9hdlETioYlDVfIW8XVNs/2g3jrATMw1We
Qn1JHdlU0DXnZI7en0FBMZUFOQKJWW/XGhopKXsRJ9Mg66zLKzUI4M+BCJ4Ee702/ikFK0oXw9Az
LA8a1UH1k2VmiFDGxgZMewrjfk3z9jb4U+7udiTrtn/Fm0yd22zWVyaICl9QTHPteww5/P7HgPLD
4+fLHveY37pAx5vKeKSBW4nu4Iw2EEjB42alTY2MklRTDosxMWcGnChphasg/oLsyKur8/ppCCiw
kuLTr2SnFmrDs1arlaGT6n0lGNOijOyVPHLRrUTG4yF1kPdXxZEk61mXRSZrpF7rSOGqAKjmDt4F
uSXuryFP08Z10rQHSjBRYg6stU5OxHd2pt/qkKDJSSc25cr4doLOCgMiDy4aTKYAilipK8Mm6OmR
y4csRqcTj+bqA0AUoBqGABqFdNpgDK5wLLfSnUpSEc8PmT4Ty5pSojBU2lxHrXDw48jZao/tLIPj
C0FJscr+cRfVesvlTC4l3L/4zniHBWxdLWEZn3WuQMrly2VjsFEnunREusDan8IpgeW7dM8NJGlR
jinOFgGGaksRR2S8JSkB5QMoCL49aS2GBaG3C0stLEWwRBZ7QJnboc5QaHyv0TVIpJgjyQc+7GIG
Ox7rE2oHEscS1t/IGicEXwdn/BjOrFQHcfEO/viMmWFuUFuYPatvDIjuQYyMte7ldv/tl4dw5T5u
rcNAuQPETjh6RlmYOMn4RX2neBy9FXv6GIimfLS/0Tnpn6jj3B+yqhHfHNVxWQCqVDIQisxef+84
dW5w0/O4E1lu/jbItgBI2QfJP4w9FQH5h0MR2C0Mp94zmtwE0t+HKCBt2vJGF6sWO+iLUkwO5nrb
btHh5WaNbpQZgd7wtpH6KzoT0zuhCgLQQEOvdriAcEGXGk7F6JNitPNGGjn0ZcxyUqqRb+TJVL5q
x3pDVs6jGQ7GBT80Oirn49bwEg4KHCVxOoys7uA4zcyXQVgTJT+wTZ4wBhnYYRnnm1/PHQDfReup
MSd8QHo1C9shwHiMJnvxcD2KpBlmRiwTCWfto4YRPdQDNW7r5pv/SDyLUL8fL+Yw6VY49L6OA9Sd
vZ33OJvA6ACmfQoQZOmuojJ5Pvfn817AxBODmhfmaOTTjWW/WvaQj/aFShZ9FuB7CtVO68bAevTC
RGm0WseXNa28Cdaj94cW0/8dXAj1xLd/0Zj5CxZ5eoFhVfpWz0A4SxsKyHK4r0bl2OKgr3SfgQX9
iSrXCgzwXnE2ZhMgo5Wsn/B4KEMkkSrU2PlUdJwRKy1u7gGGcbCEfQLvAqn1bLAERrfgbnaCilJT
j+/v5Wi+YCSpn0IggMJPhit28XHZEGSBloS381Ins9++ml0xPduVLX4pnKYFwbaMCXeG+KuJ275Q
Dv1/RmU4ja+GnuGjjg4SN+47TkNixj7EelaNBb5J2EHlXH/aCTPwOk1F5fE7ydzrpbB0sCtbqqfj
SrNKfqf2xSFKOJ0cYeSTa05lomnvFnBDx/n9mIxpKlQcEVaIpfs/Q7Qyn2S0mphI1TBjkztAjK+z
FbahdLRw5Rj5mQeem9qOkX6AlDrziPhXfxKSRO57g2pd6urF/0mr+7i+XZULXpWxrFlO1xKihiol
9FhChJq7naX3IhwQsKiyIwIfK2hXz6BjxH/LTLMn50afJLSb40oiSWSVEyjdQ9oZWPikVqfuoqxT
g3BNERdQu9o4Y6Zi0mobtbmsYdAxXLhooMtnPJXT+c88fxmJWS1tP3V1Otn7fw8Lf8MWhuiRXmzl
zxRokvnen2fWULpRC3L3jAbO1luYjtrKIGyKmPi12g7bL9PYpXaVeK+bkaevje7D8E/XjC5jaiVL
yalECFnaLVhJqhCbTxUMJb5JMEzMYI5po7jzhCVFG3c1VJCOI7nd0rQuLu2YH48WoxLbBGPXPVo/
+gxjgzZ2l4AMuJi81g2y0CXdqO+bUWZcsqBhJLmhD5El7NpopMXAdHaR+/TJZMDiGtq/LsCsindm
fxZGOluFKu2i0a0GzOJWj6yA6XnTrvZBky8Sofsw1XHqoUC9yvlSyhcI+e5ddw79CNnwoDzUm8Zv
HpGtBiRDin7qovrog4FlRFQIc8a+MC7F3k8N5K66gIqKugWwy37B/6sR2o4M3wQGAA+6A5TdT2DH
vLq3OMkmJLkuJ8XIAj4XmG3KrvjY1gm/+mKqsp3KBPHbFPoyJ7ZozHGf13Uu+VbxWGkBumug9w6E
t1bQNC9yAKF8Z8PpmnE/dBq6ZfAKmEmLissBbwQo3oEO+WXApaCBnEKpAJma+fhgNUh2FEz0TaXH
NnUGy4pOQGpTNlCfJw/SY/jxCFvvZbAIrezl89b1DLU+pOl6oS5RvGHLCS0Hy4//YDRYNoGsVZnn
iLPCCDgZAIr+MuRQYaraSO8jMgq1bLK4JJ5NwbOznpgdURDp5uhdhDFnr/OfqySATFKVENBZjt3M
pqy51v9Ax8EgimfUhpJWOhgv49wx/3dLfKC+P1lolWveVhgKuxdNq3VZrqD6HzUBSxPkjgSCNUFB
hJIusSyEX/VTr1j2bbH6aqnPeJSm2y8cz2wROnEmTOTTrk3HIESmpcv8Rr/FHzhVPOEzgBPRSxJE
196t7GyGyBpFQz0UIfU4tNwfRvAD0ruy8apTs0dSpwX/4qDYvYCUKUQBysWkZvVAv80U6epINSQO
S8yICEXo/FiKAGoI8TgTpLTN5TUyZh1jDyD7FUT3Kh9t6p4Hh5U7DBAJDefSmhH5CrfRIwib1eMN
hzVg5exUtBWSSnIFaHASWAWF9uoG1u+Qg+IdUfWYpFQD5/7zlC+tDf3jOzXUbKlcnOpU7niJbFti
/SjKhCNU679XENGP4N+AnELQEdJWHOApFRh6b0QIFGQAyqXvazgHqaY5nBPcJgYoc0gbHB1pKFmj
mvsQVKHeGrMeP5EgxynNUzeAwIg6y+1br2nIfdqlsN1DfcsLgM/HHOnvmK0RvLPpGMQv2PAnnV4n
6jpzbkiY9Jvea9/lY9rORbJDsvC1FHodTDjyycREQRlbp7/qTwv9+oryiOi0zsRcujuQDPecw0xr
tHr6GCJLdd3IhhVhbBD6ULqfO8x6Q4TJb7H4ceLmVwTJnASpP+RxQhSsRMGNAsqbnwdiwg47teC+
vPtveyeHIoqdoR0KXg67zEWNR3uDurf/DWqsO1wmRaP5VlXeC63EUr7lvU7RTGBe+NLcShrq+nuR
JyskA7gH2uTUd/ijvcoRV/LJWIWqszfvjRPY4Iu+x8qEYuNEaFv4D3mMJJQr1/mpPNnshKSLaCYV
7qYHUiP6hBZuvfJWsysP11eZcFXWJv+x5Fe1TCS46x9LHnBJ0jVfIK9X8pXrsLcK91lTftKnaLgs
w3E8QiLZSjWAneet8RZl1aYpO2n6ia8UXSbLGH4SdeaHuyAJFsAnoaVIiUnEKcq87WZhPwnPyqwN
YJ/gVJgEej4JaMgcJRS8yennDFzqvwAbn3ISxHxlZJb+LSBGPMnB3nOqmUUiX2TXP/ZPwWtVYl3/
PYWPQCjj/uoFjK7aPNmVXeHKz8zy3lzfQGdpgXwQosbo6DQ3H5xeibje7l6u4PHyKJgu+tygSbAF
d6fo13NXuEjwA2g4eVFq3vmPgT4qPsbKCpFVGt3jOGax0KElIPeltY/AeAjrRD7dP5HkLZCme/cH
EMw974Ou7e9zCo4r3fpKwVdDCJsaBerDQcc/J1EbUWMLPd2jttPyqdtP9ZKOqlAgzJZ8Z3cEH+Ez
tS20ygGi7DaNApiq9EWw+Kd0iTG4ci8BHiyISlaUJbEGDXf0RSPE7Cz73dSiCkUARqVW9Tk2wQYu
YOE2oDV2NyLcg6ioglK1v3SfQVREo6QOpZRbP/z4DXo6q7PXQC1Gq6UhwfJazfMjfrnjO0x1CxJx
dwHkJ6WKGL4i1HdWnxgRpjXt49PcM94FZAP3FdeiVYxo04XmYzuukCc2SsdgMepo15ngYLzZE/kg
XW83M6W29Sv1yREghSnSNCB9XLmylUj4hjLOptQOJYg35tqeShUMENrcZiyoyl0o4hZqPoSPqjdG
QGlQh0ddqHwdrV7Z/whJnmtmV1Eypf7nAThFeeGyTJ5j4w8ffnccrAtd1rF69C4XFKWh2H4QePgW
LtEbV7wMsDoqVQIyNqzMYcgHM+4y4udQ/MdxF1IhzLRxHOB5OnEcwpJX7OHX3nS45lnKs+t5x/kr
s84yXOljmjn9C0h4NYdEYc2U6jL7+yqe8Kh8aSgtjdrJElA/xqOa5cSFkn0Cb/V4n8XXeliIMxkd
iDgQwMMMU24+4B/FgfF/53ULl2CtrqF8jPgPk9h9yDPCrmkOD+zN8o7NshnNhS7i46fuBGtXKHSm
x8BUAZb/dlnu9j8reWzp6p93ZETEnfQab83jsKO8d64qUWoMm3G7HqJv5aJFQSmiLbmwGSI3xf0A
djYD9WZ/7pzULjJMa0/lm7exa9ZaxdcU0T2Ufve9UXoIl75A5rpmlRSGKs6cZSy3UlBdhmuanhNp
XuXmv3WleZZXg2YxT316sJQtztULNr46KxzVopukJK1U3glNZRrIl/iVuEykwAqXfmH9A4mQkxsB
PqXQtyWHwWKwDOkE83/ufvEpjtpjraSakrgYij/bcccH+5VDiT7SDRIAr0PknvkaqhmhQYDZqym+
u4mtV0YbeCny+V/+aglpcr+jG5xNMH0XVrOWZIp9/VA3aGrWaiG/JIXJXz4r6x6QCSBrJ9Z19qaR
FrxYw1EcUW7lQfFpEWdaTMqX/zujqB8VMWOEDRAwWH0dS6YiySigquTkUr1On7SqmP7EVQDi5Ank
W7xGUrrPvg0bfse0viLAxh90rUDCiixuQkcv1iQq6WJCY39Wrhf97eaOKrK5nJyu8A5AclqsNVWR
uhaZnpU5Lg2B7midOZkVjAj4wLwJT4kKxM8zS45+0uUWvTONhkanjv3wm9AKDaR2BXBcgdKu4Z8D
jj73emSRD2MuWJAHQ6WcTe+S8AHzEw5plf6Je4V/LFQWAt5xH0gMigEtmGFP6wsOY1puJrLbmimj
Nest1qj7dSZCBzAvrCu92mY3tIhDjPXtOG3ujWDu7rcrxJwb/RzitG6D+i8c/SrIc+YGDFiR94z0
svqTSUWabtYWfMYtGvUWCQ/OrtnlPae/yMQLHTWkG1kov5K3WLw7bK+LgDQtIeb0hfKBPyYulCQr
nU+HESvm1bpt014z8uMBISFr2OYgNx6jtNvQ1Ess89Tegb/Asw8qZkwZ2SZe5QVVpQ6hAuxDZdHe
wRV6vX6DF5+bMZXVgtzOSZueCI5bqj1L13SI2chD+po1PejXFh9cbAbgLO1Bxx8Nofkzx0thNYzr
x8CIU/6uAbedSpksdRx38A674jzhFigNBV60z2ElDBayMtqNq082phc4JpdvIQT9c+jOhSMnna/4
wisMEMwBrpFIrILU2whKHkm9kEf+6lA7kcjabDOu89RkbgnvrdVZNh29aPifDSZO8Nz/fzk26AXT
POIlUw5n2vHjo7YpHX5ShQ5SMLXm7fJ0OC6BvyoG3EDhALhkZwV0ywlxucgRLb7s2ySYp8Bfg5g3
BK5RHQarS46gRvDjNt/1XduGyXgchTPSxDUjRQHOt+1+3gJqkqLYLIE+vQTDNH+4avN+PFY0CClz
8zz7vInftLFBSyY+OdHLEc3WanwBIIWGIOFzsLSQ8aP+ijBbZAimSBL4W8zAKwCirUnMCf8YESwM
ssaxdIDmK8K8FPbqmeuokwBXOU1EugGRNIkPIzldgFXGI6ANgDt+4PVW17WoS4iWaMtwgx7kIS1W
V0muG7g+Mz4huTHybAq7WUom0Hw5SI5U1YdVT9eA3fhysw5NT6wmap98YgSDpwyIgnIdN2awSXVp
3wCFAMBlYTjLcK9FECmUzP/ScZ/FpRVbObXz8zY6X8mBv0jeYfK8wKt2dbBiTx1rRiOD0E6CMlQB
s0b1pvyYe7yAVsMX42bWo1jj8hl9V6jixe3bUHNd2dh1ISZP6QqcT5Bl6hwTPO3+qrofXRNknYRt
z1FP6ujV6KIrDy7LwOCrijOeirWLYImJlA+Zgjdd/QWKdY6otdWfEe7gzlZZ2caII8PGFuJna4DR
msBeEd1wAkKJxc/PtSkYC516FnXh46Xy81PDblJZFQLRP6aWgPJyXsY4RzLgjvi+72FinFlU79mi
6nrPFAQc97Py0Porke8NIuk/Kae8n9LXQtpptJuYrofrdyLnSrOisMDhNUENhNMPnckYqOMSdiCI
57MJrmWevnJzMr0pPwjkeCwh9RWY1fJziGtxNxUyj2UmiutxbUJM8862XIZyAk83vERQhaFJlM5m
XkKFfPVWJ9xMHnOfGEldCZ69MyW3zp0jwNvlb2OWykkey763wnoMTxUpawB+e/Rylc+dJ+OSnjas
72cCxzT9p6aCLVZHukZoJY1XunDwPla2eAo3HvmlBGMhvZR5AgDSUPlmj7IIEwe01trantpKv52R
Bk5lZSfLs9mEDSmi+kfnjVJphBc3l9BCTQFT/kgAAS6sn6D1flIp8glG4lBYTDVNHpqomojqlWnr
DOVQoMOUsI4iUH7EyHGYJrLmGmYCI3zISUpGzsf0a7Nma8YIvDanZpePry74G/eAzEtgrh/kD/2e
vVV1ZtnI5BVtgqCMSFJ7uG0iNyLNf8Xa2cjGria9O7jprteVogTqwylWoVgMi5dwD+1kBJFmIoI2
u8+BqlXR3J3MjVSj0gs+Dvcx29TQa5ecB8bvQnVzq7266wFwLT4Mv3cPDSgkaze9gVoOKkz1cFp4
exALjjxrxWFDME570IBIUMZuusn2AV6BaJhc/4o39g195xzEkBkC0bmGN4W1GdLF91cFm/Ld9YK0
Te0Ntz11Cvux65w/alzwc7AmHgNRXc6ehBki2AAUtfiZ2NV6P8fNCtFmAZget5EwgyHOXVD59W/q
jMuW4omtCGpFZ6wu7VCahb/wiz7s6glEN3XdV5rgwLQmvk2t0+aLcIavU3kvmhv+2RiLvJaqrOHf
ynN+O/m0nNTJGUEuk60Co2K+GhsQSRExvP+cKMduBaceBPYbG9gVxFUTkWTqtw//VJAP3I/huXMH
u7JpLOUIZNZWDahXHxIgy63fUyiNUs1XRaY4qTBuS7Wy+BYdbc5gnh7Fl5eVlA070E2VlIxnf3e8
9bkhlD5sJ+jwg5btbmLw4RS/iVsEte9mWXx6yMZHlLtq7RBLfy7960s2A3aqFfJEHR8lASf0y9GU
yLwSaOBLKWmF3orvc5t8Bg3iuNu4M5Ke4s7AUnBs6vyoj4wKTn8ID7mv8Lq2i2aiWeyfub/2J6xf
OMd2s2hGFQIw7HyPth6rw3c/vr4tXKGfvi7tYlxyvaX8R55WUV9QV2CF2grbi/uKd/u9Atpt4PAz
R+Pk+bfYZsBFOawZputjU/JLBVI4xdkN2IOPeFsdfwVX84IgR7FyHSlZ/aKjG3K/kxCBfyRbWEmA
o2GKIARERK7PAlxcRSaVgTIHz9SveUJLKwmWKq7iTxm2psg4zHGC6C+y8/4i24Ens2F/a5kU0HJy
grmqfbNA0A+6VOxIug6foYqUlh55Hn40IyW2bkFNCabn9llijg5i+gOEqXDQJic4eUe4/rsTO+Lm
0HWEtQEFynKcH+HF9EhbIAJb3ptrYKdruy/ImtiIDChIbxGR23VHd0gmlhMAeChX4FdOGXBb5zhC
nouSVnYzoNNb0MnGJifgGeIWqRfBH6gKavanLirXuoFaIzU0gbg5/tvJjnT39DlbSv8+8nnOfNYj
+kgJzrAvA9eUplNJiCZwWenP/uvXglNjykJt6wYdCFZuc7jw9v9byyrUvEPKnnK864QRp29DqG7w
IzDPtjtS3MlTJ8aisp31Bwclx1lFLiWn5YbMvlC/6uIcmu32jTZceHhbNhRbMfnSs/gS0x4Y3WdK
QcYMt6Qz6Sj15XYWBThqBseHw17CuK13gvv+17o7/SifhJgurei/AG9RIBjfWZvZg5YMvBDPPr+H
ndYFp1KI8gTp/e9o5EdLPUYEIR/c7xziMro52Hpas8Qf90kM4b5poQzMu2ENhF38CtieNMd86MBO
I958DluvOkIiduT69HdUv36OC9lry5gpncoAK/ya68EL5iKwhkXcMQ3sxj4UGkPI5H+KGcZsg9aI
Q7zs4wlfZgOlNYCMxePxM/B0bpPCzLOi13WjI9KkH0+kyRCuN4xtOSVA+fN39BEc6NMMOteDf+xH
nw4VcA/ZdDrq5ycw7TN+sosxtgMdUCllF0rhMJKu4gagB/SS4onvSPmFTne9OJDoF9qp3GjmHoSc
VJyyZGzif6gJA/fvpG0fbihr++FvKGOL2DNmXj4KMzh1N4HqCdUmQy7a6mCN5jgJ9FzPyXB3bSKW
yKPfW1nZFxfxGnFqGtKFZLtTaRGzncT6LkipKdAZrvngmqh7+Jy5p6q1dXWokbo0rqT1m94UtIxL
rDxI6oAZJhbpYqdhqj7qgEwSJ1cFyiGh6weYSKkQ/uyR2O9S436+0xV4GaYiViY4j06XOY/49tM4
R5CKGpU+1A2QsBQpE8fsQnGbmVDOoX/cjSW7zLB26SFcpJPrxF15vYmdT3470A09tDR/ekt+85/A
jIXCPKh1MSdGd6wD/vE3v3rmkfuYqcPQV0Pk8+ca+PZ6uJOSzWBzND0bGtbDhdBPtzOLl6bEWIpK
VLU059mhESpW21f0faR57g5sA2w0z8Jushq/aWU6bzjgvuAnkSvGOd0h0v/m5oAMxo7PI1QAfG2b
tQTq9vhVRkXMPC+GW0Mj6WZpScn+tRNGpIxpxULuzKWCpR2NV6H2Sd9xYl5yo/KWCPc70ShjFyE4
xtMCV5rkof6anA3semZtYNM1lfisQ4wUFmpOfCukxylqSMhySNsPipsJQDaeNOAF1v2tgCtWHiw/
rA9UyJ7hYBwFhTV0mLn9sh0/G2/ZjJcVEt+WYP/N0Si791YSMXdtMiFLdtC9/lksu35XuIqgW4Ja
iNBOPsjAe/wsQJmbULizIJphd3DPSr5dV1Ht+cUOQ7L4MmkEHXNu3x0/irCUHXSZmErMxh6/LwYA
1mDoEcJMnk6BrL8iQvYMr1HcCppRCS7GhceT+mkIFKSgRr54r6FhRmBKj909ujh3OZAF0/8W15kg
jtsRgL44wkFfow8K8YKVpDb8H2zlTqa1ih6OI+wKQ5aelvYfkj2rIaCW9Nsjxt+AFUsK6uxYoL6i
/ncHhRDX0Bjqm9KgpsJtBMkmx0T72qGwWFUJNqcEpkkXgophLSBStIGUMxyl+f8+NNWwJFEJ5qPY
8iV3xxIPL6viyoqLt8VZoC32EQXcvDUW6TbSw7vk2mMAuLzd0DBdAAE6HOe93CsfeWeqvh2XjkJX
hSuPaxpk19q9EpQCerZBiMEAJ+2ZgGeKquaCK90Hemdw4dz00IU/nOo45AH2Fo0zc/YYXkxF+9sD
omKrjgezL6EhXKHsRUzyrOxWqcWj+bRUUsLgb/iNJB2z8lqP9hxOlAK6Usjc1AxQWlrIvJIWkxP7
sU2btKfxOy5s+5rc5TyKC22a4WqFCx/EWqZZMjfypJXE/cIL7smeDGWU5CmtnuSG9Fd8eKpBH4n7
9yp9dQU3eNnbnvqWYF2T0WbaHtq4UVGV5dUc0DT1C6wWqeQ2ckPX4FpKAMJMyw5XqZPn4hB61jEJ
Bm28Cpdh7AXEEDFE/YNAdaVzLoILwCt3zJ/eZG65wYXJYXbPcT99m9LVKOHAa/YYpr1rFDv1ZYaw
7Imo6G3hGvEuZs1qPgkAvtwXFejH/JcVkLfn5syeHc5/wviJf74gnNwkVKa+RX6c006UeyD17tTO
jhg3yOqgv2j1yKgXTZZnY33RkmRn02eCa57XhXAzap9KckAlddoIc63sCsoZfjGK6JSN99gYhXCj
BUZJ3MDCsvIuknImU/nqr2rrg1yjSI+mMVu3lghfAvLQnrj96EMM6QHQ5NvLS4x2LDVpkmGbUHvw
HQPK8e6t0MdhSxF8O0QypUElsi/Z+JQ5GvqTWdz34X0suJdfZ1K2nlOXlhxCxUnMvUiDr0T/m1iS
PYFPTfNRNtZOimYbjfp0I24HB8BcAbumnUJHGoWlapQT39fr1ty9RYpkKG7koWjzmecYI9MxRLNL
ZhEYFvjE8bvHRVLY4CANQRx/BhUZWB4Gtxmzt320HQ3fknxwm8jMX0A67UyffmxK92XMY146TwDH
wlsRI3/2UikBZHcQYgH1tFGcgvrj8+v0KxItYNuODtfFe9nYchaK6OMaqMx8wZ45a/Rgs+dd7u7q
6odO+z77Azn4OqfaLH2GHw71S55/nWzrS6mozH8rs7pYIe0gRjtDLg1QqvhbpcWOqXmsrGyFJSpA
u5ydP7pNxeHYmo0H4EiwBBzk1tfPgl+5iZ6E7WxVfqgPegfSCqIpvtznBoXx77arJVrH7JfM6mDx
SvcfkT6ymZ9x7WKtLRwzNMbosQ2hODPH/Fppc9oa+QXZzJtHvQduNnNuHbdtMEU2G/rLe5lYpJq2
4VTK8wKtp0dS7RAHQoS2A7uJlXe751Kp1pfRfjwzKC2rHjzfJ0qU/B/E628A7K7R+JvMhfiAlTor
/RmVLI4VBaxNdvoRxfgcrAV0LWp1jPrAfRn60cImRfMHIgmUSEtMTWhRagIKBtkK9t+pLR1K8nYb
LvnpiCzef3RQiTwQmfsLIpBt1+p9yxWlaSL9oOzc6Yxvoesq5b9PPsB5EJWsKRkalSy53XVi+Ugv
BJW1RaTg95OfG+CSYA0F4PdCmmf2NKFmY/NYC1lC06Q9IfdEMeGekvG2w2aKLOdja6mvzCLhVG6c
rzQsjnTrCIrDJYgHtJUSMR/ybyeTdaom+R1IPGehtMKfJ89/bCHgZiCPNYbKYvNRmFuMy8FSLywS
lBuq0pMxOwU5xcmBSz8am2DFNvjB6rHYGbDzJtpRfMDcMXM8wjOmzEg5iUelz07RA8/jTOrtgQb0
ttBbtHuDTOLJiHugcGV4RcC7m8Y49B3/yinxTJNcSH1NrnyNKqQsPlToUDRMEfUcKEk5U+peRZ/C
Ba6xrFPvFRGB3rbe8vpazQvyU0Vcls2tUpM+Q7UwgEmjWEvQyUkil/QYDQ951ShOzcPyUhPPkoyW
OVUenCTgyfbta9H+ETwFSrV/Yv5d75y0V1ETIIAAh2J7Wpa2I1/VB+gBEewbJ5UkGNFUXWsBbQor
iPLIa5ZNGiwjYZRpOaAp55q6BHjR6DzCAhm2utSdtANUakW9XdDlTUssfTdK7fjP2rsI+D1qz8r0
ZPTwk7EzIF+wilbgi4seDElHN0a5sXB7qswwx67cs9+UPpT6LGHv0BGjQhmiGQwVeG/EheJ4cwoR
efOGYC0Q7KIK3hc82RBDtQAW3HN9s7+AyWykhtUF8mBt5X2LFEWmFiM3bHqthDvrBNb1upvRSaGE
YG0h2vRxv6ytD/vJ968GF7/FztQwKAGa4VvcC5X0dYMuRVoFzqS/NmXUQ5mhSP00v9zKxaK6qYVS
w9z+ocNStRtVz+VOtAH5PQv/XgUzYulVyv+zH4eWAbEsv/5oQ8KZ2j6oWsiLF+WPEFp5hKWMGTjV
0aqhWHb/hZKfBR91uEnMmv6CVRmSLDe6CKykhS/AtnkzchP6lDpHSFdSr9YHrX5uZB4V8SmhJ15c
P4iGjlJuPMxY8JV0F8/Ry9odRaS2ZZGHUsW7c4E0OppwR8amFPyTa772P18PtyC/IbtLrdxwiR8w
KE8xZbFp3vpG9MWgZiBXHsG4kZMLv7axiqjQTLMcq9ZFktTIVjooMxndetTPXYn/k+PniohWXIxF
oohIzy93uYGb8a7hHmXnezaGxBn4EbmBT4xjNXptwapDTduaQZVAZFDROqMqS4MNX1Nta5MwLXRZ
TKvtAXaEs8QNjLJROO7i0BCwtPX53VgUThzZJlnR5aaAaf2+Ge9+BHuQVYgTkbl/lo+sghpRmmpT
z4EUF/9hj34TGTDRGXQiBy92VmW9ezBpQM5TW1h5EcotZzfR6SF51a/CODt1DHbQK8WXlCB8QVjZ
GO0qv/o92Vog9QS/nESMqALQnLWR+eC+Oc3MPDLJn8ealoZBgJaEnyqMBl7d/uQJdZEMIXhvxDyW
nYVtAGdDrZknwH4B5GlTVZdWpUljnfYtvM1LsrplAavgZNx2VbzqDu7N4idV9WXPw+gGHgC0KzgZ
/yReP29boFklhgOayeK6sAf2QHTQ9GiEY0P5n01LZdb7AMKOE5sSb5HYi2gttV2qvBVLe62i0UAD
UJgqNklQNfHvgVf8wPQueZLeLDBqQdjTHkrI8/l7ky5hwWFb5IMqdA5dkkIfObFqvwZ/yjAKlLvl
HbmK6bpNUPm5tLeR3k5/4Qf2nVEIM3eBZD8y0r5gnMz7mb1hL9YFY5er7Ld6Ll5TafRSYo9jrVz8
EOWD/fzUl8gDDqKNhbCz4vAqZBNd3DiCpE3RhVW7oYjWmLEy5hGP5ucLVDdCrik/BV5ko0sDE6Od
kH3v+wXEH8xNUwogD7xc+Iri0XMHuGx2ViwitL1BKulewMsLLHJM1Wp7CmmRn3nSO12qFnW8htfk
V8nPmnj26E7MU9NY6lnY6IPKAaUsX95x7X8S1V2I7xRFO81aK/oWbRcZ2iCqV5nN6tB3HZQV9PhL
zzH3NaFX/lJcM+RSAZSskNnmQ5BV4qIdOYaLgPard+EBeuo2RBqpOlgIG3kV2UDADUBP94GoGKLA
mhrbpQHNdVaRZBEX/us++ZozILdO50yAaH/KK4sJD3q5dG6UD4rGDf3A+8i1sEd44zAmQ/bCZW/A
f/eB1hYXqhgToqmuW8gM644IHkqPzrvyXUiM2fpBu31cJRYKlOP0HUJSwaojzq7NAVTUwHGXPYSp
ya1LsAl1XCQnUQO+2YuSgXoSdh4wVuf5BlWclRselN9HReDjR2FymSXBqVBcwOTueT1eH3xclvLU
/2hqbnrhSQU65R2RlkClOgV2bW85mnoUma3Mo1b0HCHfSq5DUSDzpUWg+zdWFmCFkMgmv2g9z6Um
vl/JpFChUOoXMYgTFvt0Id9HH7rQ0U0r8v9v6VlDCWW1g6oR2da+u8WxtUEDaN/b9Ftbx+I/i1N/
EoJgpa59fDMhafkGD78wFytw3FU9ukD7ao6tP810DYAHNa1xtYjb7eyrpVQwmjVmPtDc8Oce4qiC
l+1OXDRni2U5YeepKkBDw28N44A7WcQnI1NyKAWZLK1QCjUNM62SO02I8Mu+hvRhyCr98QSpa5nx
ruqLrRRhZ5byc6v54v76GsvuWFVfu/C65VqUueKyh5dyZNRqu+HI0WSqBLfHC1m6+NTlxlFgFkGT
gdbRynIZizDudVkyqC5GbxmlHR/IObPyZkzrGTlyJKt2rrKu/M7W2pCYwLQyrei4Datl5aNTwM3X
n91+5H1Xe3OSmFElvI7ERu1aY6hybTre9jbqhlr7V7MZlMxnCXbtq96ktRGFo4jvTDQp2CcAancb
z8KOhCnh9E2nWU7HR4UlIfNObNAy5epBjkMB5p6p3fuYLVV1ncPfo6LxDsr+et984u7qzG1TaEHN
upRrllMI0wch9Sdh1swHWQ7Q6+ueTfP+N2CTaamfU+xAlUY9A8UiBmM4HppLy3dlxxqJRaNPdg5i
Psw5+92yULrk31qEznbLPz1eqiSprYu8GtCO0BmbSzBKEGNQqSD9D+9hQiUATa4UEFS+K7oFONE+
JZCgfDo6pBHkRWlBJl18xcxDKBjl3WV84Cu6Sm1of+PzKuJ4pk82xppaWooJszy6xCTa1cjc8wuv
Acz3UBm8qc9qMr1Nu/dsIjbNpTXUZr9bGX2j1bVpgPEmQyOcTYebL1BWEDSWZkNeLH0rANVGJgkW
hKK8aVXrO2Y/ujxQ9rWWIz8j36oStdIz9E+PKYbrcn6JcJwA1q4X1vzhBWoP2Rba3aBYusiXrA0L
XtHS7llmaO3kb82D9GohuLD4hAtdJvVRwmHtizXHItK0893TpsiHgMNqAbcmLpKxlaSgOs3JPana
4UNCi9MA2wk2MbzL74gTg8yTgxdKRbhjeATSk96R9/z8zRr8y63kKmsnZp0GnYcVBZkw2HEYrbZT
x/h+uBkF0Ugle1DMzhflSnd2Y/GC/uGAim/2mp738nJnmJ4OZeo2AWd/d/ESXk+cjKP6IAiWyAQw
k03Oro7xDPL48Nn2QmeFQx+iC7dxtq8pFDZvCjMf5ZDq0IQH5hnggo6coGtTbKgXFCy0J5ND3vLP
m+m0yOTRrSu/zYBfcRnRHpxZj9HQMKxfTDy4W+F4IszZikX618MDdaFMLsmKqWZp2xgR9nmio8Wu
W3GitUfFEWb9wV53G3gr7B+KUxVq8YVH8azT7/xNVg/B1JJAyNFZT+eVbJbNKppMadFlpziksADU
A1t+l1X1ZEYgtA064ifNyQVcIS5zV3it2wUJhkuVVM8O5LuYR88oJjqJeN18ub/ndJ3y0fXI+jNb
XGAo+Ucse+L4TxeNb/11OGKKoPUMVyDN0fLRAGtCgArHMLF07PRdrgJwohuaiBmNn8fN8OR7gILm
MyW+KHXlYjSIX2Pyc044CRCuEW19vnw+FnhG5DQqYOO3SX78atbLlJbQyk8sCQ6ct6yiwIhTiRs4
pyT5MtOvRm1MIgzajI2dmWJbGHsaIab9T9YxTklYTxAvSmohc27z0XNkAs6LjdpRXHK5apXgthK5
AEFlDBGRLjou5jqELISH3bxAM5d8HuxDtmg9eUwUZLDiT4sxZrGNL2Pv22q6+uNdfslhq9ExrnDy
RaCDvKLUswuAmfUtqztTthtkwViH+ZyyO5/Y3FwQipUt+vVRLCcuCfQN0JAVZAD2FFpoMkZXsozP
dr9kY4471Jh6sP4LeMtkCv4e7YSKS8OZnkqj8I6HoPeVjc0shi6W8QrFa7uYANoT8hJSnkg3RxGm
zVja/xMscoKIVSNd3fQDYLaElT4y4ZPMHSTf2a9QncN7yFukxBJaddsGdFmi5jpqGs/REqZCWSoS
hLgSY0QBHI7V3TslbdimGQgPxZ4zw68F3Umcg/T6Xuqobn5emhED5eeqWxaq+zLRNqZka+jkQ1nU
P2X3K8l99Lk2nzSrBpfZMOcJbKqcukdf4qil6N0KXklsXroHiBx5dkpiutJ4tlyeA3lAJ03baCLO
CNm6zZnRJLwssX0bXXJp2wE8mqcsjQj2NV95g0D2OTMCQkhMvAVirzHFILSNG6ypoPh9JMtVI6hE
462Ap5JbwR3mimljrhP07g0H2RWjG/qQJnSbwDHpo1MZ/Ozj1ItkDkuSwXxi3N8M9JWlxzl8C86e
FjRNcKe+Y89Y63wMZhCJLYqqgJuwPajLO2AfqGFO8qgvOGHP/i9fmHM9UGFC3B7M2XcFo4urojkl
KpggVOeozCNCtG7h9OddOyumxtr2qUq29+huLv5jJ5cH3zyBA+Rz82p+ztbcAS3wxpBUY0sDEzRv
A2yWd6wrASdkGj4WstybRBD8S70s7c9Mx4bfMe1QihQw55De+4+zmyk65HTz0pSAYc3i/RKWO+Y9
53/l9LfjWVwKY0RKEpBxQnd3DkEEJ1H+AznZV7TSTAHYAkEQkGR6VSANY72Gbgjjbr9zj2JQSuRy
VNnJAT4g1dMGNScs94FY8+Pkm7bAMmElvoVsnzbzZsWEML9qRaAwyAQNOF7gwrQKYKkYarZd+Hrf
PreAPbOwo2I+2cja/RmqQNcgY7/XZe4BzrcJOPzMdxVqI289RUkWs/iY66Gi2ucLM/2H1j+Ur8ky
+J2oh6uV+LxbAdoK30E5DvSQsH5nmfGnxry+d+wZuG5e2KYC1VuwtS0rPmN3dDqWjnxNiqQGbKXC
dHijP7Oe47PZAngoY7FF4U4CWHQcNCW8rlAv7HWkXriLlTP3Zx8cjzGhyCH7JoGYHR8yYSSLgseM
uL3AeIy88S5z0yJRMkglVojyctFc9khhRhexpC0Q9bRZx8D3QsGkHOisfLmZpmLOzC81137hnDtM
4gKHQbHZk3G/QsNcm+gXvoVeCGGUDIhaZGXH5f8vOp+7T5iNaiHcI+DkO+/DzLTJGepMVj5APB8S
Hn6N4BBgXahvXVYc6qxJEFXqcR5HOBXXKGwty16etMSHXb17q6TCCqcRC2ELsQQwM8RtEd45B3cE
W8fKtYSnMV9lv+50nrlEEhodJzbDD2psG/geUZu6ZqiCn1opdMXdPGnDmsoTeNPe8VRzOn6SFwPP
SE4HOvzQr4cMbdUJJ1Na4vWbfsPPrGRWy3yx0bt8cGNlGMdKTr4XHOAKALjedlsdO4GtI5pf9ZHM
YdskR9frud+4cQOr8bnmCFKYpTm2A7YdrcvZCsHdYEW9jLCiIdIjyptNgt+bqNyzjtfjRiBbnf07
xD3vQxFFvx4/4j2Wg/isCPf3hS9MEdCuQ7uBXrJjWksq6LNeU3if7zcgbQBIHaHKilU4Mao35eqq
Q0opgukJj8pg8EHjFnoiOaXZbxG11QhFwJekIkfgRKCFy7fyEeAknehP2keBaUKBI26X6NM/Uovw
L1c7d7/rzFnclrgBGobzvCGuacS6EinHHwI7690C5Oxz/xTnOn0fmQ3588wMzoOYh8kxpEPYZBYP
VV5COHLXZL8W8ETH7S0DRvfvuGeJrs0qCtCBoNL2KdZqccr5hzM4XLd1UBF+PhZDyYByt1k9Iy89
GrkDTOfJm+YS6cvpl+oEX4TMkHyfvADB2v9zPN/0hLKJ1AFGaSYVM+uSGhckqImSjpMy9bRGbW/U
7l0nDS9HdO+L3VgXbZCYcgRGI4K6fxcYj0RiTBitl0y+NsIOKjDWXjVfPgTzj+XXI2KgGis9dVUs
7oteWnQXpd2JTx8QLc0qtcPSkeafgUAfSjL0YlosZ5hCxb/wtZQVS4PHGAasZqcybQOUtn7FnLDF
8VTjO7bumvpIydG9t9/BIRiLPyfJ1+ekcRxVvSzpzawYwYCTSrhgTmkGoC+IZxicXoYSWMQ2kY0r
hkkSkc9pqInSaqr4jMH2ViomSyk4i/NFlaf1GGjAJ/mnXVBsQO7TMNhVDGqFAVepoU1ps18mJ5g0
NQ08DSWRzNnZ0ukvUT+WfLfZzbDLw+m5H44zEG3iNszEq55eGM0qKRSd5sk8HR3E5F9nFk3xKyg4
qy0FqeyynIPCPEMNsV4+ctwMcNX9nxB7R92OPDFjZN16VkzGd9oW3DXbdY828/Jp2CN6L7o3c++B
NuVUFadXJ3YGunMq4rSk7kiB5m04tx1QOYOTiwugCmlSNtAWS0j8R3JmIA9XMXOGJC24HsqulwQz
oY0EaWY/p0RjPdSwDpov8RvuUYh/LOKxmtbRlmBMYlVau5CmYlJNo0PDX942y7Y94ZbScqSAP8tl
830KZ5owfPCrFO+LcbX27zgmT/fwkXvK9WG/vQ5NbKS1o6t+3TovbozUSIwaXC6c376Q/7VJPKJQ
FLmuorZhg9sc9TFguHfOFy4V5+3kT1FbzPkYQ+n/V8ink8OddKYftraBeWX4pRXo6NVrN05OzgeP
2WTMYf6eIc2hyO+h4a8MlA5HBqrWsDIMb3hyY/cfEeUY0PPVJGOz1vhCG4GstMddikHfNMYZTRBh
flfs27d5/OmPecV8GxMEeANkGeF09mx+a/79uVznU+vLXoqAvyMK2HgBoy/yY0V6K0WF/49g3xNX
Qc2oVZrRSK6SM8xhsUerBJ7Y3RuGFu0kOdGImqyThLX6s0IzIJtFFRrVRbx7oPMffTEU9yidPbG7
Lwa6SzixZr6AviVN8SHKwVNIZRprc0s+AIg9vkHPGoL5M95AWdI5EOISkmBBiLChbPmRwWnQgue8
gfZgpMAyXZT1I77fs7wENs71nGwocildIh85ZNk29IKwVj0PEuHLv00/yvK33xiY7zL32Jn2/LuQ
l94SMqeyoZj2Sbk0BstOmjmS6Hw6rSV5YMtVTUwfop9W7HU1tTZsvGM5ovirwfP4h6H0txt3709B
BVDf+VnKgl4NSWydas6yBFi+MauKbEDUb7pylt6sgMzOxA1s9K6X1vfBFXRId+16H1hsKuTGZbwV
Pe+w2wc7tzzrAm2dVNVvknRDKXHX+M6xymd1OW5rgXUVEzdWA8LaDHGVp8RpiFUfNnQtVAkbnQO5
kN/EMxHuqb/gzuypTqc+S6NGCHi2+9N1ia0znD6nmDq16BVhC8xsXcGWxtYnxszOTbJZsPSw1iGl
7p2+UKft50zYeU33xP6GEcVUfvZdhszaT3Nt47RaeyOb0iRDG5b+ez86AXQpGQf/dGqMOX8wF8j0
iSyACuPhGnEnHtY0IC1PPAxj+FGqmjrLyhwDCgNxoKtJrM0Ekd7TZrqRoFIrRS0Vg6AX4Pl0OwKW
hUk0VILy3rFzjB8mhZOxhBo2m3puA4HwlbwDpjpUZ8858YPhGTuKjGVZPOOlGNvPhjtXDh/p45dU
ziIbs30NF4NWQotoxJJoXtT/eXswqlmlb596woedWT4kjOBTnkMHTzLEzbs2qBOemYPZxCbTRjzT
sZF0PMg/YCCaq5HwAl6V4uOfPuGx3BOGmlbOy5Gw5rTrDVKdt3qYec2rlkT+iR6nhec6gxnM6tFe
DS+6yGrRdF57nonUcej122FPCtUZLT6NBOjXnVv4zZjjHODtu6aXedEdfgIV1T61Y7mHFoOsbugP
7nodRBq5nrh6ZGj2erKApGMYOjxXEq+9O3G4LeEe9vlj0bNokD5597yvbc7SN1x+l/sApMYEXxPG
q7obbdEFI51V1NxgYckT1L4e+Ji5DoTwZ9PyAnJ15kgrCvucwkAETl19rcE6yiujMRJGT/vXQlW5
GKHUvKvqnuD10kTbtO83myJz3xkcSLlxcbi8J35KehGbACabWkUhRC1PNQ8oojhF2MOi1Bhyv/wr
/eleuNzD9KSvDU7YPXMJE6AbBapayyGFTceUUsOU1xYkU3k/2NGv0p+u28BB7gKopT02fY9NUb50
Yjk437ndb6TpmzW9Bul0h15LPT4X9KwX1sCFLI6U9ynBYhuJO1EXE7AJT+XWkgQbsJbrnlD28kB/
c7g5tfFk5VRJEntLcPkDkBrI5e8hNMKBQ7J22fgttzjzI7QKndMGnyodbLNsOZBECZZYY8OBXqL1
AdVUVr8XX16bCRx/BNSYejh7XndNaL61efJqXN3mW5PkyQzh+C9MQo7V34oa2sQyPIKBSAcyLxMa
oKuJXzYjAWhyq3c23TxtWixPlznIHuTnme5tZoGtujGiZBst3dXJkCSu1QcBo1/r2DGlV2eXyRVn
k1oNV1Xfx/JpX/uphrQXr8Yqr2L4Bop5VgufD7GJskH9JIpzu9M7WpoRhzUIRmhs1uYuu3XGxrRV
8OUKzCCtXYvbbdLv2y2oUwB7Ch++ttTQLh70l/4E1irqw/sMrgRTpfa6diQxOrEqf2VGloM9Qa3r
ZAoiw5yFHHumAyuEoZAwwC9L0Bh84UaaMdIN9VI3OKdcdb9V61Jugen38GgeBNzIrH2fQ+RR9sLJ
dcmkTipz7X55GfQ1EHpGgZeZV90ffUtndCkz2HkvS9neoUxHyeuEV6V2/BAupG9t0wY8RmpwU+E+
zR4aXHUg6/WJUfs1enc1baHtdqOIJWLveF/UTlLOa0vMjtfXIl450sjIAu4Vxsdbkkke2xpef7OZ
UVhhrRavs8n2fxSbB5x5IPDI0TqXAXwBPJWj7lArIAjqkjha+zQWQfiujmUToPaXMsE+6Hn3lIoZ
pV/9rZJestDrpwhY5VJT/cAiZluMJ0a+vLtFFXaw0nTJuKUa60PCYPuFFmvwjDxE5T0ENZnW0mHY
cb3n9sq5AM3aBpnX9/5yODkZaby0rphJsGMFgSDW8Vm12bAQwRce7j43LIF4hbb6kJNoc7l/WdRw
U2u38KGyQTOysS2SyrkaTX9DrhwNwnjF5C7ipPBgMaz+lrWHU9/Z15KXgykkxEnngSei7JLIDrjD
aYufOKlQRAM9MGJCUK1sg3D3HjvEvRjDkNOsJJg3dkmxfviEdhWyxxVeqL6tvHYhbMwrIVi/XjFN
uK6fnt3kkKxdNuzRFdR6GhC/NJdETecqtiQ7ioaxTHRAUICKScka7Qqo47TrnBO+FASa81Ozg+yG
LHxLb6lj7qGAld4EG0x48V53f4ZJslJKakFmU3+27yRl3adyAr5wlqs92vjOcj03UBbFCXpl44pf
jqmtJKQ3WmERXm0fjxRLGQPlnpBPdN9WCZ2ebimSkdIcK10uKOdV4Q6HyjJkDaXm/Hs4Exb/nLob
lN5btsxO2MxMghyzsCFxVvK4tOe+1YSyGD7CO4taUjwtjrfG+GmtuhgAon7ikesQYgHr4QlLlnwB
sg1qpzkqEqDet+eYcxuVeqJg2CF5Q6N5RWw1lRjZasDTkB357k6IMkrwlhfeFVkfADsl8hvQ/f4X
UA4fkJ9FHsTCqcCt8FO4wfOlTkX+sv7M0lho0dZcUznhF+z68diLLIkWNY8RCxkqOmi4otY6oyss
rsrB6q57Bju57IvCRAOzPaD7qscZ2w5K7ztr/ckIFcHwbBlQp9pyFZ37H9lWmxCfITirA20MA8S2
dn56NAnfASFTmgYYUevzpLC4V2Jq/GfKy75kKEfUOwkWNQnn47StHNM1dN15PJ0oIBS5IcIhpOws
zCxo/j4xqNJ3VKe0me/FdfIttgLLZDXQqqdiKt9CkaFGvZ3vjseSy1dB1asvY2j5u/rmpSBcTytW
qSPd6Bj2w1W2YAWp/FLLSwsGusWN1PBmdMV3eFyW/xd2MHn2yHNcPZFZMJpy1bfShZvkxqrl01/0
AlDeLco87oh205ae+jsqJDjljyXyHVpFJBtcXA/TUrAV9nfpeci8L80ug406SlavgfGeBfLgPCB9
WEuntssias1w8IDbtUlwS8/GxpNRO2LJulWfgBY2mxGtJ96FAAA3QrFB6zOJ1KwAT9gzbYYS1Bru
48GX9i7hsQu7ygBm0pseQktifcbEUS/nhD2h6avtYk+cBddm/LjWEofZzr8OV1z6AuWsRRlzHZCA
2TxKV9bobYWeQ98tuBqJT2jW7bpP/lcZ0xBmwjaZcDjNKfEJX5B0tzZjKdQvmLV0t2zdlrpzOxMR
cZifOMhCTjGWIuN8DftSn0LXou2ysNkAYdheVuayHJoAZby71jlv9lV0FQBoh5skTL6Ns/FuLMeH
W4TfEJapjfVhIvRL/qV3/pBlXk0ebD2FgvMxSo6cJZ6OuDVsHvZnluCU7HqR4Zj81onR3gQQ8VIO
pJWZ4pZyuKZwAryjuzxerDtj2iaLrJLa3VIHGMjBVVhLdYw1TrFqAbttiG+dutEUSx8I5cwcR3dG
Jtv+SBPNUJlUYv2rNCyOgIhyuKWjp+gvYTfZ1LjNIBO5v0lkNdxRB0iHkXVZ6d6yvkvYPOxc4TiH
jEvl1vPKcNDJkfwNdEg0wB509cNr+oEc227uyxWK7VSQ+JHCqFPkq8SBsxzCys6Ezk1j3a286yDQ
85zFy5hm9aqY6yQPiHVz2yDkYIZ36U3x2cOxGsr3n4knMCw7FkA/AE6GVy82CZeUF6e6uODmRG8N
tR+Zz8Cu+BMFUrDrOvFCjZN/GhaKj5dA9YDAts6ndBfmuDMdXf4zk3Z9XfanRG0dPM17hHG5FjPb
3PmuPEjRVCFbCLqmyN3gZo7ircyaMFVQ/Mo8P6P0zbyqP1vMcdD8szH/+Jd9L+DgZFr4cVhOoXG6
B1KPpuUwMBnuf/wCXGrs9cChJQZSbbDJWTY1IS+Gorflnl9IQ2EUNhQKYfE9vgANJmSJRmjGIKFG
mqSuZYez6Ns3jp5TsHEJEofNurGRg8T61RxZFNWw2U+YVxuhJrkvpCJ56iYVl+nCz4dLA6svLUwU
T9uPhWodFf8/u4iY6v+qOGH9gjH7wRms9p8pS42RN3KzbPFAt2DY2PzuDbfHdsraMEkeoz3xGeBQ
WqFZboTBid2G2H7+/j4su0PSs7+ySz8Pi5cMHarX8XbZRXkOIa9ZJxAXoOlQQLHsEqlZfaYTKifp
Q5NFBRjwtMVRg+0Zj5WQ0TpTC5+rVA7hku30vjsi65eLsA50k45Mlikuccul36vQUdPa4nZQ5hk/
itJelCLyykcC5e5CE6XcUYxKIth6i1kgv1WEqm5fa7cyhekv7PcHAOJ6ggx0E7gnlv8eznjX1cZk
zQwmPcCNyNr3hs1uzEVr5hCOYGblUCBQzej09p80aV6U110HqVOjaY+9bHUsskMAcW07xu+0EYlP
WtlwJxvFNVCPc8HuK7G/MowJDi6lkhM47CcVi34lln4fPqTIOfDLhjKmUULOyTiHyjxPf60ytIH2
wSODZfTPMsoeSiuGxn/uVbviIu+cZ/Vx5jhsf4Yaw+MXAQK/Rgo+j0ZVAaMZwk6H1lOgPdRLTu0H
LQrpvfgLvNp7iqqnLj6r7Ms4no4++HgP/PH7+812o5/CRAUxowu+7Z7WK4lvdLAKHM0nWbI/G/ds
8TKzU2JJjV2XcaSq67n00za4gSEY2WC9itBp05AGEfQF56SI7IntozmxywRlxAwnO7jzy/SJJJl8
FmyaYCyV9ghLqJ8K/FNfvDXZYDo2uXUbN1OwKPGakjBxWAyHNqRc9jg9osCqxSIA4Hzy/JbmRpSu
GOeEuJG4lhm/l3z74lRSv9/HX5rW+jRt89bjayKkNYyFtmHRNhshHf47QtQbzwDGu7a538LndrR5
HRWk305UuWLIBuNmPcSp50zBJ0K0Lw38R9u1NEc3Ymig87YvbMlsgrBKIpJWk+8SEYQh+WV1Zjln
a12eV21EMJbAuTQBkWlElbBNHXSljhTuhSOtm/KoOd/rxenifHt4AvdLb1jgS2SHHg5rkT10VJRY
/e0FTPTbrwG1XNNrP5YG/EmFN6PGREfxXCBAQjO1/6YUpeZG3zLB7KlhrT4vuDtVn/3Xs1bFcr/A
9H6M5mpdh7mAWw46yNeWK9IswFiMh6ydwfw84rSTqx78n1Scm3+TDZvwnvlaoYNevP/PLF1S1Gml
NdCeEV5O8q86MRSMZjff549dyAtUIosWsPFA/N/+RibPhw3ghM82XrvKB4xcCxNbMfWQNt+Y+qeb
VIhwlvokqAwUkpLcG4WnZM0NK3gzwMcY2DqO2Ay7x9dH/INV7VWrbbGXcLbd17Uma06JHkIjhbUF
EHN9iIrZuA1YTZ9iefzMN1MGu+2gOpw/rbPXioR+UrVRqVAm/cub8+HACxfw5lDivO6I15VjSRNf
HJcg1e2ReKVcaz4KoKh80qG1V49CR/OBGDbX3u9HlNdO0vrASjc8m9rFif8MwpMIwuiEx561u+r7
KeFtfXJW4tz8jEEc4VjyHlP0pJtdsRGkQ5d9KPLCFHWWNh5yyvgXudG6oVIxJav2xwi/NByt9787
FMDKrh9YQo872ptinLPMDW2JSi6U08YegsHR3v+CwwILzSpDKhsrJkIG93tP7fCpi3qW7ZiTCAB4
+sYxywDRFxQalExPcRtmDZPLkmGb7sxF+CV1DK44Cd8NIQLvB1v0rpukv4JbMyCYmLHV3mclonht
ZrsiOcZbTpv36p6PomgzKJTMV83mJOmvz5Zk24qEXkbBFD/Qu/d+G0AuxnnaFpWiye0UTPmYBFMS
pOXc+ban7v36J96jjvFskUvD9N0OEfXvsdLzooax9BMt1NQ6aXMQDByVeRC+q534ynL4baHNPpEg
kMVI3UD5Q2fA4RMPgF3LYsagKSeA3vRjkVvPVr5AsMR2lyn3IuGwuLmiVIqItupGpx8fV1CdnFkV
9vuj4ivDSNz3sQJICMLL2zcgRf2unpMieEC1e03/mPZtNF+/Fa5kXC3NJ+1xhOyDm4NC1LzSlm3H
m+qXACaQ2J8E7frviXsRmU+wZLhSrZkhstiKfy2WTMqfa/FRvlvzhPAJQ0JVxC3PEYLp4tI4woZc
95LLNH+yIlvPAiounMuWXhagY0N59W66mSgMxLKSAG4HqxQR0fPptQThpotsUDcQ78y5kOj5Vk3L
fpiZVZRM+UcCxowAjAMvLR2+cbRQtMpDLOZommNcMzoKg/1P7yhanB161LjFiRtyAYfzibMEDClK
WfWBMKhPO4V+qlC8AkbU+CWBXxtVJil75TjthCLHGY1HB8lLKjXAbJcSOKAQIC3MMfX7m5I85yPE
vB3zFe9FaBWwBLJ60odloOC4sczYmysz/k37EY1iIotKynSf/t3aVVQsbFUMBoO4rbQjBIxfgcUJ
Px5FI6WQoxQS2MJ1EHHOVynX51o682Xr/r0jcvTIGZTwxsfD51SVQGOW4dRlgnsg4I+9T2V7Y6WU
e8TUvUsuXFjnKnuDx3hKw3pi72ZJKJ241x1ERapSmhTlik6DlZYGHHlbOcCHLESjjYWoWaCpst2V
40ertFmV7pRY7sg+RiNNYpvB759yr4vgouvpfbTAiC40gVNDNy+gTePBJHCfTqibcFgniGoGxiqE
H/QH4mr0GCaTno514qipdQGFJYt800Vg9m4IAq0nMAQJB/BDivGcddNyETE3N386CdpDQrVbrox/
+Oku/iSVzybQVw4r5TH5V+HgIs4jxF2RHFiTwHZZ68EQ/n1OmCMJ5A95K9S0ZejQoYgZ5d5mjoPM
cFLHf1O2aWM9EpYcBiULtOSxvbtkWxceQRZ8q0WV4BER3wFS9jaSqNaonVpTZ6hp4sl4Su4Ll7S0
Zi8GFY/WMViW4hoNcq4RqKAb+9y9N6AV6kegaJpZotcoVoRksZiD5ZV27bA1mKJ5co7RC1q63tB9
URAS88fJcTUq+DuwsRnL7qBa3POGvedj4CuthDJUohfDTJbqsnHXGvA6ZwP1JWuwzqSzkI6DKJD5
oeAcXZ4AOZSEVzUpHjHPsBRzwhzs/PYQZhkIfxMzj/6PLt/1V7Vtvlp2j24Aco85ATW21sh9ShTr
Ve0EKcxVLhhtmgc2oYQvmDplF4SyJ9WgFDkN8ls2jU7ayUyQ4LgNg58L1BItXc2pSLumXoGRhHfV
oYPe5vBNEiQIS66Fn9TPGZVihCmBYT9SujJt4SyDYex13gO648h4rPngvEjlw/NivZcFbzTK3lhm
UakDWFi4qd2AMkyrqP7bnxFdr/RaZf4Ovt5XVMGSYyuo1IaUNhS3Gu34kDu68ZhJzyaUPYfII8p0
ugZ20G2xCr4NwmiH58uhCYjF6tbHCqmJgnU7sD4DyTdXwGw5JNDdixJh1i88wAyXTEY0d2HnbYU4
L4fg+BkWY+5cdwSlZRrBDGDNpDil88cru/4HmSIAcLj+R1cGTM4g7OlZG7R5JeYqJEvxrK5175nw
Rzv+X1NBNYRPhh7h+MTgv4Tmw/OifmRpqc24GYRYWc3darxy9XGnLxgwpZgqVYrRK8nh5HJ7pZTk
ESV8yNWM7gqgtJ2k8gScy66lEthTttiJfqlRmlr+pRjALT+7q6JsPh6nHMgXVWpK+Y6qKrnwlYf5
8+JyPRSE0YqckiItJv5/HRmWC9QChlxcoymGnudZjYlZxPgD9jASdZeaXYZOHB75N/aq7iWmGlx6
zX0Jo9coarRqo3ETrF6y2CxBUs5yfr7OjTFnpNJ/+gJpSrfh+kR9WllWhl7nxJ2CgnbU82n0fxpu
jYzj29BBQRx/BPQTGJapRnFWP3Vs50bbL8X5ERPDZlXiXfwVuNWw21wRmq9cQnk/22ridow+NP7O
sVU5W+GYVPMwZHyaz1uiCR0XHltBURlr2Vav8Vx9oRufUQm5CvjjhNpfyRZWJ7jYv+FLjuAcnUet
AsLoQIMWTg5mJfInUOTuKq3swzv1IJPKhC/8pO4KfHH3HeUxZA6BkCknvwVU2WoPkWbZiapbE3Yd
sPjEGNfnXWfxZ4tSUomcaA5823EFUvcKSEFl57rcNQxRFtIiA0bvAJ2w0ZWPw9Ae9nwXw8rh6H+3
EcuTlREMb125H0O2gLlhedn4gpdDvbYXx4YLn7z8UwnYC8Yxq6wq2bDqRgm3V411ihebPHwO/V3m
jjkEUBNfxJpjVNOBK0mecLL6qq7hzrf6I/IL4avliLR8nRCcJZ5+vqbUOXjSA0PjzpqL5Pg2Lc0V
tHwQbeQX0vYJHThmIpZEoI3Nz8jiSIy6Udyo6AwCyzA/eH8FOLXV7TbpMPrOE8zuARSRUVmFbL0r
Gq9GQa0y9uUslNHAFBZKj/dGOib4/Lfumsc9FAp3MEIwiwEoIzEWvFsWY3YsHc/JvxlctziOUbZK
Trh0M4h6DQBpIaaxaRFuZgGBlRMDbdybV7Gthplf+R1+7QhURmvBecjqCqsJQ71yTD3SOFd9Frj+
djTuehKNBELWff+/X7Tim1a3xvFuMYQYIZS/FxmE15LYNow8l7Wk4/QuaTtn6yxVKvbkGW0MEbhY
FgynO/R3vNtLxPVcgTFNQ2qinPlF6a79wlT6o4IVM9BX+7Y+CYX9qUU7+eNPlTI3UjzCNIXiFGjf
sxduC0YHjwlBh+em3mlB4y5mY/giEEF5gEz9SMJJ7C8kRPKQ+kbkYrL5b97VcL6KjR4wQMvbyY3N
YJkHknYZYf0ML5ZNmabKFWF0M9Cd5GlYJ4IsUYISOHW3i9i5F3QA1vU8H3ylZLw+F/L9YyFg99Yw
YHUT6yQDBHH7VYhv3GVt2mrTa7obdaUPbrXrDnOeLxlafccY+WpU91pp1A/Af5/bq1Y3GVtbpVf9
NNOv5OeFv2kGB9TaL6SRIHqD3i8Nr1ahtNSm9d05rvQf2GjkPnDwVsbHi6CfeIb1RJsI3HEBT0DS
Goj141nqAEZUD/5ETtueuezZ/GupVi2Q3Yhwuo476poQe3O0E1CsKi/UIFcMkJNzoxfviQGbsjUc
ihVje05lZoIOkCuJzBYpesvsjtZm0lBOmbrtHQmJExd9aHU+hhGyn6R2Tnyl7A5iefB70PmO1mv0
bE05qx6DMFLsrkwHY1eSVltqGcNDY2f8EM4W7tm2R8w3MsowcSj+1clp3ds4zQ9f9ZiBZ3JMwKb/
nw9+sdP0WXf/2aZi50jRgLNWcC/JFHTo7JJmoNEL2HohTI2o8TBXoTCGpoF+X3FUsX0qNOBYCPZ9
YUiNmNkF8rMaSwE3eliwVuGDsJJIorVHI3ddLsYNdH7w5xd17fXe9QYWQuTotvS/vW1UbEsSt2Ez
qy8d4LWi/aVzO5cLPKBJb3hpY11Fngm/WJkTHwQdLkpds0BCRCfGMOKeFcBD8WEqmwYfH2cQ/dWb
fufjOMt9QrCp30jXCY3iUbGaAKOkG9xpi/Mhkchl1pncrJ+yDGUKNojD99Vw3OftDASDjE8b8icP
DYIJda2XmM6Imk0UZYadKYI9N4e0WRY5NDj844M0OGSnd8b0ujCwvGwGdLhpCKuhRU+RkT9TRxR+
ATLBy3RF+gfRMdBbVte6/Yu+lIjPcsEtfUSv4zL1BonuCXFFVLMRklWCn/naE1k36iKkQaUL2pG+
/fERBpcIXK6FKqvr5zSr+J3rYgIlEIAc4LKFHqFag+7VVL9zE4uz9cnmMk3AXC20/ZZx+CuXBZcY
qNSlKJ1GYA//mBZPH83vVmghdGEuzGrGIKtEcrj5aaN1tTVXNuVAyZsF5NcJXZ/kRD4ZqAGL/tGS
e9zrnGGRc8InT/jmmB6jjMom3GwINOPe/iO71ZPq5WS9yVO7A+xhb7MWoFsFk88kvbiqTm02DT5R
YrKTuoX1LEIg3F2o94+afWG10MHlNl8zN9o251neOYAEGb1orM+U8DklAd4GihXIQ28Oo3DgHF/z
HUXjL0+T6FK7+T5eh2xsdjPCOzoeVuX0oF34DEpxCHu776NxcUZgRwcN9P9sfqGy/yQShHHP6dcP
Q5H/U6XCUwm9UBHY5qWIHLR04SfLywZ2WQMiwqmAtdEwUa+FQwOdZzYuixtEySJlbzP7vnofiLNJ
KR5mKJtc7AGfAEmXQrxMZ4GJXVNevNWAInQeOK2s7IB5gswJFwPE6v+Ww0ygRc0S4BKPU3+W8Lxn
bOZyISDXusJDvs6onmE1z5GIEwCcn255prWuSjvPD2s9BSIoj7BywpL/gQlHvpPN+rg132VorBii
uR+H3+yhrmD6MEvq5EaweHqDS83XnT9D0HAQNA1UjzxdgKMmxLsXm0q2ra2gYoQLQQiPll4l90Uj
LMJ95V5GzXRi4qMGEfLhcv+xihk1iLj8BJ5g0Cksq/kEpCWqc8ysLZiziQVwmuCl00IH9H07vnpO
CFYQgP1/p5TV4YWoza+QSpty4uLwnkP+PsmKyNOXQ8SV1AvSse8nsBEAbd+ZXi2IkonzkbMvF+9b
dEXn2pRF5N//mIX4tyLVuANvmC2MYgFXHGrmhfGAJGoFdnBnx67ysL0zQXhl5bslzc4Cf4d7FB/J
Ipzace94PQjgRDCRu9tS1INacv3PwOpcvXmPdirQAQL6IFJO9N/kh7jJDMQ5JJcGUPwVD34d1s7e
vZZglQfMZV808Qv+6/DicVmtPWxwF9Dp7R8u86x6TQ6IaxORw7c95hyhj2knleNbhD05CebeBpQY
wiytUnzYQ2aMhatps7E4ZTcYlcy5YwuGL3+tW/WdCExge+P8c33hoOITuqNWIBhjKBr8N6lNldd7
JuFXxBwC7LacWtlCSwJJ8dAS6a3dY/q6luAofpMR9i4xD++bFDmQIIvVO7zPVPNudqfy+R7KlDw6
ZLEh3DBbEq8JbEjoIdDs3o9mEmarWHCKNAEiMD8biN3W/elqGomz0T//pNcVx21dsNIBMNOWvUw/
WmaOcVi6RQy5Kfqk/ndHrhK1jlyKRVf5r6XyhFi90WGVquiLm6ex0/BtjawkWgcdGEvcq+tlWqCB
0BJ0VbMXjrME4nMVO8QNdMbanDt2lxIOfQpL5SpkfLTAQ3NKssI9mDG+1ue/yK2HOXWQYOjLelh/
Y4q10XuLovDr0qUYSmUpadcOqu2BwBpjgOzZ5yZ3VdeNIldOM703VEldfIqeQLY2iqBzNyHUd4MQ
Eph+4ODPArORs/G8wi7uZrNymNh6ra65jBTSbloUnMfpzDw9uVaO8/5DafkMlRj9ulY8ZUGgkCGp
R+CLduxeejHh9BCQGV6sAk7AvciXhqj4L9ziuC4R6vQZCjipJKheXZAwXiTt0Np5DcjQ/+ESOCYN
p1bYFol+vJXH2f+tO5sbliT1C+FnojhgHoG2zGzEnFTof0KKS8cBrQPD1kk9egZiNjUfRH2Uw1e7
w8O5blFDKAUGSPagzMOP65kjn4DtxYe6FmsN6CcVrzJR/1XAzGqbTJzaCbXgP14uXOKhzDL4QxZU
fK3/slJ33Q6XCT/YLAYnwag6BFDTYbUE3EtpRQWu1qDA1+8Tdwk6yfXc+ec9qv2b3LeKLkI8pC4t
P2STbudtUh0l8mdIIXphSaK/bV25vpF+EqobmENsaJ5J+pOXl5/mKeCfflnwBguY0FRhKKwWRbU4
MgnoqgQL4a1Fov7ytzt+i2/YrBUkn8TDXE+VSSvjJ+VzjKAOhQDH/p4v4C5yGQJsqX3n2fWakBsN
3/tlz6FMiWdGPz78zb7paQmnYkml/R+Sy0Th9uR9WRMyyYx3dNWrG4uT+Ta/p9lB4Gc0ctHMHKC5
Vlj8ByRXVMuVfPHFtCZiyKdPPpEgwdMLE+ZGSvO5YWqBrS3ulMgIjfNc8MRPGEYUIUiTi2KsV6ck
X3OmANm+b/hX7It3yNG6K4i/V6eQDK8nHIA01fOfZHTKqsnmG82cvR1unr4YqSne/4LVTqmmjsZj
X0bLox0FGysuGVrZFnkDJF8nGesnGCYdNZ6th21kN23Jd8kVJzzLQTsoe0DX4MYPl8+WAns81vQ0
hfmDHaDHknhCaEVdjgDeHPDsSdELU5qgHaP2mvnls0A4m2cCyP74jvrvpC3awLcGdIcYpitB1NM2
0RNzi8r83cRUBGdnpmFeA6HGXFxiCjvIjQgql1NbdGyEN17mCQ70cDMfFaSbr1YTCOQhlpeWzjE2
q9BiRRkMaGqK5oS51bi4PhGggqpMvgpJEqpwVUUDyBrt7KowSjdD7gCVTkqXADclePLS2RsE/Bm+
Yo9k5O5DNhKWWDGB9EJeiGisMU1xBZrwGQ9xwE2tU6OiAvPo7OmKqqdJPzeP5HZTPJzsTo8pqQoU
ulUWpvmK9Hk9KK8vLXTQu2AdWuXXobrP4kThbMtoDTtcCS4X8nS4uaIVvmk4gNtPK58IiPu6hP+Q
w9FK8po9ZaByjNm8noMdCVLqj4q6tOrpdeSmO4zSKDHwJqQWp3ov81DXJSjm5c0cLjoOzg+x572H
gMeIpFUdMFIgQBYtRl/ldCX4rsEE+NxpowhziDQ75cmLUrRidLfasqmmnvUpUfingkscIuAlE0b0
OwsPuGNcLmE/eq/giaJrvjGfcF1VC4Umkj/jJq+IkR/0dG/eZm4vuT3F5bOTZW2A2eG3F1SIxjU9
p/CjLFFTHZOhAstnj26/tZOltcL1ZvziQeaH6h8R3yxD2hhp0Gx0hHSB1wsfOSUlkWYgEfcdspVJ
EnSZH7FBW5d4lFealxtkPEiW5LPDpNKqvQ9HDlLVwSkcZOgkO6cK7Su0hii6OFP9nvwMNtJ5BwiZ
ux1i0emer8W8FdLSuBhaAeniSBeDVGonAleVtl81YCQeeSccj+mS1jf6frGOaYz+pFYDyxOdFYUe
hLW9JgDi6G8pi3hAy03KJ04Ge5ATmjnyIKpMD5UnW8vMqlO0305VLCLjTN7ouhuoGHRNU7Gld59F
GyVCJYsiijXsh25Xf4lHm7OVA/P98jyjpC4x9UXOsyVOrgR+jZPLfo2oniAhXP5moDKxS8wpHPV9
5R3jjWy8y3e9nkxc3SXpyGgLL2FoLZ1HFSa4Hbp3El/ECOvOJt/0wfLM2njMYez25jchR9LknbpF
c+3KG4mYx1GPWse5uZPg2gmG17a7bwjEVlq6gytTBjrocQnL6O+azWL16ZwHYtcuYsQ8LA6S9cIt
XzhZGCUYyUrJuGEG4gRpIc8CZ8Qt9yU5qabaPgQ/RCvlITNlp+9Ydr5UO9prYth6J+oWU9MkVOoE
1oT1rsXKfoA9bbQqVapHOsKSl1JOdhKJ5X0vUdfxh5pmtit4XGuWEjNrlJwJxMHPz6v/DAD1zAW2
4IonRU9qVuJD7VQY8xc+q7y5iX3o3AX/bWH4C7JFmzIqbPIeFfviX85Be2FcCAb6rXzKmh1G/VkT
w/aOPdHPkjcMqV6t/MbojztF/QWlzfiiaMK7OUszm5oY3ovEjyUsvDPsFK56sk3ELgMe9QbRPOtU
q1B1l1zCAOxYlwiTB8wrQZmL6yCeESkqUj7leZeSdqQZd4m7M0wjTV0+gAbT5hEscBD/Kqp4a11G
wGVDOvEgYGefrLvLGXCMeCfHQomPON7Hj89foV9CtckG0BjrewBWH0dgKMwoKY1cWALL7jxCu10h
+m38pHu3PyU5OiOcdl+i8phd5n0lfleea6buV9Ytl6m53NNBe+xdh06nNKQCLvcifbmrg7p+/tTt
yRwF3yuDKc32TwYsshFNottdQN1E5Ya8VbDwPFtVTtgUFqUUck5/k2peAjNahlIRjAGD/bQHHAU/
cEDspbBwPcDYfMCMRPlT4f4Qw/ufse8eqfqxcKwIiqPvyDto4nsyYRcDeRrW5t18O69ruVUP2UaM
51z2wsWkp2hKLizyO5sSotMrQe10NX29XEZXGGM4yJNRKbPNt0Kk0Y1Dczv8ONMQUIU+fwVRN+yR
hgjyQRrXFJOvNelXt6X1gaP4n4iFga4gLnFMFUbmG0tvuKGdqpOqvAebmPus6NvUqPGY/uB3+64A
NJr0kpq7wxuyfyBCr657S8ThLpRkpW7U6hDs+lDubN12fWH8g1MqCdlIMjP+B90dTMMZwOHffO3y
5sFtvcuTlPlvEOhmhn/rtXs9cMv3Exr1uVG/0gB0x5Ru0vYIv1Ut33bFIqOyxoyBYkNPM56trR0e
hSb/lUJR5aR0LmT2zz7Lh80hFTdMsJOHNmTk8WYJuuMtuHdgIWNyo8a7TaAVTiBYW2ti+JzwGbFa
+R/Go1+B8ylPERHoZnq2qR10xxiEIkSWBLhf5/AeiTk+CgStQqjMv6JN9rcxTZIq1xFS9h2H4ADC
GTHBwVT1y8cmtPXxZQE9k/pG8ss4Jssv7X5oCsnj7oIZN+RNr/Mi7eeAtoSo+rMuxaG3IohI5lCd
6un60bPGJKnyhEHJgfQKLyWrvAOFIQ8xTMvTcQhsBmfLN7xAnMRA7BSsIzEH8wdQCu9m97zVAFdy
nupui6FEq9ZZgiXhXB0ZITKEgZPA4QM2IraYtdlXaoqOY0U7lHO1GPAQme1+9XxvXEydBgpD8goS
HGSG9RthMsgGI2nxb6BNhsYmivNH1l6YGjbVwqtZOMWTs3ENiEDv+6wq30Q7FRGsuYhOHrirInhy
GvDNn1uY+kcazP84mz+7a6UU2JSzTwxFsVx/lYfJ5sSLxzmjW68USq40zrZcA3ZUbs6IaEeWIpwb
VASknH5hcmz1EPQlWgOv/QLJZXqqY3u7Jq6IqVNAtHe2Bn6r+YrT1q9r78tpyuT8aEUpz6bgn+X0
QqdT9kepSUBpLwCx5AtxarNTMBLL0e5m607hnfXdHa2GUvizDYYKILiAkBhCGbtOpN6bVx4bcxZe
NXKJKknw2f/pWnoHkQQnJnUeJ0g3A0gqyVtlkY2FWGvbuRlhChlXqKMD421IlciWprk4DUC20sko
qtDx5bJp2lYJNbX3pP8dOjr2ya5rJ6qhbXvo7duyTPCURcghI/QH1bX9dZLoubiOg+8pCovZOHwy
jFW4kkFX9QH7iBFEJ7ylO4Rfwnrdej45paufhI6gjdUUFFR2MPQ7GyjXbxUqupKYRJziBQLnAS4j
ThlyP3EnPTl/qbdYHhhzUyhxdfeBc1Gx4RDhR/6giExCRkHzKw2bwTHC/6EFUVH5JdcvZpZtClkk
gwb0OhXB6sj116c7T6rfN2siK7R/A8ZzYpOCJsqxMrAOdU27Dp17Dtct8wbw0lMuvjZj0NEj/yfu
shGkSPYwGJWiEkYmAFuCpP+tqNt6mkTlyOxQbZP8zUceHjHL7qtfE1IbFggSIguY0uj/Tun4YSc1
1wenQ3rVUOIR2J/4nvaX9Kx/FSD0GCsjYzR73cVQjznpZL08ra5wOwWETr8cAGn8u8JS9WDNZzid
yyIhkR78+CMsG3qgMeZ9xEVNSTUZli8Xe4BiN8IsmOW05arI5N7q1I4pWbQgdP8eTJ5skqw8izOy
AXVshuSso447SYE146rqwswQsfTab9U5RzLziUgO+WS1e7sS4/8wfJuYJNUfAv+gzik2IEyKc2GH
KS+u/bmAKNZD5f66RkvzCRPp3kvtZ0HWQ7aTvF8JDsiaNQEGN4OS7L3w7texFZyOI9I/EcLVG4Fu
XblGmTrctjnsl38bZeuYYdEdLD+w5GnaWLvyRb+XZHG0MZEc6PZxhScDB4HOn80cVPNBgSCSKw41
QzKZ3owS2L5ZdJNHnp7t9wgqNWmOqwogY9RkB4RGJCIJKvMFwz8X9wSwmWqMHzIfDrF4hv8CRYvf
Fvtk1bS7QvzyMwTSHGfJKH1fmRTnjytTggqKCjvSPtKsLnwjNN4CX7cr2JSvUqrQklx8q6RnKVpy
PBQ5JYUHHO++sLoPRy0cUt0SMfID1TV8jPLkMOgbYf6mbcUsDp2Id6TUGXkwYzI1g3CP0r2YvfDJ
TGMMtSYokthr54EloiPYMM7tlRB/xXvOgCLg5ARwtTuCC40oM8R/UGcPv2qsolLqxouWLz1dUKl0
m61zXbOduOaJbeNKgOsUz3RnbZvqkjDWMjWHrjbIf7l9Q2b2ZEinGZT36XumjDAHwJc4KGVlyGSq
bYDboRt7bcnK/ZYmqJbMiHvbQIdWZS/hcRZbRD4DaThM58u19G0xnOZEC6d/o0l1Mmqiei7dWWw8
44dL0zEVWCTHexKTKHyye5Yh4XSPDAmgOnHdl9eS0iczEMZrEyGE/J9lsJHUqdXOf+JMvIH0JHFI
Bfpm9ZDYKRREMHzoqL4nmE0ow7QOUtebb65BPBK9W4/lsvyKqwdahXn6iT5OBVQ210pX4IXGpaN9
WoJBLMNh/N06gs2U7049VX0lmCVZMXjSedlCHhkHSa5XeBZpRafrUz0Bz3BubxI9FyjEthUShkv9
J85GvKld2NsFxsrBOA3JlMyQiNjB/xdTgcWShHVdqA7+bUxB08aYc9KXFNPDoo8CQ7m1o5Ame2jF
otcmPgMGQbKNB6637x7uU2pes8xx/IUDHu5mMQszIK2XJ7MGE4cL2V0YBbK2yzvtvE33Xe0W7Q5q
RzReNfvOyfEPhKkULZre6JXLQitwy4DcgNPzSUxDtv4gLUGV+fbank1DR0LkQlLI5/olzMXoPcpL
/i53crlnA6CC+IO9EDTGtxdjWpulsQP2Dat9fZCMLVc74l+l3HWlQNdUCmkv1n2bBo4w8hPCwjjT
1VqyFW/nlnZ4/s+LGpn96phjQyblejEmw0j/UkWiPoVVqlSKJHLQAtJ4A455cswc8jtsCh8QQQUR
usZSEewNyYMNDqjX7LyvYpj3Tro7DZSLx2uiX5jbs2pzTZX0myb6GBwACwNB5PifpE+oAHa32LlQ
WgimI8rO7NVH0HHAAnPZxlQ5isjJ2z1Lp/QbUWwNXlCN1ASGSk1Jmwn4cntNNFAfFWr4iGI7Fwxz
JPCzOXxXbMohAkAP5l7TErGVmblpMGE+Ce/9b1AA0Du8mQnTiv0ZiQu8q092OFVjUio4Q0jLxbpO
RIzPfKqnhGyy/+nQvDKNwFjCBk1RZ0skc4pm3bUO3fsIGw8jNxxGbPqaqzCUijJ0EIVhiNBgfPTJ
FIJXMpI0t1iB2GFoJYgUTxNExNBYnA0uT3YGaS2fzzMyPH/CGm4SXiSIs17se5BRExEoLLv7se00
98lGxeJo57CGd2Bt7CgDNVVYo/Qrsevea2sgUXCQt8BaMd7S7E8whU7ja6oIoS6j6txaOCNIk/VR
aySs+dnGdS9WvyNlMdrlpv4iHJjulzFFlmOS1i7Odt7WPqRdyC+swuLx5WXO3rpss0UTxzzBOdcW
dKwi1i/MllNt8oKf1EHkwr4MarHBZSf9xivoNXX2jm4X0JOKXEhD/zvL52++oNBBR4F6HLYo0dzX
621p0UAFrjREDne8DtQHO4FSCZYm8l3HOoDFijfh/iw/3QrjUNk6MsXjjOyYBA89KDeE8qP9ibhH
PVRETR1iQvC+QS/0D/BPvwlOfvtsgWLWZSo1/gvvocGM8YsV5pAyC2sHqICMCCSie2hzdTJwtmzE
Xi0Az+nlb4cEef6ZxEBDQMCj4L+6KAoemImP3rlrMjVHfR9zaV3cUPy6adG2Q5rJtoQV85HOSxdt
4oLw1iAZaHhNbmV5yqJnFGkYtfvZDf3Ck51JdoWxqTXmZn609UZ/HJ8l9ZWfevoMJbaHKkyMm7hr
q44+7krnHj5fIsTxiaSs+skX9Y2fqF1grG73t/m9UWlKsOcy6fr3jfsM9wUqgkeOOm2e/bDGLqNX
/wNAGRgDlWAnkm/Swzr94cZGnsf+7VY8ldvDutafxlRsY1ieAOEA6CfeDfUZ6V26jmoJqwM732ON
i1NJsj8qhgYWacjNj492WaRpreE6qU/B00TmB46UNU+JFViC8XV0AJ9j6/Y+BkqyL+9BYS7pnMTS
IdJcWyX70BVU6X3oZVwglw1A3H7fhq9jDD140Yfa/jQgZiVJThwMezYiPmsR2Sd2ja/Kv2eVjUe7
Cz3/Ly+075CBoepR2SdMk6TkHfBgx0DMuOFqxSc9vxFOv1HcYI7iEEbcSq8dvU6fvC6WW5lDNbps
PKPtvaOEpRoVqm+om8c+ONNf3kLkgOHGeE5wGrTEabaeVOj0jyV0Hz3QXSRQahCRH2kOrj50IqDy
5jSMCC0pDX4ZCDYvTd8Wf7RLBgklsNZOfQx3Uv/6KQElrA8VhAbb/PL0jtSAihGuyonLNyDAB3zY
MotN9iRgbU4VQxp+GLpOuZpxHHbZOx9ytdJXqqv2H/mFkmoMChB+Xgz9AChkpDEfJCNine/PL6cp
ntbU4rtq/L3QKP8w2FMxqw3WgvCdimdeCokKWhH8J6VsAgdbQGQzZ0zgMayrzCfPQbLGlyKC+yNR
0c+D997E2B651/DI9uSBaDz2Hke+pBDMNP4K7RQVVVEE2A/mJOAXCkJ3IkPPWk+AxvwTXKs9vMGQ
oh9nIzU6GD2Y5dGtZW44kA//ZDYkm2UFNqZz9Tt/D4KcINoSpdR7uWO87z716IWcSnea6Tjn8jl/
1k2m7YTVe41AGPL06NJSL3cDs4DzWl1rsiP4YxD2A1qn/ce/6iGjjxXTti3+GNmFXB4p638uKcG+
d9zRps29KGcEaF+Az3O6pHCuYV4dywPf9k2EgAf7ZIubNUIDx6muh87/2bw+15HBn/9Skptsjg7D
LtL2nQeScz2qScK6oy4WiICpo74f/1fM9r/s0M9ldT8VySiOh4Yu+dTPLO58Lg3UXgJ+8yasAt4g
jb7x/RR/X6KrRC6f/UaUS4pWna4imL/Pe82UwmJuzApoupnFK8ucGUu/ED0txQmSqLO9Oe2BbVE+
FhF1j17KuiTf7QYwv1UCpMuiQfzNOzV4hzWXApxK4CYFYvhSZbdsrXaWtllDbGUr7dRIkzc7+7DH
W8gE8OjG2TbxrrDwAHlcyhGtvRbKtRqCFF5PNuYaUasxs7nQtXHpWCbHNoGHfCVU+q060JYSqno6
Bhav0YBLMfLA3gc9PRGgKcz/xfAGvzix9DWEBDgVv/NPwckKZklhCPuTjAdWL1Tizk1mVbU8XgF+
3rWaTHkXKus/mpc3/w+tgYzs0gVTgYspjA3FYJiytnipSO0OtcsGa0njJtR+wPF9cLdFFtxplQl7
0joTlD7IB67iVFAR7LPmHJK/A0qJwlUKcSeaaX1DB92vgkYO9pkWPvO13iaX/p0/iutba4mBK7lU
LP2cXB1l+/tYZkayGB1vJuwN+Z+1DawByixBuHo3LmZR7VdbbX+F7vB7mzhgpHG93gFV8SpjMQgy
u6S3cbxGKFXoM0nVAZASLJTHDpCXzdfyqFjw8a73jixPO3A7npWcAaKzQ3JKQM2OVylNoZrUgAK9
T+ewTnMt9q+Zk9ueruqwpHmp92AIm0jYnbigs5fI0jdh6b48Vraz084jqKiuC0XxGsvrZtrGeNpw
Bd+xf1ZPw6DcE6th722x1X/C/J8gcUAYIR52rD840kx+chQcYRL66uCY0WNyiK2jfgACqjDynv2n
Hg/x03AUZz4EmJI+wlIOz0Vzcp/0LmeofsQwS0GwRDcK5neXzMx2+DimuVlW3abswaweTwnUN/v/
sQuAOPUlKUhyAS9TL6XuVZODlj/wT6eEpk1vC3icIVWNqBEoCLU04i3DEWXE5R6wLlR60yE5CHnj
5BANMfi+kr+Z4RsFhtxbf6a7WnofCnpPXQs5ao1Mpw+J2221qU0WxNS1BgbxbGRb/sHndk7Gh7EO
y/XBbOdUyqw9LjRuLWEzhVhn//mCXjS8sG89Za4nVC8RfUOyJLeJsVzUUF0fL8MixGXGKnd9QMKc
K0GUc9ql+NkGtLWWHYnY0zpADstNJHxVRZykhUR5YFbbaWYA2Wbg3QHPdXsV56OlZ6dn0/zuARl7
5hr54SKT2KsL81QLobKV/N96yySFebub7gZLUQTAHAG7AN+FHe8xbz0uyk4jCedSWMx72haPnYQX
UyFhz/fhYh3jZ9dlJ7HxKpBXEmHQiDIOa5hzUEZ6JNCg9K+9JEmBMrRto4OS867eZOCi/J0fpHTE
w1CSlU3RysgEF+AmjihNL3TMJZJ1+XVciLLXIZbmWJOnvx5OiRZJPfQN1TpkmDI2sPt4314Taxl1
4vISyFfRZxFfpszhMr0w78pDdPCMDVCxWL2X71EXWyCjy+gILEOMr0DdRiAkG8/6+RbgzeSENhZ6
sY/A5J/6vKsYPpb2Y/4Ilf6p3agrFABM1Jdf/KK8Fy4H9oQZOY5Muif3RGrlj8uuT7jgo+lw1S8G
2/igMGfNnv4w+XtXzH/1XzDZ2x5/xL4Cjpwi8fjYBpiMmg3khHlmPkHW/qjnLvwxAhzUClFO8XqH
2V1VbJ8Vp8BPs7d4Gbdqn46KpEVHvuCKVFchu+D/Lu0ZktYwFZ4A2YpIjrWsrwfGQJKmE8us15/k
RDYdPS5dNsXDzs6vZtY9FM22behDX9YMKmZNPlnyNTR50sP4+tpZuJWBlcLQIhOSJus7nYP2RC3Y
Ns1QwbYCGfJqmnuLRdh7aju20U4tuX6yUw+TYhFhbW7Fa/As/URMj6yc2k+DslosLopBoNx4MWbI
txXdqZgRmXyGhSdRKL2emKLXQ0fd5D8j8XqeaM0xyxbi4qMUiPhebxwi2oPQJ4cvdXT2wa5v/GXI
xgj4UbsQv/GLq0SthSCanUOJkr3mhx3mHMGx3OiYKQznvqltsD9oegt73+k3D9YbWd8Xc+GrpPOl
EK3W4POfXQdpCydhj7q2LnUgwaKO55EPDX4deJKSihvDTYFdHWo4FXf2lFm/vqpcneFd02hPCZvS
qmG0sOOzLey0ChEOn1kJh8AnfX0irqCyx4KWnIZJ2pN6Bqz9CboCEuPnmBPsbO8GA9ydCoaUL6j2
+hN9Mrf0WM1MJQ5Ws0GCz4v+nNQObuho7uS3d0wJlgZO1F7mm6k1bqo1YZDBpRwbMQp4GpXYnuH8
iGDlvQZmmbSejc8lGGUPHiHto6VR0H2JfMOeKeTXkB83r6Dm5sU8XgWY/QAAsoE1NGgSC+cu6Cxd
9KaTxau+zvrGWIG9WslVOCpUg5+lCohF5T4nH6c8UfR0dmOOwWFsRpGzE1qI4+Wl5iLQrmgViLHC
r2MYcEp5FmS3+pI3j5tQdVdfV9+7ZgI7bkn1tP+5uvlSVuGO9kKj3BkVAa4xFJ9+xIksC80GJl6T
9JqhivdJycvSKDot0/RfVnuDC5LxkzSEEZg1UKYnVhjXXNLqJX/QMb+Ht8H0JZQF+EhFEVHC25Gr
3AG8CMpHacJo8pOU2LuUyy4DFzzt2cVnR7fHfojCuDeAvUJ2UtO51Rru67ReW7OP0G+Sm7hxfeOA
CgAuBQngHz+SEDFe2vHhx9f5ubD3iFWcRQd9ZgbFwfeVkm1TtHj8ha8apDzgrFe9B8qSF7ryUgbW
lYS6eQElpO8accDgQWhM7sGPx9OFUrv/SiTJUrFafmUPP+QTddXgbA26SDNIVRQ+VUT1X4w0AU6F
XbSIRDCwICpodj7Mo6Nc7Qv5A7GCs965jcWzr8pg0fia2k7iGcr+eHKmJFxzGb5bz8KDpZt/ilC3
68ySplPjau/TFnS2HOQg/hMfD4Y5IN1Kx4JLZOTnTtxDDfwxrzeeLVHz/TeBCN7JKO82cEHInyHq
xs4Ch/fVqD83YVMT8B9b798RsGyI1sTu8/ZVdOnEpw6Dy7qQysf2tOxtZ3pXEbqgh0Bw7q8edok4
vKTOVEAcPp3UvOyUNiyd45nba+UkaYjvM7UJwjR1Uz7QIrRaJPlVelHkTNXhb+/IwtoCQzKuTLEV
h9pc00nfLTqJF2Zc3Ufx1QveJE1nNR0I8HxlPHe4mkYXFexgnM0M8KQt7JxBoCK67zU2H5o8KkHI
nisbkwt2cGKDwFPhDsfHsEIYs/ji/NtQikvxEly32vAOFF8zhkEa6PFPzcTQqWwNo9RW/j0uLxd3
qRHO263RSSC2NwodqWMJl2LPMepYLWviNUeGBvKQejosDUUQLaFVVgu/3r06kzdbwdWo1HAH+sSa
uisGsVcnJEZi/4YFO1AVZceD4QwUydz8Y1q3p8Hdc5UxhUYRw+UxCM3H8oiAc8UWGH4zCj2bmC41
Kw0kjXu2EBnI1HYFnN/H2DY3OhaFJP+mgTVRyaMJ4sbl1mfNibtG0dcwy4r5PO/H9mdDPHcaRw8q
vBp+mClXa/VKmPtuvab2GW0+QZ2U7p15G0J5AbWTFbCNSTS5EXTHv3chuwyZTeLjsL5wOmrtO0+2
q9eOC7fliLQ3vFVMctACw4K7JZHs8M73svXxW6q07T7ygBQkMiXD/Vr2A2FLsWmzeLI3/uK4bGxD
s9m/5Pi0JbjxiLtqGZhXyHrgvSVoCSwA3yKql9p8gJJw7Pbtj39DF9kuU2943XCf97GmekXeW8nu
Gl1ftLXW2aZIuhujNglVbtjLnJxaH5k/KCaNQsXpVEbr8vFCpTQxjnpj0faON+CjxYM54bKVWVLy
PdCsE74AWju6GSG6MzDy9X9+ZnXdSvHyLzf1RHcLnK37d5rKl/GajCRCuvBSYfMUJ6IzvzxVLrb/
YFsLEZiyQWLCQV1imQmbqYWHu8Gf0kQCXZSBYhL8Lh6KZy8BzNojtwdnQUHF0KddA5HTIlogBLPD
yM5a5Tp4yu/1Kf2JyATFH5StOT0nHAmyMIqJPNoNmhxG2VwVaBlyH3b61NhKkYsgOJ/ZQjezVZYs
o3u2crB8/D4DI+P+IAv4CIbyXaWACPdd6tBgexTKiFllt/T7Bk4PZDbgiIflcCLy5zA5KeEtQq6I
XbrZb4dda63ehzjvARMJXI5CjMu0Mqlb5c//AxmUMHNoZhbbVGLXsAgjw8V45UN4CSO2yLvNsHsI
N+5QRNEeFJvkolBcLvcM8ORKwTn1YgliEV7p6adauNNGxb4RPvh2IrBK4uBVBWXittMTMcmTPmB1
x+8HAy+k+06nOweki+LMoHryji4a2v8bHxUpVntQj9XWsG8zKGH7nyiI7UR75lSC22kdjQfz6XUa
3Ht3qOxniDtqoqvMrFl7y81wULJBE2tBm8S+wL/WmJinViNxwMSGIj0zCZ6bbMaXrPlSFlbKg2MI
EUO3nxxy72/HKqNDCpdjnsvj4DqM7iuNh5CBrYZHG6H6Px5+0e4T5dPod4ow52KO4ksYx1HJYFJ4
SijKqTQRymolY12vbR+UGE3JEjU9RQE8lBn8uOqjVexdzRPyM/uHKM2T7/1FfOEMyOWi/byPjlsk
X9jU+eaDYtUq+bXkHxhmOTEDLroRZI4IfrJO7CxZNgyCPKa4KBLdQDgg504HbVTAMCJXBE/jGbJt
HayhzdN/d01vRr2kcDwe1Td4L4a/veg1u9mKSKaX5z/VGVi5ySx6LvTFA8umzYmGC5efi/a17h6/
Ezq6Rmfp7Tlfg3trE6gRF9qlXMEVJKRuR0B1jI49ilxYITIihvGwEQmzlkp414O1xI1EoIZRrgRC
UW0TX/sI327lDqNPfpUva+jO7yw9KD9cMUoHLpSTfglkuxULdMZUt6BkkPTfqW7Aikr09MNPNtjm
sDur6Q60ez8UKqU81Xs7mXr5SeLVQmxWJjgSYv9EM4a0ztEWWLirrPAvLZWfFuldnrky2CI4RFp0
blFkZb9IMBfMIiox7BD15VTu5uTVk4p8cF5NORlvZk9kkucoFC+5NGX/QLDkHrjAxQvwBUIgWgOj
OHMoWS+HnQ1FFjA3J709dy56unz+cewmlUJcur2efm2wBz/JjVHm9AFZ9fHdl8cfYSKfdSvj+czg
mldP1AjWzTXD01/vxe2nizDK01CpBOW2aU/gu65zDtM79kH5gI/yyRfiV8nnp2K7a3gP6vM8dUjj
0YuFJKhIPJUN/QKA8KqlggeuOHQA53wJexZOpudJzIBmuACLX7WkoS1L9byic/FDOoSvk7SluIqd
3uQkWB04GbFbCmeZI3Rz4R02hiSKSYMcfjuMFxCQyU25hC7icXIP7RmH6xx0WVfi+b+g8YVZNmoL
3Sj/3/UmGNiN1eI6pXVzfhoCjHrYfM9ZENyAgy63j5hX129y8CvubFpbhyuS+eyazLVPrAvFxZOo
ndJvrknqWU7er59aiQkHo+Ow9UMf+EJB0Mh4y9KRxqrKYYfUmMSgNaeBp6XEJf8KSCXFILBrm/en
qKJsw1Zw3pZp80VNf9ML6TSWCFVqHquA7pta8N8g39cmXZ3DNs5mgHT8qthHdAJWZNEZvr6b2+Er
GTHh/Vmtqb4uVfeKHEPFGl/Sz+JTaPYU9B9Lf+mbeN++Pe/ZvsgI5K58MsO7V0SaWK/XVgxqc5vd
rfh2UW4Xb2GutCaYcIOHXrs1zQO+yWs/jme6oQ+IUiNMpPVUNsXC2Wt0cvZEOsyVhveUBhQdw1FK
XHxnOCWv8uXUuGKhhmAtrcGxM41HxfDoFmJvFaYEVGANiHv5AQwAuY6B1MYvOSA4RwvQ2EB+rkbS
QLYTVbO11eP5QDd/qJy9pJbJL7OnNPlt8bST0LMi4A+H9FUfDdyIeGd5MpOek5xtlWLREmIP3M5o
7yDKKRJEKn6/os3fGdqLuIOfm5TxpQIXEHWXepU5xtizbuULWXMqq6rQfQSFDJynOQlRMFepkN+f
bBqMOtAV1TtcWOUNNUCN5WxJBDkT57PctebJfo1dS/HbzCoeTluB7Xbo/jeQRw/ae34//GBF+3kY
S5CpAiE2lN7AUhdg/CdBaKvx7TD3CEdeQi+4bYTlQuWHoYfFrwN7YClYgTjT6o2PowkGGEufSnoF
3zIyEFvM5teHfVsz8TVYlXGHaqYG7QIuhru5jI/89/nV+bwwQWbQI4+mn9+WLqxbTnxJLjyJWFUM
zNzazkHE5r56skO2MCV0CqhFpx3GBkBMQSQR53zr3oy5Bi3JurqoYjgsZ+c1arkv4mRXxdr2Y89L
p2Un6tktI1Hwt+8pu2yjeIl08Evvfxxg4s1zbhTt+2ISkxa8TYKusXsMnqja7ZwXQszQ3US4/QEs
r81Q478mHWdokl4ujNfroNY9RAlj2rMpR63OJsOdJLJTfcXV23fgs7lYD+EC/oiD7PCXnYKUK1sf
VGgdzT4VnuxqwBCzbAfmQUmwqDnk62XZtfmnnxAd7yy6xjnYVfHKPcwO5VReSkE1RQapzV5TnSyT
de+Cxo1z9qZbqmOH+vPHn1FqnCqZ0BAt31C70+XSh2E3ng6KeVooT2PWM5qYO0GecPZ7y4eoYSPI
bUo+0y/0YxQroPziWWqHLyGkTd/M2Qz4DDnJileTyyqCzS0drOOIb2RESuvpOKDBi7Bi35FwsoGR
+QfVLkK8NHdL/E/SuUdC96Cc/FcUpmLsaF2qAUxvOuMw5M9QxvRn9O5lQQS2tbcuc04C69ZOZd9M
WVOoVsaLDP+47QIdpvzuQPYS0EJvNlBlUAksNbWan8coG0j1z++en+tybNX1LGQfZaZQrozur90l
4NGRzCViUJhcP4SvlzgH/qLz7L4MGpHIalN7X9bfeMWDoQH4hG8RFVIGm5NSmMcbTIsWHj6klGhn
jbbfex9ke2XY8ua+SHK0qloyrPSObLPTugR7t106YTPE1yHCNq34ye5QreDjnacBB9C2LfF6/+bi
52eXl8flpyaZeoCZ7u2CBexgFHdEqSC6sIk+e5E22xPYC5+BlVplPO6iSb4KG6MpGLSFFpPeimnY
4ynxqVAy1OaLXOM+wD1CtUqbrF9FQ6Fc5t7mzZmKKfkSScB6CvQI4uB940rNK5JpbNRSLEj172rt
I+aqqNM9jxDWzKnMXTMooxYCyqXCiBlPLPXWEQwf9wbfSmQRvZTNaBucZzfiag1oonrULRzvog5C
UKSmBam/Uwid8N7ruYO4EOVNhccO0Lrs4F/bkRSh/zX0Av5PQ/LPKCCQS1YMtt4UhAgodXHnwOLr
6DCvA3+hl69c7RN8QaeH8nNOfxe8DM3AgWXtByu782Kw0k33V650QLQ9y4Axvr0A4oYX7/d3rYO6
fSlVNyWNZBp5wGA4uA67/Sx4XfpgeQRhsLPGC76+8YPm1psd9tNC8q1aBuZpzSohTgrvQ58rgK1V
/JywBg6kP7GCeQiGOPewgiWE5hzTwplFsSt25xbDfWGUk6o40sI+0pUAFhz/1cgOsJtP/Toi3bYc
tL9uyhRX1vpp+RC2cSQFaz1TyWj3WgFxJTgnmVUazwhYSq3NBYcyV7BT/TGztSz7tJhd8teG0qhN
4ImirWJMJ8IKS2PDLLFxx+EoEhUDwgd/32buhiVuVjbrldEet7dec0T4o12twYwAxjfaII1vLfPv
D9BTWk4KsL5heNNgWhKyplQA0sqZZLdVxqhWR7crsigQmt3cp5P7hWzjtN5oIyXIdN8823KHzdML
yUUiX1frC2qoyqOC1V7zc7J7K4gJdpzGKOeXO4VCpkJMFaWj5DGHdsgHXx6M09FIRudaQ0wSDz7/
x35lDsMWM1IfMJmwLbZQyE+eVTNT9b+efPVayN7QZAJrmDdnOrw5xk5ZLNumdq7vCaZ0SEo+/Ezi
h+J+9RfUfCjcVVaWUMEEhwbo+d77Mp9KKb1kInUnDKVCvyAPmiVI1XGAC3GKRAlMTWAIe+8fCdnd
jhl1woAcJWyUSCYApVk+xqOQouMGzpVyv7NSDejeHc3uXExnBmmTg15PTus6hi6hycaWFuceL7w/
sx8WtuuLCGMCQd3Z2etRkk9Grqqn/vG4d7isTAUiR80QMbknVDXvhOOK3FEEe910GJFjTR3f8u+4
2/LHeZR/j9nVNzoCEhD2W4odGw9l+XAUi8zhUJwBXSfqw9u4qXtaLfOVs43EAU/lA9OVSwZ0BGSd
iBjLMQS2T+KS74UVJ22N4Te2z/xabIFRDCy9bThaXeP4NorVb0ynGCq46faxNM+ECFJiV9FUC8z8
zTlKUIoyr7PezjbxvaLcqrTnsPFaIuGVFrJWQNhCWPx/Prs3mHFiTCzaxNb1lkkyGUq6i2Mjuy5P
37lqIZmBr6Qyonj+EppSOUqYZXYGQHcnVye5ZTJGsqsEcOdaJikHdD+AfVV0xW9uHZaOcbU39v2x
hVoj81Tm9ubTyFXASjgJGZ77XWM7q/UIsxxoRuIgicsElDmh+AZpwHg+HIp0dNiSwlsX/0nsrIIB
+RrJgpb4hiAliSPDOP2zq7cszyNSvxkvmCz0Upds7EKhnR+YnuExghgdQUhyXA3LldOAieOedVCu
0uBKgxcDlRFsHE0bMruy5SWyemFPJtjJF+Cp7VvFUAzMx2AIkeF3XnRBTXmA4aNtqpNgObo2BKNX
DDMOzUW48fAkLPWlCZp5hEdERtG4ARPRmebRH/ZwlaTP40vlyTbtxtejJ7IiSRuTBslmDz7nLpGH
yVYKphe9HlpSV/jNn0Zq81ygvmPZQe3V0mF+3NdiUwfIpQDW4hhW3A8ON09r/WGIsQ/iCHEA05oX
GJYL+zyFqj2JNdkKFfyt9fmPs4L39aG9eOQneu2zSJaHgqdt77lEn0HsZ+yDP/YRBMqgqQsvMdsD
MG6mKukTQHkZkyKA81O+JWsr57TL8fv7naUvyXq5DlU1MDhDNBPy8ionc6EFfu5OSdWPhzWSHV/3
q7vQ1qxEXr9P9DLA+REoMY+2B4DYX/Gm+SazLpiXERJRYFq8mUNKAuEJjumuzFP9UsbxVH0ahSFc
AR466wbV0KsTn5dce2+c4aOFFUqAZ5oxJeXGOCRXdf4SPiVmQFhUsG57OZYeFtwE6RcH7DG+smfE
3Z4mgiBdAu16RZQinMmwVcJveS3CpLQ1YY3vTcMJHzx+Viu1jy+7L0bSB1KYbnBFtONrDJSWXxnt
+CYPpYmWkf01LyR8ipgvY4hE9BeWfdsqEo+MCWxT/ZdENt3aoiMdJb4422hHRBk0fMCV01LzWWdk
Nw8pOOy920s0GwW0JzLhGOzaxwnogi2SI/DWhVpp6Ja12mUoMcJY9d8RsR0rSMujPdfoYf+ScHOg
TEACjMJ4X6+eqT0fgaVSLVC+GNH9o+800mF3xoLWXgXGB6jFrL/OaGq3pkGsY5rqCHn8KnMQipki
YsZHErO/Sozj36MSrOIS+Wgk1LSobnT//DaagoH0zKXalY+NDq5HaBPrpIa/lI43nxR7mMXkOMfL
wttou++Xluv/nWreoijwmUY8rD/ysV7DHzh/aaQALmY12UuJ5hs0/5rTj0rx7sj4MQFElSM+O5bW
L7s58kFId0sEJ9KCoczVPD0znB1KRuSSncw4DrPsmRIdpBPqw1Am7I56VxD1XjWT0AYTZnMnCiTz
dEnH/vNNvza6UgYFkNHD/kd7kleIJxWAAg0cl0zdaNM+x8IoFiUe4c03CCrrln4c1RJG3mITHbZb
i3SgNT+ZPnS+by1VWfMguZ7iG0SNAl+nDAmx3dP9JLTo08H7P5L2qiqRolxR+/6a93ZJiJIiaQ71
uVIrXcJs90E0npjAPzdWIg6ohh+DaPoL4H6m7xMxFwMzv3bVRnIpoedyoaJNM1SmgJS0jVNySpb7
35W8wkEkMS5y9T6vIlOw8aQvVta1jawy03Caz3s9kls0hbfy8wPZ6gxiNj8Of6ELqYpr1Qdazj9k
SXBOl7sfQCK84Z17cKvVGO7yMn3weP9+VJh17GeDy8yXxD+7k1ykPC8hVVZCn0JQe1BegbqaQbhT
xA6YNl0dGB5dn260w0znEM335hNjMkSHVVMU6Cfz4YROZ4/hTj9XGGbaNyRvRUfLFGfmEsr2bVdw
psJ6Fi+sxuKnRLdhAe30Ku5ZLSywgxQvJLM9gdyctn928PCOtWmykEoTERlGNUQ0MhJtJge+bPgL
Ueu9j6pzcTAO1dtklopx8YhePB7GAXheFHFHCg1pBAfeZXq0EKkRKg2P7SquE2edDMzNrRYI3PoR
4pHHmBGJbvAFD3RgqEeN2nK4fLz/nYH5YMcdDblfHWfJ/H2M6hpabRMN1A6mgA9txlcF06EWIdiK
cpp/ZH8R7J4bfXlTagFhm6bVr3Lxn6Q0adYiY+ht8lT8jYOb7WjyafAvjngAlybLDrgR7Ld4kXWT
NID3szVw+yXuYL/TKVMWoBCBk9fbQaDLyqZ7HBm+TTCDSeKeXfoMJpInt6peP+vHd5o+wcvEahUT
fcfoURkGjeFfeRyzQLAu3UM0zmOz3INouF+NPtzJFfrKOCyak7UHSvcMemDlfcQTZnEy5Euqzw1u
4CNLZEowAszY/xEkfecWluzEZ07PMSq1ygBKXjmF9HB7jlo/yQf3CqP/dFooSw4Q1dEDvqPOorkE
lLJUu4btm6YPytrAI9MdotSzS3g65NxR8HuAwOpk4CV7zgfLIaWmL5dww1AJ4Aa+ZWLGWvQOHSsP
T3WnyQT0Kpj5s6SQgfO65uvlNM2ijT1jCQ2J2yXL7iwzhdbHy3UqmmsnKNUhSUmTfWxbC8t7ZVAi
YbXhTFD+Tic9hwzFK/7se/T3qAVeV3FGSWp97o/7IXyIIlMV7cE3IT98FqRuEW29Yi7lfjyv7uZQ
9LhvKRExUnb+cyBGAblbNCsrl8NLvCMqnI5ozebqfIJA/RiIdWKQ9s/6QVEG8A1IYCsio6ZV+E+Y
JPOzFPSCqMrJQSsfxs4hqlHPjZvuv2Le06ssA1gCKTIbaly/fDz7GCTM30KQCsU045Mt0Ro+l/la
l7LbPuzpQNei1FQ+tJy7pNMd33jDkkcHdSOXk3jlIucWOAwVyzy9B41CHEzSM9raYJ+bGpzL7Tmp
fkq8Lcn6bxE8U6CgBjCoRT1hIxkjIdT9ivjQ9CyKDQrbj6Z12FkDqLcampMd+SVj9xTpo9KaU+44
BZvaWt+Q2zDjl2XtXUR+8RpWd9dAq0BgYDgErHKKEkwnHMM2S9RnWMfwtirmRr2T4Owvh7QR5LRN
82UhYO1whrqf4jC4s1SzmKedY63Ll7U6Phlw4zdDjfTteBcmEDlrwCMM78fQ69vd3nMEn5mX4C36
ueqdZmfEbQCnO9RmEEpfOXpc7m9xG4xA/YjAqx5cQYvaTEKlnbQfOODy8R3Hf40nUg0jTRF9zBJp
9x0rns/OQmEisQsDE+sf0yt3BVZ/afn0HnyPLyqhtg2wh97uFS3s3zH7cRUgoBkgSLRA7sUI6Dde
OVgJE8RTjlYKPFEt+gqsXgYMfbdX+fNLy0TjS5qFbX/VPIxBLTAxNihSitHdIThkUIvlKr3Wyeb1
ChjROqwyO5qZyHBQpmJWfiSHjRb/eOKlX0W3j9mGirKdfVRYJ4UjVia+eVnjhVVKJgcKkcK7FvOY
YEz9dT1KfbMDWMIzIC+agTFvWuR4/wjWol9hN2o4S32ppvRQmk1jn4lXpVqwOUB1NP+8/7e2CO8k
EqkkbAvajd2vFj3n4ZMuzVXzdAGppMXOWl3qnXYLz6WL/eXqAsFJ7HQOn2TNoPxxPuVOSXTytgwz
9ha5euURZXXtS/cF5qElewQlENnX9oo5tOCmx9SsBTARBXYE4O2sXMQeO8Kjs3GUgR+ZQxK/n7Y6
0jHHPtxZj63e7vjDpcq1+zVxOiGLj3gObX15mQCJLn17NTOVPf38MZtqkws8cGdy2iwTzvp3Zhc1
3kl+3AV8refi5u40t6tvGFft3MkjGv34jjMJPEaPl7B2BzNznGublCaYfAb67FiUHQvBmzH02D9v
7Wr1qYQtm1gt2nYWf8ppLIwOaTPliCb/pwJn7c1RSnj9BehGQ2EYsQCH68zs8XDZS3/9gjjJXUh5
ONHotyxENBR24nCzAI3oNfRxpXXD7FAn6M5LZM3LEUO2OpOu3LBy5/CtSiCZ1UpwGP0tyxAf7w2l
z+9t1LXksYElo+Mu651KNUH+2EJ7luiAgviis1JAJI1Jvzb6lrV4HWOMJYqyqc3eZvxCw4Xz2Kat
kLiKnwwGqB9/6+zs0X5PL74SGJpH60mOMEKj39eyuRC+0+1K4m+bYieqO7SCNmN+OFA/5Yig/emM
6NelVOCcXLGEWcfbCJApHvso9/LnpdrEA+dqRk8/kAr5/jw4cLQxXKT+GO3v/Fv3613ixcILLANW
9v+L31EGPRR839reFJomZKHMEdILV1D3APKVBpRwBhmEhZ1h1WJWmE74k4F8FJvRwkGS7EqFbPnp
Iv1v64MLrieKeXZDf3bAszC68YJGi4iTHbUE/577ckjyccB9DLdiD/zkYUVywbcfw16HQItYejOG
053/vj9IhOQlgJXn5rbZOo7fymB1jDer9HmbT+nfQD6TpxCk/tNy5VueJXGdvBr9SAJHqV3WPUFi
vVmqGinF7cbgcZspXvRPxyoF5BbFAQ4TDU9rNRi2ZaTwTshDoezQDqwXv3bWzQTCqj/4Y9NUlrOQ
ve9kgnc3q7MrOvRCufLvhv6+IANGBP4I7+hpKkJOuwkXpG0hzbJg4nwFDZHDE6wN+EtHEMI0uuQG
sF2t6fKjl7Yy+4wbFB2ZNK9nDB9KOeYeci+lKI3s8Tcda76vtEoCbxulik/CwBtK33fSvyBcaWd0
038manf3/Qpruj/OIwC+4xnu0sp4FP2ssBv94eC7+8sC5+F5j8QjoCo6VJUoCXeAUXp/Nq6yugC7
cJVNCFAvCmn/mHqbTvdY2il2Swbxpqv3NOKv1PnymPCpL5RZxRIGrll6Lz03s9PZtHht1jfRpZvA
zKUagebYLpfu1A6FtCaUnGL3yLYPb+wriA2kDSSFN5RK9I7xCfwTsi2gC+77Am15QNJxjW5BpEvU
XQNIs3Y9TdPU/7k1UpueKr+WH4CpZAseBJFLHLa39Ep+wzjUrzFvMf+O0EoTPSlKYjxeXtqKkBij
sK7OnzmAtyqDeb3zCW7izcoHR7GQWcHQhuD3JmPIXxRBN65Ao91raTEMttXEnXhT+2ALwyg/7OlQ
pjsc/XOtjX8yXa125kc77DYBJp95w4UXoTG/SYG3A6gJrdw5xzM22ZvLuo9Iu2hoh/9R/YTxfoWm
Mv2kACzncC2PpVavjtBOzPpb9AglGTwyTmy2axdcJ2SZyixgDNJIjNZijfMJHqijrJwa6mc7BaxA
wAJCnLTjRKRq307ge6Ses0kT65k8bLnxo/+ZVJbxAfHTR2bg1m2/EGPTUTcGqXPZzujjuCXPZp1x
bcNn7aJjH/IDqNODHq/uOPUtfGV18qUGFxyez2toR6bKkjF/CBFU9G0yIbpRhcwnbgKpGENL+Aoj
oPTk48UdUYhZWtYGxV4b4MXwxWxjlU3EGnIx19bw7Fz96aJwirkYm76tXpm4gTyA803cfAuUbdiG
eAj2ru4/tw06ORUEo2JMoXGDupek1GfTGyYhhlGMXQ6v3xAfeW1YK8ZPuS4/2+0Pu5Pdj267R6LI
Nml5gWPEcu+jZ/5F+ALdcbGE6e9cezNhyCgZlW43TSul/+s5HvFehUBEPa8+wilyRMNQk2WpNloD
unD4z5hLxntwSZarfMQKSCcsipU3QLg5/O8QVSEP7FHhEBxsRtbAK1LWGI4Y8C7apUU/dUMdG/Z1
WiMjHCBtQGe5DUmgFk1W4drnHjUiBsagtNlOgrEy6IIpXYiigcID/p/8G/URCuGc9C2ZAR3SUHSu
2BaPOfSvLQqqfdEJdvEA76dFjL0Au+dvPsD0R40bYskIHMwsksGj5l6N9B1dkrgLZEwV+PQcXmes
zDQwTSvhC6LRkoQbBnO5YMhJMHJpgYWk0gdZYyiZEG323F4nkRjD+m5jDKrMNasZ3a+Tp62oQERh
7/V/OVZTgMCXDg2alxbFjalwRJEtPMmtiX1nPKAqvzKBVtelIJ0dGiy3K38hz+rMywNH9qxb+HRN
lpy3eDxi6o57W+aoUXamZKMNlNTyqVXqVC7LQgLrDUq16wSdIQFvSiSxVBcIGcUOmaQbaNN1BviK
PchwGDKte8KrcvJTUZFv5HtrPyBfWl4rmqBYtZKWJcGysExRqBMh1TEHgiLmwmhhUPcqwdVyaj6a
Osh0tu3/l6GY2DwPO8VGurGXWncC1OD0U3mq7vMUkNb0xf5fRtPxREg2Nz0GKegxG2lS/vzqDMis
W7haab3Jf+lM3d22SJQq6y60Klj5XeD8kuUvxnRCIGkv6jOOtxl+ZhMomrV1QELoKnFvim9+ToJw
uhIndJRHXNcZHPJVDuOAlBBCWO0EbZOeL2yVB37anI4VFlDJl/rHmn5q7JBwjnKPxHR9q8/KIrQu
Q/HnFIJIMtwwZCU+obmBsk+ZU2OH3DnrAeHRFloimTEkj59sFJNhDExnc88wC4PpPzF+1psQr7Am
vwpuqUvBSv+wIHcCY1sU+s4FQxNLCzzbCXmhIz3o//jWhz22z0NzPbJmFiAUndqQZ+FqzO3aaTc0
aygGLTEcUiPbNwBE6YDZUSk+wZCkDOfedRzV/7pxIVuWxBJyIYWlWLAFSXhAWxDKFK/bhgxgfSqR
vCaO/qdPVCq7oykXVv5oI7r14eUvkwQyQLCmuuRv0pmCx6RXzFpeEeryP+lNeisLFfvaJEzu5yH8
Z2Ib+yOktocDx3LmLQtqL0jMIk1HRsNur92vtoaGMsuRzWXoHdRQkryp96ZESQuILKhkEmQdSJBc
tKSKE7J264U+elBDa7XX9Ko7dnniWinfiTZ+JoAMrRG3ewmZkk5CanqENPjrFmCAxj9yubQ7mhar
8t73nrVH/nLNw71HDyNgiiQl89Be3Qit/Xj57sJp7HTndPXULrqZxKEQvGa5IOi+lg9pbM1qdx6C
/8JC2UFpb/ksskrTaptG2wfrHsXMXqj6XospUVnJgrwAU+mQRX+XPfRiiGeMC6LYJwAweboRVhqu
A4MitueN2k6SlQnW9xE8e5UnO8tks2Skorm3rdEGcu27MPQb7MAjrCsvYhax9OFk1JanAUc3HmQM
tCtd1LRI1eLVcVG84SwAmQW4nhE0yEZAmYrWq+AicdAUP/R7RzEtUubFss9eT8iOz/27MXsFpn4G
lBkzSGV2gVJKlCnfCu+JRaV5kD1hMo1YRfcD4dVIrPAERkiNMUWoGX1O/K0SoczcqcOeLJDAjz6T
A5np39s5qlidT3BH0ertRBvcHaHSSKQEc1Z2DypEFb2PibXBzATOpORNjF+zXh3d5nQ3YqKV1KLY
wdM09/NUFbYBdnB/0SR7dilXL66EMEizokCj7ryDV/5v5K/VNMo6yrcV+D/SyDvgLhPiRhhkgozu
IAR6BevkJkpuom5enmiGFUpUPHWosExmPVphG3eQlWQHOyN6IqNqh+Ti/wZRQUQveOtD8MHBQyWg
EQWvXCEMs7tcFGJcG7J15IFinS4sRLdRVnJ+VDvHvZc6zeTR3Tw7jHKIC/HUQTxnWdO6J18e4pBf
2mxRXa10vyCKO+aInf8GoIoZNpZLrtXFgHWBGNpZMRnQjBe7yN1Cdk1KOM3VGsSssEiCvWPkCDD+
7qdKtz0mdYPhmqgLU2VfImBv9WYiOUSqURwsepi2j+2nNHIIrgwZHyKyShtTP34GY7pjhxxTzcAN
pb07QOflWNWNFLCenO/Wq+q8Hus1qgwL83p0qrV0m6IS4iyMF3VsyRxWSeze8mUU5JJDbazWyh6U
1sVbCiZcDW8seFRhlAOvH6weEVbSrCVYUjVrHI9nAZX99+K8R3gy8hSSmS1VVNEQU4m+Hn3OYKl1
fblyjT6ojV6+0XAUbx7iapwGTCQe37R7l6uuM+IMLsDj/+kdWsYJfvStVyzlphaptgydsUluEtcs
JetJcKREDfSWoGuEl/+IO4EFNtcl8vwE9DC+8ujYp35T5J2BHle4Msg8jaAsn8M/hIcilUBRN61/
EnRcfz7rHnoJV/++7tTWvY1lB08G7/UKNiVETDC77Uud3BqwMN1mqWfAV39yjjxee3jlw/lGOU0M
ylEjIkhgkO02JTM+REVub4vIY8Sa0eL+/pERPP7TXF8dUfUl8HDOxNmYCFVLglqYTdYKVqiXF/aN
2JrbmZh7dcI+rg/xolqYOTFwIiR6nGptEkMhBn+ST5ycjuRTsX3gP06yk1ARJZHd4QHJFW/qS3YW
NWaErIu/G1PEfHMEtOMTy7I3cbZ83fthMpqgzqYc52se/CKXa2IFYjP8mcg5AOk9yuXh9e0bzCa2
MN7TzQ2kC51P1poUtSz/AK6EnPmJWUO60TzePeDktgN/QL330v6YqAS9I/si+Rq6RjzHUmnKx24V
dwqTB4l23SqJE9QGjsSGkXkkZlk58m0iHsrnbyg1AJGTSWU37wtD9rb47baCUg4QY2jMIgZ/nch5
FITZeEeJAtfepu3tBQqiGaW7+FGcPcaniSaphr6IkWiBxloc/dFP1Dumpg0hvWUfZz4izQw5+P4P
Oe6xTTxJ7Zj2qzMngyLZ0s6YO3ZT1S68vu9By9CC9FGn18E+/PpLYWj1Z7JTrCwHkssW1Mars5sq
QoFgHynzOAx0RAfKJIq/FDsVXR3tl0ASbkSv78MyKHeG/V1PV/uQ7bQDL3kc3ym13rOOUFJHfMKA
mZk/3g0twpUEoWQt2WWKa7DFzm1OWKNUrcbDBTpe+uUSo5XTvrT7/mgU7TEN3jPDYdkNILh0vCvM
pRTk6vs+EbrOtnFCV80hig+7oHIgne3h36rm1VI+NzcdE53Ba4jF+gq+3LasvZD681s4pgQLDDZu
eMACSVR1fnXtrrZwcYOtt6AA30EykT4pVt5wK3R69DBJ7NJ/CP8bIDEKiBkBUmuFmonJWeAFNTNu
8uzt2eFA3a2kH2V7PBUsXFmzugW4gYbkkCNvZobFlXwFehgsjZTAPs4+UwXxtpRW/kP+nkjY6Z/Y
zhAV68pLVdwj4JPATayIyM9XXKWNnqKkvhdq38nOOHxSPc/0qMGDN2VNULiyN1OjG/udTt5m+5Fo
LpFt9XNhGEu84bPoMQTaL1LeddgF3iGl/TiUFWCU2E9/pCjd+9F1J38Pwgbu9XoJqlJjUY9jgC4H
cKRv0VbqmeXCQtkrw/X+MH3/QmQx5ougb5fBr+5IF5vROCO2ixxfpVmBumFy6xwRdAghp13jGim9
pUEu0ENyXxc961jTxhbLyaxcCLsyK9OO3RBw9FkhBjG0NYDV+4Pv5jvvWJRevIbnvhfp8yd7Dr7o
BysdSaSyGl72nWmmszpeG3U5tN2o2Hd+zDlUG2rvEGK4xQjqdDcs1o6pdbxT6Wp36yBLYNAGutRz
nYMvxENL9jr9SumHX8kAGGBgSbENMGMRJalC5wWd6Qz4kNhop7XsFJwACmNASIz4SCN622ICuWQX
axmlmj7HGiL17soU44SDRAN8s4Oddvh2PtX9npwo0WW6mPbEN8VHYl3Cz5zh6z8TaqzmoKOaOWwC
piedB6qtYHDYw0QuWEHBVGFxKc+5DHBtiaocCEyn6810pCa/CV/kgJpKvFJo+/O+CURv8WdHIqKC
BRXHTnOZLdsUg+YxJlApNcc4HwsCWOLNC7ZgPikyzjxUhaeaWLZQrW3BkxLB6SvmaqXMZ4Ox9h9Q
XXS6d1lODsRiqDcl8tCEjaz3rVU1lK/VnrFSAw+40kkbPxKXtkoofQ3Ek3Ym9wd3c9KsMQ3qAAyd
ilnL9k1bBShawATnqrpk13A9lD8YF66Pdpps1XbHiso2wf11bhVoY9hvQ/WgcPfkLp4aZlVlYbNF
/bKYt7DvXzwsHzCE8lryBYobYLAANX0WmBD5COWCjOUZziqmELAY01LbfB8/g41gQpiuG4P64jZV
f8x5E/RbnKIEDqVuQwi9Anw2JrQgf0OAQsvIw2l6x36UxgnYFDoTGbF9/YfdIpkya1Ks0T71LkDp
zHmHtCN9HSM6TXns1KF/Y+fKmYuAwFAlIoy3UCQD/FFVNohynN/rF/3e+mlAHM1LXfRIjNGf563Q
g6pygLGCEavWFR0Y9bnZQeq1Tt2B2ERN0tOOw+cYFSDeTErvlFms1k/ayHG5OPAJRgTBQodxuXQp
KrKtCHQT0OpRUHCaZB+HxEY23nF17eBDKQdUL8d4qTsBEy5CQm/rLa3Tsu69RzGnF0z0Nrh6uvlZ
PKb149gPgXOWqXIggKJNVDwFDxNwyUtuPqSoCLqsCTkIEhvRUeVJe6skFFpTlUN7bdUoXlHlN1x5
PXDDMO+Nz0uGJ4BYymyrtjE7lvePzBY3Xg51dI2EMuK9pKMbXfGTZjnv/j7yG6it8/xn+4QDvGnv
vUjfjl3P98cgj3DyaCC36Q9cFDvT+s2Ymc6egOMeH9fhFFWF6UpxRmLlr6JEMdfBH25CTPcySrH5
vG5kmjty/KBnBITgOTyhkqBkFFzqX1aqh0MA8MriXXwT00+i7KPZRLgo0bbJ+zyy8N1lY+WkfaQb
FmxdJRwVszC5fD0/i1fnbhdKxTU2uuUg40y3RF1/U6empBqjEXhpqzA7ZnRbJzg5E3zWAA1Wzwrh
PYKQmvdQrcvO9nTqMRD124YDRS2vzHHgDft9bckeGz0ugxu1y9p0htxox9IJ84kClAdGPGDg0B9k
u4+crjlbfHms2CfBTyPdopjf8fVBF7868GUrXCqb6p3t2VFYkvXn9m39sG3au+tz4lbdeoLeX3q8
2vWO5ZEzQv2Roueb+BTJBQoWfpggFnczPgJaA9Ur8ktAdeORr3nkrAmxxjiss0zu0bXbb/pdHZPb
D6llNJ1Gv1K6f+Q4GR5OX7py5ieuY0SyKnm2NyFRuzBpsWZkhU926y8LSQ4A9/S1om5mENnlSbQ9
j8OfIQiY3Og4AYLO7F0XFa8/B8aDfUah2fcWjW/Z0p5w3lfJ6I8jS8FaYw51FYfbGVC9h9d8y0ib
HowpQ0qkeapFaL6f6gncTvXW5g39zncNYJxdDONIf5v0+PmhpQCtzwdn2L22rsrm9hYQTmQnK1KP
kFQSQwWDwde6xbIxY1jrPp3fF2SKtcwOTW3V2DkHOqOg2bVIOn5Tut0ozYD6Y01RFfl08uAdn7YE
24rvK0GBmJIeAb+uIoE5PdTq6Of/wEQNKbFpK2nPGMkFlGGPFrwURSSgT7bFSsLtTBw0+hliaPpS
gf3OWcAaq4cxvvtHgKrv4yygEA222CJQdwGhjzsCKY1PHUn6oSknswpORDfbpsiYnMgruwFIpgtU
tCFOUFuuvumap8d2Zwqt4uFJdmt9Q0og5RFWB+i8FY3NTz0Ih0nfYcjQUA8stDiLEuMWvYdFfy7K
ERKm/TrP1YW32s0S/iP7sV9LDSt498S8ifeZcmMIZyisbhSSeN6uy29lVXq9ghpLzTeVejPUpLMw
Xi30HqhFNO5PB/BpjhmzycQ9dFQVQdo0pPUrJ5a7g/mLzM3vm9UHFQ5mVYNHHZhzIYoLDmM64Rye
vPYOVGptOykT8m/AExcvKORwsP3hSYgrS+iJdTt9YrmYEUPgaTlxGbsMDY34q91jUBT6uxulYcyq
DkrWLGybX/+GpFNf5n6ihqdjOlkQo4msZv4897p1FaomZmiByr1Zl/HAjPRnUXeFUWUVf96nGBYM
bybAqwNidqb3nbjifbRj6UOlxd43WQy5YcXr8xhDZbaqEShY1fmr92q3XLLY+4Hz21bEzmqzLj9o
4u4HlxdIrOleElU6gM2yjT9Weve4GMPSFp3s3qPUbZx0haaXnRvcv26dv1TlF9Vpp9SggiIFeDxU
z/is1ux2ji7wr2Z9QwYQyBaVfl7tNiUbQFM3woZV0tDvtNI2ER8DJupG4a5J7lOhaIX7CsJcXk8o
zD10skmmCxX+saxmVtk3Qv29sQNr3ai0+97X+DTXtIe6Y1slMI3KYGxZ82Iio4PQ3Vt33kcOUowW
qrmewM2ys5NWU0VUPnmVeVnHbEaSwWhzobSaU7v7LxgR1vrm8VwmsaKKjxrqNuJSwLwuT7qmTV/f
3iuxfel9OKorfgur5xs9z7QftfmAnB7HOmnP62hUyA0hGbfhzDJ7Soq3grMlQwzNfwh6asPGMN3J
kwzGlutcpYauhEN5TE+zHQqPlWvCMJTGF78Pzqp+PFwkg73+zSLcaJC82Z4gMQLPQpM/isMK9Xm8
sCogu7Lw9EqD7RdbM8l9sGTaJtShV1SmX5SXDY+KQEH3OwTKeQWq+O6Ec4bEvW5ETwHiXOvnaHZt
awJyZoWaQO0Xi4LrhdqtQr7cfGbe9gxAotGEdFjMGu7w3oreUaeRtOIM0mqMfphaor7P860PBrpk
VthccqHpQ0chfiIX5J0vL5Fr3sDipVFtbEeaRq1MeB6dYke6r3qdOmipnSWUDKNqSiZckGl5kWEc
/ZKK+DHvlISO9j9rcJGDA1nLcgM5tnMOGGQvWyoZsxHRNmGYEsutTXbcE0o/ctMLkgUTmuNSUvdb
51nu0TwMeYwiUOxWBMH7fil2Cf5MDrTrX8IhoOvLD0nhezd9/3Nc5H5mHdQLhRcRbj4MrZtDK2w6
0MCcibYJGbtQkm+b/vLzw9hka3t88zRvMm3C/yxOqsiqFZO6/9GSlSzmgJEQsgjANuj/dwqFhN0o
r+w++MOXKsDuKXe/pcnbwzwgS0PlwJ02NQhlR9AaZwhwXzvJymXVaZJrCXHhPc8+mXMKjGuLzWZN
FGv3vRKqsWCBdW7mKXWOWzNazgMf0xEVFN6DsOB1ceFamY6Bp89P5Vg5CREhcdfMDzoXMb/j0RZa
9NQcgRJq7FXXeSD2c1YkCZLIDX7eFzaDahb5x9ykRkbzbPefyPUe8JGOaZSu7+A/jq6hLZXYPsJ5
tS1jiRtaaEovhvFZ+DOE3s9yHW5f7+vt0nIibX8NHkwLln7uqy/8HN056Wwl8lFayFyECc+CUPid
AL8lPBODL2DiAOcbHq2BBBZjcZLj43/ib1BtBG78W52X5DGUbOrvQJKui71ACSC0qp+jf/+DzPA7
nktPWU5/jAjgwlikAdPMs34uzPrLW4VXT4bx4YUYJkoFYrWd3nhSC/qawUEmtuG17R+gwvPfDhJZ
ZwsA9R7oJL3IC7/wMkA+htVPyIruclNGyDWxiZoy/K0/F0lMTXtdniHgPf+Vh9+XzGhOG07B2Uv6
mpCt4LG4YX1Y8Tp8F92GOdeAavrtQ//bjmFEmXdYU4XGgzpXnf25/EgCjt8E9lSoCUGp4f3SSH9a
yTGgTfzGNM09Cq/V7hhQH7qUxrhQ8yo2jWtHYhC4qLePsbKf/w0cIJ3qg8PIxa7/89eL13+ZK/qn
qLN5ufR3dAfuT8hZGtPZ5GiOnkHi1rLPQtpsQBZCVDZZ2be1eEltYL+aOe7o75MBwfIj3DARwTYs
oAtg5lBodekgVn2J4+3jLYGpdepCrQGDX0HXb9tMubcxy+66hishVz6VbymThvBqVA0jixabqQyA
ZhTBxAv/giMe4amyx0ve0d9cMQg3Rsv20A8SqcyJoVVH4cjw+isAzia7lu+wVQpYbDf6uHkT+Q5n
jvZGr5CFp68GE4ChN4v31R9oLQLFIjZ6jwoZrJN/fHcuXDbwqR+aibvYrOGHKDkRyO2ta32VpyWw
DLnMz0dzxmyt+BqMTNXFCcYOLb9Ma2ZtfUDENRJFbZZmA4zJ/pi2modLb0X4pCborkN8BbRH2MOo
lifsGEujXJOFcKXVn2NXte+HSVjJt9X9cDjgBZMKGzaYzSHW4gX4JXS9B0mQB5ma2HKqrXJr1xQS
afwIf3pPoUJp+vqDe9rwAd8k5qHTtTzczq6qrH+d9/6DX9vPtQh/8Ka+LXbzHu22UY0FtQI/T8rS
daiNr2f4xpNhDjlNe1ZS5oRtJyZ4m4YmrjtLMoiYYZrx85Gd25yUxC1vxgZ4O0H3BStlbpR3Zzfj
2sCI77TkrzGl6f28RylfBzPqu1sd545uRiX1RM0IKMo7sllAF4RZvwZ20M2rBPUdz3k2kWiD8dRQ
/vqdmgUSrxqzLcYNP31K5j2vFBzeI0vlYb1ZSnlA+YDepkWU4w1RNiChNHGbfRG7nTeJA4KuS/vJ
7FYO3LGhNfJB9mTR3ECj3/w0ly/y2nhwqLmKGU4BqVR2lNaQGDgPQy7Ls40JflCXxaH8pBOcnGAK
PLCTQKq54NhLdkY+JGFKN9/dneG/OJATJFzsfG1c7zYAImiec2Mldk3lKLZOuCcEKHoGc7frS0dT
n5OqpoVT2RxFzacg59GgFvSla8bthKCSfxabxm4iIBOsxwwqZhWn25DsbvBcxgby7MMhT5aOPAK+
fROQIqs2mgkiUZIk7F07AkRVbJvDoD2F0xM26jq+rojNDTeZX1IZM8Wf72HlMoE3gLJxxLESOC3l
RHyJJic6hhZ1i+p+/okU5+g/9h62YwMU9Rc6cAPEC+YeolQvmej45NxCOL+E6NKLOEes38IDZIvJ
AUXcyqNdHivOqHwae+kVvAO3nzidJA65mjWzLjNh06qlw4Y8cEKqbJyvW7C7EdVRthC6EYx5A8Ri
zPLFbBLUb6SQjiTUElR2RWll9YHyZqf/ggexArI/EW9CYqiFVGH5fabQPdc2zCcwaJntdkYKQbnS
jbPDULN6FnL2ep48UqqeQsMbBVpXYOjlR4Oq+5rD9YddH73NY38lTNHlpnZIw6Fr7F8SlUydYdcE
VcrP2WA3MbNroIIpoNS7XJfKe11LMsQ9FD+fIJlEyfVjHKy4VTy7/X4iDi40KzboKTi5hrRyJISy
aVHNBHQ6HXCaGgJ9+5d3ncLXOaSj433LwnX8ch5sf4q+7Dxf1iCt6gNwCkkno9AxTqU7umFWUQkG
Ii2C7SY++iP+HWP2lEMnQmdiV14USOUHDbc0LpkD8Ym4Dix+byTrEQcLXJ7N+LpkS7Lis7HcuvJm
HSGJosM9wzB2eSlMqfuMgvdeg/BJJqIEPjmSDI6kwryAHd0xLJNH9RpP8hIy9FVuUi7a043s1hcx
mW/8XWxeWUf5MzdhKif0MeJ/4H4HGQc5E1k/tU08kCkjHGVVv8oj4jQu8xjDJ3kt4CSTVrh+Oih+
Znkmsf22BaJi5rSokZm8nXLX+dv0j4ox1mU/ywoAcZ8MUQV+YJXgdkTvF6HhWd9vmk1FtbmSB5Ln
Kiuku0DelItPpQg5+8ZTtfahBPAB1sIDw/qMUtDRbBQqtenGPSWxAg/neiL5JFIBqua3cpqtMPuk
c2rNU6zIr1KZ4zaMPgm3vjyslQ9qYbvp12cwgKG+RPwRKV80aA1yuHs8XKLCNp77cDYi/0tZ04py
zy1yfWd2gLywZHH3jWfBCCVqlWutiRUbwgTG9xyCmpmOB0XWdf6bGRzfbCQWvAQ34rUKuoqsZX3c
2gcxLv82zghFEQUFrlsZitS7c/bveZe/JDFrd37JcpSsaYzr3TnLVZbLXHTpWDqtTWzrBU7OMhvw
EcV8FqQdlcANE1Hvtkku+8Wmv4gjB0H2I+5lpjqjVwsNAPQGen6GbS0n60JgRy9nTRmknQ6CGT+h
ISGnOsgymKc+vNAoCtGB4THht94n0Mm6JK9ePQDcOQyzeDtWfsYZz3TlYvRGzytXVuIvZ+ceTypp
RqAaznzHYQ2+gh2mc/ZHf8ey7QkbsJc6QZVuMnsS+/SvMBtKV2bDarrdVGvsWsP8Eqx1FZynDRaj
lmlkhRNQlNI1rKLR/n7thsL+iwYrLlrvj3lGK2X6B7smh3Uf//oBjnsgeUKn1OUEKtfMD+CXIK/s
BK9y/hgj+B4qnPVsejhBwDi7KlJjTQIRts7pEtuv/YHijAbFO9hOb1mvx+a0ss8bwtmH8FhiI7ML
/OSw/P6jkl+RE3tMPprwlNcVerP9dMfmsRHd7ijpzDe30mTY4yMPyGe7lQvnGXtbFn16dNmDbm1b
HeKEpRQjffn0mDYENlG9P0BSoXFtqH34KfLXwkcG5lTltnHbgyesVL5ACj1fNriHQs/2gX1umiDE
P6oCbg6cZj9rTapOEnYLSEzJIj6c9DfRpRsSgynG8qeVuHHcaw1oic9ac2Rh85i70UDz+AkuhTNi
gYJD6crj0mQAqRblqwmx7idEeE38CbY30OczKvwwlpauA+tpcQSnTx5rSOGWPIqjDaffKZKp+Jr5
YGm8oqQMMerPbvAao0AvKKDv7TXvcSg+CWl1lLeAVX6wzzLRbv2+PTnAxhcuUgoze9kHKX75OQ/Z
A4Tlqx60Qv19HXsHJrLN+mk7upnEKB2Tui1LiaKcnagqPmya9y361UQW+WuLTmEvqSgxJuUt7jUe
j2kKBMvvrjiRl7jF6QIJZtI8jC5lL3vMm8eLUkjOGyETWT3kYFGRR48aeztgio2CcWFdwzXfWDis
mPZAC1rZDQD3FcQXrcpfbInrAHJXg4Pk0nNOU7UKEtRzZLrP9qvlmpdLI7Soh6HQvfax7BZUwJMd
TlR6tdlB2Tu8Xq2I6mYeDeZ2H1FryCIt7CiZ/5WP01l1qnxIOpkAjQbM/NdPmr524li4DoCNX5Ol
bPxx4YX0lsTqWHAdSQJ4hHyFDJmyokXM6dHpkofCCYXenOaQ/NEoDvrzs/49TSXFxKA5b5nSk7n3
P374fXKMV8XNNsuWHMmKqnpOR5Or27ZdgB8CVmqp+oOI8wJBV67XYUNH6dZeQ/NdWU/wjjKmq2uo
iJQkD6fi8x7KvI5fU3fOi5dOLoC8RPgRPbLtVjIMoFECpa6PwPo+LKEtPQ7eowPFwtrVs7Aq1UZ0
awfnOk1rD1+GT+YxVuARPmcwgpVrIZNu+1s1W1Au/bNUHzhe3axi0USNMBUv9gMuboz3jkE/GsrN
Lr0T+V2zRLRqKf0nKnCKUin/5VfmZ1HvlWdcvzTqbNVoTwqmwctZwyVP0/bRVvaq4uE4nf/4pNcV
M1pc13rYxLHtcoBKp0bYAQr55arsTiZdnfEtL/fhLG7jTQkToJkZF8ejWQsni9IetBtvVqnI+Lb0
dQMpP5gNm/WMHJ2VKBOkau5cv7W3b2wdPtFMK7YPk2u9nPjRChWRs/I97okx37dpeZN/kTVDTiVp
WpEHENIYKrvHHti6EkbJ6b5GfFfDfcRu/wyRNmRfAdPG/Jkyrm+qADKn4QnbTKvJsc1SP55bTwLc
xGzV2o6uimNxOfLIUAocM9byFkFhknvdMsso/y0h/9YH1mMicM/Kvoen+cIi7z+DsTV5k/4a5V5B
vsJo3xqFkg0bMjg/cx0Qlg+EAcBDmqq/c7bLgm14OgOVvtZ9MwxAkk8QJ4bLJsHUWW72BQ/RtNqm
uIgssZuAIkkgWKmbEYwEHt1eCJwGgowQoMOg7jHCLFKFwzUn9yNTXD7pQMeV2xgteuJN2+x+B8Tq
Oc2/PL1HXDAQUXIeAHi6FsVRLenrufi/Q4iyoPLzxcxQ424aAoJ62SgElBuz86uuQEGof2hhqfJZ
+rlF6lXMwMav9/6DPx1htC2VLwfZ9Xljr3wXtKU5SBJgCmEleUYx0lO4DhgbtdQdhmkbY94a0ihp
GRjCW0LqBqo/48bqUKGStK1mKs8ViXRqtJFX43iVHUAk9MCOw6tyap3m9XDS38kGmxTy/fAEdHdX
psn0K6q/cwS8cof26P9rKx11KxqYVYztBhUNWSvsonh142E9KtmS6dBHPAosAy/lPYbhobaeCsit
/b1DLNjYWQZTca856jG4uUqrYEL0UZ7i/DaBg9VEugpuKhhJPm132N6LiIjL1tsLkGCDRf1jcNZ7
LqqVjsnRrh1DwAuspLZ7MYJ5kXiWTkbqMW615Lv2X4aK9+sVD2+2UuNSd5LoYPpFpoAdUQo/0yEG
d2z2XWbFKv5QJIAhVIkgnY3/nCWniFqCyKXm04321vgRbnYskBn90ZrQDANs0qOniieeKwOFTh2c
m6rTgAHC0+4/ZTMri+1GXOC0b9MRl7T/i++ooHfZ5HcM8C06ca96/QTQaYuiGm9W0iHY8QExbSmS
CvJe35EYI34goyNpm+1Yi9+13yG/onZcwOUDj74bNEpE/7DC/nRXkhnhNrfhCUfMEG7QR6CuobS6
Q5GByXZaGQrr628PKDcXaTfOn8Sl9qzyljXlCtmg2H66wn73N9WfVDedZwAEa124dNmiOrCatKqY
Cv97XAVr5d2RivhcPFCOJKqnOZ9/vHa/DXMFpk7xx/gHEgaJEcd4rIZxanv8COV0mUqBtHenvdfl
oefMq1qs5vpr2rTvTQI9k2v6da6Crk7Ko2CLS2XmYAQAjpnVauDfU0n3E2Lsw5UXPdxzjoVZTvYj
UJXuTbg3TQrtqMufHEIpk7x62+JkXtcZPxoqR8Tffj18hENfzOJFqX0bbuMXyHj4S7GPkq6c7Ybs
J2m+ReF3NOEBwVx97/xUmaLOzkHef/FKBH01eNA24CWronxYShI7FsYcco4pP3jn7HDL+WiSYnez
i5vJbQhccFiDqNA5r08FtfuJDC+eaPas2jK4i6iNErkyslErkXXFK/zC3jkX8cehPKVH6SkP8t4s
djyCZ4mR+LwPcQWZjzFJOUc+nKlqw/4xzN+BDyi3Fft3tcM4GJe1GjDCyHY2GQj2gsJq64CL+Nr4
IJUx7kMYLRny3h/a29rNV57k2BCIFp5Htdu9Y1BFd86jZbZPudGCVYV0DBuTY8o1+zoF4MtfX2Q0
l+R2Le65+/cXKVJYJJm1mWRhfp0iXfy6MzvlNYPxITpn4a9Joo89a52PQBoy9KWVn30tHk1emkMW
kbjFyrGOz45gBr9pph24qszcL0lHWHbDic8qvsS0MeZyi3907o6OAeN0HEfYkHcNDKh+9mDRrUjQ
RJGt+HLEcvjc8e51ARMDejJT2Rsrbk8rwLLhUrbv49Vy7IYdsJlbRPUfA5lMw0EzRXbGFpgT3XQ8
RzWh5ujjMSzTv9Ds2St2BEzns51EKfB4jnRS4n16oQV3C26KWVAZ3AVCyHrdq2kwWLEHwQ2j+pi3
xXULFGOffh5I2dOpuUbEOJWbZvZvUQeTx1Jb49p6gBNQn8nNr2H00nlvXnWh2+XEsnkGELzr8UCR
rTfkEDB9IAyq8H2xRBrclOLiGhfRMdVjpCTafwS53CN0AM+4T5pWHsb/NPhV9tSdKompzqXNNxCD
ZY7/PWBacGpxaNDUtS/kYDfGedsNRWAiE+lLkS1u59twyMlL0s/9aylLQKgB9F5m6K0RYjcFkqtU
lvdIYPz/70LpQbgykyNhPveWVMC/Ivi7J13N8CfYrhrWSlWHZxMU3GUGlexdClVjH+JNRxFYgfI7
V1vmxtyruOS4zYrm9Bu+kQRYp/wjKDgg1GqS6kPVHGNxwnLR/TrGB0tuuc1z8NCCh25a6ZbBhOFZ
vtEKWicWMAirqnhInYRs6iPwX6pE+K5vfLLMCr+94CD7oW2TWcY5EW2B6AWjrm0A5jCdW1iVjKlB
JWoCIBQtPqpl7RA1zFi5iNVzRIQIFg3JvOknSCCTu//IMKZODPo5BHr7WS8/85M1vLSAweF3rA0t
Rvs/umuU2Iag7NsDRimQRMIbRLboMKoQM3vWQDBBBKlNoprbmZwZLpaLSGutUWlIUzWBdeuWXqRL
t9ZLn4opSH6CzpDmp8L9YHa1APTZNKAAaiSicXoNSsRYMWsQqmzGIp5lHSXj21TDG/mfA6JGjCLO
vtrAElRWxLugdpTOUUoPYWnUmZR/2omNbV4IZCdsRflTFxBagAgGTteQ/aHYjTQ/gBRmhbsYKjhB
H0CzAhuy3wBkNTkSeac5VdYNaz9E/iKZPmGaXhUIN3h6L151VHRDThfiZifIjuB3SYHvFmOKdUFR
mad9bVBSTBbb+PEcw3ZTMiSzuOjr6EvgI1UjerStzPpfSjIRZALeqwmHaYXt5Lhu2QMCtWCRobiZ
OlMTpyRMWkEme2SmOqCv3wm9iFP4TWm9DpOQx2q14e8YRtnIL6nL8gVmFl1eYnTkodQCInTGcb3L
VrAlX5fILGbcLQ+XZXCQuObjNusC3YX8xZIQjHQyIyJyo0RdNagCOpqpn9uz7Xa5kp+qWfly2aOK
XHrjYoiyDys/8nvlG9o50lNQHqE8pzHA2tL8H/gtYReNAaSDX6j0/Ga7L6rSaDWaFBiij54/WfiS
e/1Ztlsm8kG2k3MS0Tf4gC1ycfq5Y9cFeb7KfNE7185CGuLwp5LvQoVmExE1AeDY7URxJIqMI0Xj
UeL1//KX167sLOnrTNINl8xoSRwID2yQNqWoBV2/SwxVpe49a5qTFrEZRDNlMAwzHSYCz+ZNsoG6
H4OBm8/Z+nhVgyRDV28MrSZLLIO5mIVJL5xkkCNdssol6VOStP7Rw1y16rMCg9YsTUZl7UanZlZP
9a5ZDYq0O1w493/6y3Y3E86FKqpahJoHHXdaX2J9IJfEHF3vzM7pXpJNl89b5r6pktAS/e+i6VOJ
ethKu1bqf68n9Y9cZYcmecKo6Qlbg1efXYYbh9nIWBNX0JZhLHNRt3OM9INMK1ghrQBS8q04E56R
6lij7iK+tXyJjVLGeeIyUIVbji3XbFyDqCoZV59YXbgKF7olqv6HtWhRGywP2wYRf5ugLSjpCA6b
MjnR8Ts4yBXO+pa9CvTxaES9T6iy65T7mdhC6r+x69qnikCr5ycYPL58d2uY3L8A+AeodLeq1nCN
OZGVuKDtCPUQAAEidcmjbXYLT0uVJD/b05uIFMvc9Ho9OtW7MfEsWZI8BQVJHf9paj/X+KPm7Mqn
pLnJzUcgVBBys12MHCA7kai+XfM1Dz/sSwFJBBwPap3t7C8Vf2Aq+m4SsM2kcPnQAQlMouKuBEkr
hFy6j7xHD0widoiqXiCEB/GUi6GRq3BTReZ5MpvGxTCgDiu0ewaToF3pTBFJwguI+7cPFyYK+4pL
ooTxHXg73i9j55EdFD6UdzxcVk1H148XXT1QweHmiq+AfcyI3VxF7Eb8FXU4EhSl602MHmkOavj3
bfEGKr7TaAayr3sK2MjybJet5N5WYQa+JjjI0B+SX02DcVwrnvw5qY1f+jK2ZgA4q0WJLRo2wxGj
/cV5V015ebNXJ4f+x4bkNx19rX7ltxUsQRoITKW92ve4KOyHo679Urgkuu4q38AS2nXjmCoI8JJ3
z8kroZmd5mN4IqDxrHfJDcbGa5zorAqQZ0pRW7NyCzmr9gYvBjryJpbRHHbX3+LMRvma/t/mEsMp
SLhoYKBeIdBNvjqrje3X0HjIzJ740OHUp39xdkk+FaqpDRTJGaQ4vOkW3DCQRY15N9xERTzqA0+S
voq8lm43IbFpTLEWPNTayor7wXmlNnt0EF2N0NboA+7zZ/UTxSbC70uFwpB59KZPRV7mR8Yj+ait
MnkiGTFJYrJyaOx9z9VaoST9BHhx5u2MelQWIevkkm9IASWqF9W4wnvrT6Vnb79etG0b34UWjek9
etKuhzrSnW9ccQmmh0/EwDhiHlEaGK2htjSAmfU8cRscw50trhCgSZgB/R6zYIONRYJrsMGw8jgG
F8EoAZAXG95czV4NMb10zr+/OEDfihUET5SoaLphybUAQbGq0B6HF16eegjde6Th+G4QROfUZjO+
C2h5d3se6o6khdC26TfGsB8Ho6RtkuvhEaL8KjEvAXMIbQUf6nol5+JdEce+kCPZ1yXTSFUFNxvo
hH2LGdOdl28R9bdDH/86kNDbdAzeEq/L/AK1xTktcLlfXV2O7Dv83/9eBAmVUW2ZhCa0rS/RBcKi
qoOP0l+FjlyNXAVF6t8fPFhKrn2vjn/SWSSQZvo/Ynph10LeN+w8p59mNcqyyBUD+AzrZHTvGbx8
v4jBDis86iiG7f0JATo2UV+hMJwxfWUrEqrJ2+EKmyLpg6A3cQzxdvDyV6i+7kW1EcVvl0O3Ate5
V82LDSjPC8uVJUXooqDXoPfNX9N9Q/YWAXdOZL0GD3LZbzZZlEZ6tbMD8qmBSqEdIjtdIXhRAD4I
1qWYhmZaQ0DZFJt9VUw0DuqHojYRkmSJicnCnlQxU9bq+l+Te1asp7Wtvtc5s0BxSIB2TIY4RdFQ
sdcoylfJ2OVY2pjmtzdLPRNdxxUJHCKkaGU1P/uKWu8SSy8RnUESq8/IHikp/LC1lroUG3nYIOUh
5UOhvVWsZhwyY9hNFBE36MIXaP87/kuKNOJu6eiRCLqqTuuLujj1x410D+PZCvdWbJwGmtSQCVDh
2irZKMdIL+IqQf7aA4OquDBulGRqTv/sWakaWZfdBAAgHuoEPi5UvuxS+fcDaOx3s3bOPxvW8Z5C
FTsVB4/LBalARlLN2C0/9rb0wWzaYmlsfLzu+mSeCng4yBIEFcicyaCrRCS00qM7zbOMPKFp0ZDE
JbFkMuG5zeT+qxjcCIcHfG1xrIVOzosS3nPat5arGoWaQcF+adhV8jfi8sH0ED+JK2AEWaBFN8gr
1IbStbRY8ZuLhSa4r5wq4Cmnsi4zbruOBNPiyWuTZSIInPjQcbaMj3yfTHYMNZO8kZsaw3PqWzgT
AVnoKttDlMwazGbneed7H3ihYKF+nY20eGT4L+LMeM3mMD9u+VoGVSzhV55W9JWJAiy9uxzDHeXG
UU3g/3RCulpMo6z97DM5/6B/Nb0GM6G7d6DRQebP1osi/yuf2YJPtVwQPA0CYKVpSX3daZIv/tbz
vez2t+NthkZk6wCAxxsSo7Ok88P9ZBKTyw3GhIpvsyJcLZtw6ZkhdD25IwqzMkxe1/hPQ12y3Wnp
PHGkyck+zQLdPAaLcug12AvFV0gig7z9L+H+7OCAeooZzyvNVxNbkxTSV5kneIMxVo4J4gSk9amF
BKlhVkvn9S6abbFkbtrv3uehgDBkkV4WZhxMnASkZALQIwmvd+yUXlBSORVaRujl1Gp8IrO3zlwz
kn2gCDwK1JsZtlq0+vi7z4dzmPB16nxLMj0M2TC+AGPWSl0Ui5qAR6DmugyF9iuM/AEjoTCB3Bz3
MlZOlMvXifeKuSsXm3OKiJR7kKKHRjqR2/QynFqL31xuhVvCyDkdReyNPme1i+fhJa5HZx3Cclzk
RAPPvfxJEf3PbLrqQeDZgRCFvwnq9PzjZ70o4klmpUS1jHHqLlI8tLg8v6zAlNMd0Y6YHPY5bYLV
tA72qgty8Co5Z5yKsMt6NKIqOhzgYN9YaMQBJgeRHUnRpvvKKHxFsNFZzR69awGam8i/f6CSQjAW
KiMqCGzzJsJVCWpN/gtBqvH08knsvZomxsumfn9xwseCCmQpblen+0BiMSSvNiH3FgAOt/a+Q8gX
TannAMn+4jd5JpiaF6sYgNNKWp/pQMwZqGMiXZLrDJlCqtH1Fe9ignZspD0JIW/TsMtQ4sKOYBWi
CRgrBJAinGsFQqjzxD9WkSaw1gkybNi1cz/CJqkIMmS9Rlp0S0wSeCgckOAap8TWcUeXouCso0jy
HLtN/+vL03yTKzwH66+OgGSHdRvPCb3LgYTLtswUoSyFPi0UeDijpte/QLfSnrVffa91BEg4k3gL
RcEKJTHVbvZPaY3PSZ49ojzTKpNzfCesUzpBIBsTl4ANqjTRHgmXdmXI5pr6SFCTuxv4AmpTp4i3
VC7Lxt6dQP3A8sDLEsOWQj+3TI/fAHQHkmNzvP9AP+vQMHaEMlqvOXCRcnfgeOI++btz6j9ZWYSd
8f2vZVfr67KWunz92Zz6HJjqVvtSQlmE2Ig93I6L8Ql1Q76qH+PmQ+PM4dMn7D8L2FlO52yYUoz2
J/OVVKPvnbfZFdrTh6B2+IMvC+u0nVs6OT+IglxAzjrRIpS1LhiU6bs6qOtbLzhBTJ5urF0XW4pF
Nf/TwFkFbAioMCgmWSa3UPasHEgtvtIY1CsfXa81AgBUth7WcuokVpDJJS9mV/dFEwVelYOp/w7p
idH+p/eBcNNng3+UnNd+13FPNmG0/7IZu/Q4xUKBWEWPdW1vUz8TrcDF7aSknHvJAopuxF8KO8pP
0zF6s27JOaf+DMZwrmvIS6K1Sj22Bm2DzGV6sPGRjV2CLpkUfBotuk4sXZjHn3ohZLrxL7MqWmhT
dYuCanWu6Cq8smLCynFtO/CUygDBf4ELow2mdfm1cOlLUZf6KVvIv0N+HqIXbhK4pcJJVv+O2MTE
T9NhzLlU2iPZ58nkezCI5DW7aUVhtsv+fokHpAVk0FwdjdDapEyPRzizWHGhqDPfo7a3tJAi3nYg
ObUiHupLVYs5ZZSMTeivlgih8o4+KHVweWS1dbd/Ea5KUUBkx/sQcHqa99/DNmM1ul820dXIlCfT
ccPXwzoIJUuTMA7X64c5y2cd9bjLA62SlVXPFLX7TIAiOf7py79zXcJjaAXN51CmfFXoS5PjelNn
Ed/3Ryp2u869QPCn013aG+urWCXHhd4ux1nGW9xhrBKloe+AccVoH9Dvjs74/3P8ojF0b3gKlVb5
sTRyrRt/9Ap7qyVcA+Vsx7SEJheBSWVZzYs0Ww9+bJQxBRn7mX+WRzV/NJiqmjSCOD7HRbyxA5+M
Jje42K7Bdq5C2aV77APfjRQjxDl3Z7n/sHYWc5qix7ZtXGXyNM/2H1mTZFv8z5q4FK7MngweqpqL
qMiYvs5e1mOLFvNVyumqjJMn2OISGk7/3BvrsESV3Dz3R533pQzG6R1JHYW44B4F8LJkJTgtXwTo
GHKK2Zj4QNh2CWEcQlfyo6LGAQKKJOlS8wYMwrV3onGAwoAmIxX3VHzPLqO8/qFNpJHScZjkJgEC
FcfjzXfYQISGt4frCwHXY+g36/REoB9iz3DnfyEdWnnxQPskwXguJUYybUosp2P3h5Z4//DNpDve
82xqXUDmLlPJnv44To0HAbRIz9FPSEUg+XMQNTIFcPGiLXnzZ+k45jR4LqbUFuyf8BVZpqR4Dl+I
Sl1Sy3kC8qkKXI40FgnV1mcMJlD0glPBbBUp+/Ua4P7q5IKVuROE56rqZJ9e3lsnMLbm/uVJ+z25
QHdCHk/r0eHt6E5vrRIMvaUtrSRIBzrc97o9JxLHSaVo550LpC6PGwkrc2h9z88ilPvxKTlQZ4Nr
+Ldg3oAZ4VKz99qyQPuXVgdEN7W99gXc9B4kLnBd+hfhhwN2fRCFRwqEwnmPy04Y75TsOU2mnVgH
QPz9vG2zqhDglaDuTBcWRO7mhJCwWRfOZx86Ck2gycQJk4a+k375tUXgCKJzHQ56xB2ACFzZA5X7
QObgM/JtN93tSFDvOLaF5wJyQ/5O4+7so/l4yoM2Fhw0TdGvZ5m2JwJGCfgU2ykqqEr+p7kBxJgm
VeEOg3PraefRvVfiu4DjRSgF+nIuEFgP49ZsdPuaHI4Bn+3NZBY+ky00WXyGx55Ydidkxgl1IJq7
VuduliXdqb/1eqOLmmM98e6TbUT4cFaRP5o9YN9JtsUs/y0rQjvZeDbHVcUfjbJ1hw5uNH0+3Pfj
9/TVGcV8XZXAMk1C3q6jK4GZgmYxl0kqGYiuYgj3d0qN8177z9uvuDQaslvE8xx/8iCYg0d9yN16
VXRNVPw4xDTeTe7iyvA5qnP3SLDgiYwkoVGrEGdSrjomR53gogyEp6f9iu7yO+Jvk08FvJt76QQy
+Qqm3m/tKw26hsQPAmzEyjK/WuJ6D1SNQkiyj2Djm56nTx2Erx9ebU+BeXJDXkpTCGUwF7Wpp4yW
bJ0iW2CA0fA9v1JxGbxC4/aDvQmWVdQxaN86ljWLKNXpeFyHdNgsiUdX2+PK7ivCDUYR/e3KfuNa
JxmXOhPCRbQLW+PibJZ4X4UknJfBTMLuXuYoZg98nfpkeVqgan0HMC7G8RFbOElphnSvZDtPiHio
qV+Frh0+wJf5yKH0HB1nliSCBfwYhOlgwhr3FkYkkvFYOnn5FIRxqGswzdOXxKT/Ka2hzfOlgTLQ
PTwk75X8x7G/8v5oasTDy8I5AJVSWuFoypfEfGbe5/R7/4lsowGwURdGgaDCcoi6JCVci6Djf/4o
zT8j1VYUt68KDw5vBGC66Qnx1TdhM/iHt6fULEaLsq6JRKMIpKbo2QlvgHKLMTAVem7RFABAs59z
4gjJn/Y2OwAnukvkyvbnmhjHKvLadoaOunbNuCC5faeLkYZnhG3u+ejnZKeSNYz5fmV+u9OksWLr
iIbvtS+vBx8OmoT4Dq/QpKjThjHS2f4HudrwcZn+z2yOG7e4OGFV5IMIyBviHBi/OxM/FC57T5PX
JgQQcOj+H2LU6T56owHlEXzzSGGCg8vuij4s1mQUvK5GP3ahXrhCupLYcdZuhm2Dy2IZBh6C/utB
tolLiJtEjO56Y7sl950bJj71SEoRf17IxzLSzxTXl6BnFXQ4X9pA4b8nUQNo3TW9+2RcvnR5xk5w
EZhPtR4lfAIrLmQAGsbMSvEwAARvxv8msSrKUmoy6qFbDNkeiv6oQVDIXw7GMMpgVm3c/jYOHtP8
JYg76NYnO7nMLWAkqbKFfba/uQKbvN+5xQvm8MKh3169hcPaWMbwjRcQhGM6L/tiph5CboKMBIGG
4B1A6xrIHha3BScWceT5iCqvYis8VaM/kUEtFuyUjIg5GQsi1M27Ma2eXdnw52QJT+KPp4lVZFF9
loywCOFQdUqnMEZgMFgPxzH5C+j4Tnt9ozJ74gqjy/YusxgQcRGrlplE5R/B6gp+iKSwv7ZWyvB1
KZFfW0oJtK66Qt1QjTxLL68SCi2kC/57OsGcLx30nDwldX6nXRuhtQvM1BpnuWTLPv+coibg73mW
HJSbRZ7CuHeM4OUSfwtR9qGgY5GGUOzFwWFA4mVKtTysc7rg7jOyLnxwVrHzhH6QhU6X5nAYVCeb
qulod0fWz0q8/vPtd2mEzNtvsOifEsnuLsRtneklS3VE30Qe+MR13Ghx+KOiX+muv4p3fj5G6Pol
I1qzmdjUtHNQUWT8G+Y/8OvgD72LCdGUII1oyIC5I0TdVq4nBwIAM+1D/hdNb/QNmtqtc27tZ75a
SgMmGVxjKMIIjITPX6Wusd51MTcpCuQ489GhD3GH4RwQeLPLJPa5NWqtoLyVjlZtDiyrG3ksuqfK
lVBGTWhgpja2+2jLNCh4ZAIhWFNKGrd+S7b6EOG/rpkfUoIYzIP4q5uAfp6lBnlGszh0hnrSMOPH
NyZgjPxo9BjMfpIu0vrbdMbD8u5+Cpoxj/SRDu0qhcyPF7AigDNJU0zYvmN1SxBHJBVh3rdx5toQ
s8ePpxGNwAAQ8mk18NY90ILELjAAOjO0o1PJ76IHN3CiNkUg3txRP0S4RAEB9RT037y5VCnTDyT8
D2ZoFkriID9N+oEIU7ZwOElO0/DZsVsB3ifSKdGx6N3/MOdaAhA++b97H5tdq8d5M5bu2keyMs0K
rGkJzRlQETN+CpAIIglwA80sag1FUZ1js+I+gDl7PxRp+gYfMprHEy6TtDEYV09tkFhQYGMENRTj
asu8LNmwjNdwgZWE8sThh09I8/UZ3A6Iy2VBMQowzksd+oja3HcgseNiaGV5TsrV2N+q5LXAt58N
p1cidTIb+4KcWOg59WWS3AHO418jNB0xDuYqTnolLshMhDZJmKYHD1cTi/6WIS41VXsvGivLNrHt
L/M02yQUyIDLoUwYuGMW4ScjzC641EGSRIFwvZlfvwBdyP709Wa/f+0tL1JczxM2S5OtpUphS1H/
GKONegijf9o9qIGePEEZymyZbx5dJ4Gg/F5BaRWvkdUvOl6y+Cdxvx5txo8y+Y8OV0SW3G7A9R4U
GLopSjEgOTFUPMrqaFtjhGjIy26PNqFGrrZK6af7yBFEnJ5HMisDYx5dFGYASDc6wCBls+ClGS49
kmomLcUVkH4n2zGM1ZVk+nEKLFym06FqC+rIeLiZGeQFU2nNRiDxqsXRvw+6mlkE9q4XSo4DPChW
yF4FZHPv5ogTxXEFeIHFEj0ygY2FIA9Rq7UXC/wUbkwhubJIun5b+nf04c6nH84heI45SFhBMqI/
B6vNduh5IRmSJFnSeHEZDx3zPjUQyQK9TM3+a+xOR9VVVSQBEHfJnnhNC1vL0uKub5z1WI3IrvDX
oJ8SVlH9qJKrDsOTS0qlCD4T2pJOggp02Xs8PsS47K2zTJp7TB3eQFeD4UEn3GawjQXH5HIzRD98
pWEJkpoICiu8SzA0l+qdj9uUFePo5JDamiFjkZxDqiHWuHupYWymdkKf4XVfiRGZrv01loj5ZYEC
UAEOZ7FiQlfwjDIijAntXpmXAUazTKEGmsdwa9RqJbmeOqlQ0NAZVQWwH159rRuWuBgmoy6z64N+
oNAQpIINxM4vYSutIW/jqMw00O0g2sXw/J43qlsu2I5gadAIPRIvgb8oBNRVcyWupCcz/fMIei7n
MO9ZnQBrcZQjIKxQ9jApEb4uf2aIx9PiwZZfpdW7lDzAHhtStvShlht7sZDiQCH4QpbbPkjWm1JB
R8OnL7H/nBDu5xnAT/nWERcqcX3H+jqZYE5ZCOiqDfWW/hHFDHkJXkZuannNcndHpCs4DJFzjPgk
C5Pi/VlM0Y44YcQ4alKz0WNhpC8u7EdhxfkRC2tm5xoJBW7pgUX4q2z8IICfbVIOtPnns+2wC3np
IltKGsfn+MLfPk9qQ53zrdKmaQVtFEH2tpBbu6xnO6QD35AzjoTCkisfEiYmOoIyxbxV6OpEeEfk
E9eQ9JcUoj/AV8BGStOof1Uti6EfS3KIejGsewhs4cyKMrBSd0/IvXY92vCaXSyPev2KEYQ4b3QG
aPuo8uj84Wi/G1DZQ7bT4a79AQjdd/YSujpZdu+/PtNA+oHTOJGa0aD0Vhx/eC3j26hlNVLUSSwI
IDtXHDhjXJDJjJOTfAp8kftouqYih0D1y6ySdnO1hPUW/d5QJF4rRMaVrK53p999QVWIXYtvzqQx
lF02Qcu74tGnpXeNqbAIH1BRZjtdRCzQwejrbu4F9WD1K71D3a+qB5Nz17PxUIQvnP19YYJdiNHJ
+fjWiXEVy2rSUOZbN8SMe6yWBDsNxTL44xsGUMBV93bspRv+hEXOohkQc3yfZedny3xa1+71EUYK
crg1VUQiKtE2nMhTL7imRAuEATpI/C8Mk9LNK/oDTLKGYVKtdv2DaLii4IeoQpoVx0ucv9HVFAcf
gnDH+wlsXakpO9zJY2ZBHNMx+SKPNeYYv9eF/+HT8JjmsFu2cG7JlIiPNY27g5A4B7kAlLQcSnHE
tzUAGHjAOMMW2X5jULKbeNSnnRHaFqXFx+5pDMoFBDyq0w/wfRfxxN3e4ORRG81Tu8vXGDpChtUF
zdpOuYM+c74In1W2itl3cxBOaWdg7Srhstf6wyqHerWAsQjb+lH2GSIBQtexyM0N7rN5+cS18thz
krtioXt3AgHP6xwZ5NDMI1i/aoPOTFy0Rao2WVwlVwJfLrjz40K+f0xG0AucnZ7FQbpMUy/9A1pL
bd7RmOiZbzqfS7ccqR2Zm2o5zlYuSeBQ/qjg0+U0b8NaCTVrwSEimuyUw5rb2wNE06G1XSTrZiwj
HD/9pBNvSPBpHgvFJhyTAfT+lEUhWsr0NYK0L8DXCFsO8jPt9lNge2ylfvqZV+gpfuE1LY2NXmBO
1ez3kAVhH9P9yKuMMp00IGX+nDGUOZE/Dn35tLOauCmUPTuYGw42s8BKp9NcCY3ZDLilYisBmzOU
vnjGGJLf71XkX8+BrMYN5WkEvyTniouDZF6Si+OrYZXClyj7Tcenr6UwhlxnlmGovaM7M323CnVk
tWR/hSKMPky6U9f0N6kaq18kG7pHCjyKZsDyxwOT5mWZ/ikKMZz+caLx2CSvF9oT8x6my1m5iSgU
ecCAfOp8korqYjSZ1x2AFkckXBpDn7TaTG2Iufg5qHuqLQgeqkBguZzgqvSMq/AuoEboNc9KdCWs
nk9r8on9vZATKM8NFeUs1U/JADi54wdZca4i3brXq0BixjRTrRoGy8S8ktjIw/xFdXRBDDjfB+86
q101JlqkFMOwsk28p96a987cK/1kXytrEcCCh35orLckANzIq/o6fNCsjQRa1f6LOxsOvxcFnNfy
C9n0BBahp8E+e4foIoZ28oq0WiJoKWNk9+OxTCw5QFe9ZXfsih/oJobghejoBg19o1lp5x5O3cFV
+TOLuPwvdhOak+kFqP1xISYLcuGDWwSdtROJOcubh3rol80deSNwNCDCmEKToxWVTh0rzJKt4G/Z
AbZYqo1cgYTQOPBgtD3uVWYY2FAVag6yXtLtV7bazjYb1oUArILLimC1AMXdChBmHzasrOQ35II1
qn/UiJGSnymiuQufLfa7GXYipcFrp2DCfbOqoeIoQ262vm+NMl6ABFnklD8JM9pBT8yRg2BcASuj
UIZ+MCc9H3BYKis8PtvD1CGd13fHufI5rZx09R3IQ5a4rH1+oYW7Mi0Mk51wG5jBMjIrD7iWYV8E
V6xunHRiA8+c4WA+/gNNxv8RIRCsywhmREx7en/p5qdjuEXfkhgykTvnEIc+6nvFmF67GA3kqYP7
ddpOl8McXcVMR3kmccM1Uxx8ugzFHx87CwcZDJcbhNeEgjfX6oiWgBHSDcHARFOWeDi3QxOIOB4g
Kb6KWl6Or9QVmWUGh/GuXLekFk3RU5sQIygJyUqn9BG/WPBd48uFWMx8Bdiaacg+J/8g/9NjGayj
lA6Djh+siBMf33a/bvwKJfqgiy1IjbNFa8L2Vw8u49ii8s+rteqqjDTccWJ4X2eGgCMAiK6Ev+Eg
87PhmAC5dJ7RjLwNa3V/ihZ6vphZaLzTPPJLz59FBG5708vLZdu5mVk/fgF9YIgVFODkjHb6XhKK
6ieXSOl3f5XpygCrDUnslso4hIeDzyuAuaLRp0ROH6XVXluNLy9u2IpK/qT23+zSbZSrAUB7MVOJ
EGBERbCagSlEpdwt2m8X0zuqMHXWvMWBQV8ncr+gMvsyWwydboZGHZ0/yqMmnoxSBBoTLmela6y0
wQ/foVz3f89XDuyloCB7GlKvqd3N5qNkhoj97UURIGWoP1Aj3SAotlRnyUEYU7EKIMD4z6uPDBip
YTroMVDuDygUhPXn2/bsWK4OkXjZNHDXDeaXhVUTTyGC8Q4qR3VndyiAgBH9uCBHZcS1nBZAwRjw
jG7viaDrz61cQgj+O+nYj65bn3HQQenYrey0/tB4S8Sca8Kp1RG9QpktXt2XlIBJulHayQKnRk0z
X/9BDwt3/CNsh7ECaJGZtm4yubitSyoaLX3jppcK9VeSzEIyg+APRjBiWJxGu9hzUKTHxR5PgGfg
tftLeO4dTC4ziPBnGCotnPe9fvk5kx/hGAIioI60R4APMK4j/GrxHmym6ZKu1o7rt4u3hCxWPTJG
cQVzGBt1zxzWPyFv2VWOQxtz88QyZYrfNYI8nv18sBJ5TokntnxfJ6JI3wPNiyEYVLqeiZifJaIS
aY4AZzcHSxk1MejJIFdqnoRrl44Ulle4yUfCWyX798AEf3RW+EF/oTZzOcJeWTS4bWADJznuJzhQ
sl3lkW0g+bQek4lhVGN6IBp8UxLa4GrC3bArmEtReX1zF6jl018s/2oYWnry9vVcMTylcb0ez2iH
h11qTMhRRTM63qiY37dJd3PhGqKuGdq3ApHgOkCdtqBZZLuQarwKsKDlRB3cFQfqA28+ZbLV8LTt
nAQo4bcm024FdzRQid3rIhldXb6Ifn0durpL83QyHQkIvEk1DUoptCe2mQxkCxfNYM/YgplyECep
s7XsSBmXdwhjovnkmvXQsw8jo+w81FxubINwB4W9nbeXEqkJxOQeUh2TsNypFbq3qkTqds3eok6R
wHkU7h4TCJDDbqYnOzjxyZiIWJA7tB8b3V+FY4QNFABw49umVQwr44vg0ZY2wLrET0r4/JSRKZaA
zvc0e9YwFRVzFrS5ul22s3zG9avtn9rpvg6YLaGPhPcWy0kvXsmphoZ2QFedBQjurAYoK7r06oIY
5CUj2DKLX7nRPgJJlulTnJ+JioR+MYgljCHNjE+rQrPlbOBkot8P4iej4LL4dH6yeG/p7Bll9Nfk
gF4XVP6LUXIp7AvL/ei6FLOUP0nRI9ISWsJzayHEFL5asUmGhzG6n/b83VW5IxDiR3DN+vbAe9h6
jflj/Q/wAFLPsrlqPracrvVt2UlRWx/dtAHHEpZlomHyv79ue4/pQvboMEafzTkV3lzwwZN2+6uR
y2zoheQ63a2O0oX/nOMM2E93uezurzVFjPreZlme7R9IT+Zu2guwgqYk3sp1jWVKAnehIBiYXMI6
YQXurvMCRMl4tGGh93Da/2btvN4x5bLceA/5wOJpbc3DvTrNlUfkDgAbkfSPv6HnSmV/MtJMUxEy
tt6O2xNSgQoskjQgA1BRz9z6ZP12vEgYVqWC/0yZ0YzjO1WBBKNTTMv30rBffUYaGlHg6Ck0sdZd
wntKnISJYze3iQM5G62FRbWl+DNjMeAed+eU7LGC/eT9t4Vbd4aGGrWUCWQoRSObC0ry091xFwQn
VDQD/Fb38VVuQxBQfiFFzCYj4nIRqB7/SAuFPVk2qbs7NFRx+n+YnWHQjH7c2mcDdF3O9a88Pu3V
TI1/cuf+JC04wZwYCVSeNirCa7x8UVZ/a4A9u0w2CW1pDWwO2vafDt8athzmjAJtWP0Y610t5pey
d2ZYh/deRR/VuYPqEvmvOl4Pj1fMCwl3NjO65H0HJOsZfdM2Je71TC6CC3SR+Eo0M8x/CO+H41li
Wj2jBBviwrUF+EZY8gPt36xXuY8RLe6Wwh08UrW0VUes9V9bJ2AGA8uL+82yvU5Qt3wVBCCD/JCH
KoW2Rc0SCsDw/rU7SYfy5e4zLGeiwEbSJSDyJRKXkLgJ10hoB0/oT93f0FaUHDlDCOU19Nj/iqXl
X1fKIr2fb9ggOMjwdrRz60YDZMkvB7zTmvEdpEc4weGkj/5EPhsLFzwEc3K0aVmSV+MIbO5sTZ79
dZHCBE+qoWs72lS/yXkjClQjA0xIdWNSIey756nnL2REz9oOJTrOflHhL28rezD3PBnwsv3+/oVn
7TRG2mpH6fvqpchnVHGnezpuP07PwnSMGlQV5oB/3VU+2qC3VW19AolnZgyOhVR7zpn26n3lbn7h
o+wpcHV3xCrGqkuP995L7CLUwZT3Trc/4lrekS/iX6V2ata79Y4/VTbuE2lhEQyHreSOx4OMMotx
iLLS++GxWtjcuJx2uo+3Q0szqZptfOn2iU/HtQZitWDi2KL1UUJReytas3RLaCOq7SvdEu6+cLBd
OAU+QK8Lg9th/SzvkE1+LwDrTsl6WmTktBOK6/0H4+nEMRdX7rV7hlXTpPawBIxJcuTkQGLa3eUL
c0KK1PQI9zftkVfnIx6ic+593K7PYxVfh2DcvvoTQO7lVbdaurH6H85mJ05W2gri5ryEYHES/OVN
8j4+OC3o++md6MsWYuOoWbHV+EDS6/ykuphV70bzgVry/l8LCppmgaAOSdDSbNw9xrcw9wlIYYzC
k0Ec7lWh1EEQad7qvMaUCK7IT538TWV9T00p0idMQLOKgzqAxOfO2uBkA8uAWYeQcQ+73U7gTq50
F0/E5bUqLoC41voP/V2g5y1P1tTc3/uj0uAwkU6jiLg0rvuOIqbQfINAWI8K3mE0AwIX0h1j19vY
3zBDKiVo4MMZF1VxjV3rzSPrSsaHI730nNO+i2cp/CWVvXU8RYf9MZ612OF62sEhBtYZ+DMAMvjp
+X16XWJGBpEZxxI3pt7RY0QYWln2UVtduxcZRaA5I0TfDG86994K6mrbj/o1xEoF37pV+vZ/B2mT
CUSIICyXLvYYmkuTUBNQHiBC3TTVVxbNQirDg+wfGSBAmuzlXtdbJTgYdrzSh4fPjnPGzTNoycwh
BKtZceRD6YC7BIRtLZ85NayyxoAlxB/mLmDpdoGbZe37c32XbGJOpoGNA9klTQM3Br7omN0ex2n9
OLSuSMpsAVXYkkoEs7MjDXVUdX/QNeRNrhkwXYyLE+CRg6gJA7me1+kS1SU8zrWjHI+q6eIljBa9
ukbAIUQYh/gM6+Qk3cg23XU7eY3v5vueMFiE9jrFZeHflv3OwqtthemR5+4dHBWvOfj0z3HtTd/H
L+T/zmkOMf3cxGde8cnKAs04h7uaMiRcpEFR10xVRIMRXay2nhghoS/jAVcgsPRHX9C+HVbsXE6C
5QxFUJaz3S2RMJjebIE4wERlhdTwe/4jUNmIAd4FB9iqfcAbWjETp19RoCJCnN1sQh2MJE/eeqab
KCkDvP1mtCh19RsN96Sc7YHraEmL4vKrYoC+1BDX9zKcUfKLD2cumzlFqhxj89lMtYQ0Z/yXn3oV
ZdOXuXITlImHtXawECdl0X08EQh/3hlL2+irlb90F1hJ1I792/0+QUNMfYSux0uX5/0xJUMLyUNi
v0a7TUNMkvpf4/zEs072phJfP4fPKD4NduEDdd+4MtwhAdvlrBAiXYKRWzf9wnoXNCYNpefdDeZm
LleMkifrVTFYSxQovLATkXrZgX2auCYiFYpX2pihOuqfSh8k7XngltEkRL/dRbbN8nQ9qUdGHsZP
NuDDpEFuley2qyvPf3WXe7b2KdvYH3t9oAoiYlHltIdUMd4Ul8KJRJ+yMuQUF52cD5C4lb9V2YD1
bPPAhbE8hPIWlXm78umuZqsfTm0cbRTmnnqJrZeY92+lFklExpVU6Lg84P3CemwKiJvQd/2BwldG
J6Bx+E9N8n22IEfyxo3Kd0/ZnwqkitIWJnE7bPF/HDeqOenzBgMU7rMtiTVKuhWHrKwbceqQM62K
hI1CY/YcwXgX0C5hXR+86tT2UuDxuA0gZUlZimI41r73/djhL6AMFDWqxZP7pBtA03S2HYsEqNFZ
pVMTYHcuUTzRd95UVUei+CcjBaQtPQvS2eDksqBs6dQaw2HrvrORZ18/9E7XOKFXhQNiVFAnY5Ih
DlKd+6PXmdvU6yTb8BDAdSa7J+aLEHOeBFxhHiOUr26bbtROWbRiwrIy3JTQttq+I3/bAVBdorL2
nuK55AavuowJYeojwfI/51UZ+Axt/Hb+Ee7Kp3wSxk7Rmy6x70jk6hxW+UN6NlRVKjsWm6hYQpts
4/TguYn5gsqRBdkUTVOuv3o1xyb1mw9zUN6xe3MkThwisp01axW4VrzcWjgY2nye0XAdOJHYFdps
r2wmbUvLrHsPkZJJsnyvUNu6huQV5voBXL7iODQTruf8Eib8eoWudDKQtx+dMprBJd8w6WTlRpxD
FOBuYJHi5QzQBPhDTX6ge8ioge/eXa0yjx3WhKembdkzwKrtimJrC3D2JI3fHcIfiSjK59D3FGMO
0Muy6Ih6aVOm/xG4Aa8N2zFQ8NfA5MqC59Rd7RQQzRTtBQvi5zuDfOiRebXra4a2hLMs67Xoz08t
5uZrKL4Bu7dX/HU19hLWpIUh9vayrwcuUQ2tch58IxbVAwVVH8JZGarcIp6mzIS3h/EseGYsbqZG
74e05+djZySqHertbUYCLfqh2E6paoHer5HRbGW20pUKuXP5mDu/XkTRWuRL9GvZ+rz+dUDJ3UEo
TVLiaqg+CNBJs+NZnqNORKhR/FZhRI8Hgf9Ia2nvogCXjUp3NtDQoiMWqsDQzJFdLNCKDUJkviEI
j8lSHKbMJWS2bXIRX8PWfobGe44S+ZDgkAz3cYYegbZnLMXRSqI39YgQLGIh4rJgTBtWyN4/JsWr
DI1p0PyIBF2EaEQGyGjMRfjMY3/xLIFDSVHB2GeON5Rs0aur32ndMMP2w/fPeUkaDmtFtEFVrZtW
QKc/DP5jv8L+eUMhbnOtgP57wrlptSwpEt3VEACwFEvAP+00CAUnuBHqE7ZQ78rvpI+/O36+Pvh9
9Z4smWQNRApRtbFkp0cbr+iZ/7ECXSwgE0I52hvezpOpcY9ijXyc5nUCyzUVkhWVM0ndZC/Gce6P
ZiTElPqYEaVym1HVgKnNs04mwnGZhwld0C1ovtdcL8KDrQOeAvyjupSkHWaHEcS4EeJaFNrTvYxk
U/UJB073yb0ZQOVNCpRLXByEXMcHHiV6VR/IKCicXB6QZMZW9EUpDp2soQSt/dIdF+4ptE8vZNK4
KQOVBKpUOiHC+hGmXqYQupS0g6VqDlwW68drKxzlNnuUkf+duVoR8rK7pb08Bpz1PkiQKV5au6/5
jb1URmxzcFgmhP6Odpk2Tg4xCYvud4IJzdIxn4p3+SjIKJO57jrvf08uYA043cs0ijEwj3f0TgYW
eFYKu/bm0z6NQwRHJ7lcLqOPOrvS6PaPi5wcqwff7eKUwBlIYnctMh6oAYP04GfTgKEfvyoAB2KS
vFC6FY7eVfei29kPuUGUlKhqU/JXFM7H72t07VItbnRFOOtW08KGANqP3HI8ZNhMq4/M2+tBGbfZ
83Iyy3mC63TQzERLK8XPjju5nUBHDzx4IVhehdRBvcb04uJY9JJcWoQZri7E6Z602XX4cV8Y+jHi
876bXG7UvGWJW6o8UrzTcejnf7ALbHMJPxFpPx9r5PaBBZnRLdcv9vb1IZOOIKONJyvfJWLjKd4u
9dpoFdwgVm60lsqg1nPH+ih5Egnw6Nrkffek1CH06ibKfNFnIhh91rr488bbLXhwO6eEJeVB4cDF
ZgY7SKstA397mLea9BgVqTlcOkO4YMaUWpxwtJ8Qj5iF6rfgcCGKsmsdkmy2AEgg0HRwLOXq5h5/
UnA+wby3sbAxSKvhAl9UOdUMAu0V9fkaVEpTUeUwaiCBaf5vJB5B/fZLdO3D2in7/XAs8kNSB1Nz
KRrMgUlsBeExpwQWl5c3Cp/f9s4FDabbYVMTbDhGF7hnz6uyfA31dnm05NVrztSm1OIYMAlJ8gL5
/uU+xUuyhuLX1SSm110E5KKRlOXnDxj+AGEAcpDuutW9Zw8bYEhXO5Fr8j7jzR/WAKxKm8C8Qy1P
xAsMtFUebuuxVwIk8E84H2KB8Sp8BuEE9mD9d13yOHlco4r0dreH9HGCn1RJ7+BkHiaRyP7PaOb/
KdvGOyhyMN6OXjewWduXWGInLcpjahRpOEL1ItwM0DClm8XHUiy8S0ELD/eVYSmSmPednIPSbgck
/+kn65dn/XeQmvun5DmOVrzywn58f+TXWLiZoIu261B9DgYaoKNlFLzAsG5cECoZ8YgItxuxZQVJ
6pROX69Nad981dIc/SKbTgDnPDu4v1O6QhbM43UUQ5gEE4WE6A3R5hT2iQUgb8uX1Z1HVAoLEPFw
K3uNYVBhnQermiQ+oB95GWf+tBVzSWSeNIP64w4YLKAvcbG8LuaVtorq4wx2MehBedYesmAIok0+
B0YiTFODmuqkQkEwh3DYmRSU5LnpHDgU2+gzqtohOa6HfnJttBsATQj544sPkS7TLqU+UFvXh2n/
8Pbb/uBUZhNNkZsFH20Bf2/3d0ZAn7oLJMdXfYlH8UMGkxRic57nkYXuW/TGyjamTJKFtezkv92Z
if7Lx1rZ8pQyDVxdXGtEGl9fFKu6bF3LKB9n/wBLlfjqPytglfeFADIcohZkPyJcKqCpf/oAQgXT
590bV61EVkF3OOYcpoj3ictNAhS0TWneNv7AfsMZGaybHo//ThFI+en4ccPBWNlwtxEPa+WKBGsL
kZnE3pKJW9WalnXrcWwtw6QFLUc8ntRUIlE2W6VKXVgau0EIinOem5QTn1hnWfajhMEHWD3qUXpk
iHgqG1mlu+1bIj1+uQaeS4OCdYp507iRxNK1Rz1QsjfF4s8zfnEx2BZMRNuxAv8JuL2sNuzDWFNx
N+K0VVyFii8gQuDQ6V8iRJorxj/g8jxS1MeoN/8yUsghViu69xvKyOHW3RAdwR6Wk9MFMYlRunAz
0Wf6uxg24pef61gq4CN9OMj9bdcAnh2STCyY7iSNNVeuB5Vodetgo7XbyB7Ko8Ixk0aqZpFn5WYR
f/0WtMTxSwKp6hi3Fz9ra2MMp0wY1wC5KqjK9zAIn8bfiVCdBL3cVPHOwmFdqgHhxeFmuWNrTudJ
JUEyAxC7i/tQVtS5zfjdIbzhSTrDOyIJeGw15/8T0GNOPRm8c/6wbQ6xb3SeuaMhAcj7R5W79uJ/
j/aJpF7fy1t0hV31/rf43JKwer/wMJ/+vgzcWlb3WU9kpcSxgxrecWTz1UWeDF6QvWQhVvHMQmtJ
6ptel/12RV9fTlmZ1JMbWdBRWXUYHsG4oUq4ZO4Td550Z0OB2FPx33NKsY3RZqQf5uTUoHeQL3eN
R7+m3qCudK3d3fBwiL9V+7DponUK8/eH6rz/VIGEY4lAIi0Q9+WI27AoDm+ZtNBmzX2tLtfUUVUb
5+DrgzEItlPqAb6E9c1wMaM/ph64BmZjDxUj/zWON/yjCYZXc4GshLdW6yETbZPyzhiUp0YPaEoc
yeGA5GIUqBJB84VBb+SFL4khZAwIY3Rd3tlc29bTI/tb91uo7YGhstig0M64IkowGh2loMXnXA28
ayTsBFEsgLpC/VEyiN6G6z7U3Ocy3ZLipSEfL46psFGufnl6+UIgoV7SgGYI2Hh1GtMYEb+ungWF
x6XZ7c4Bsx9HlfRSF0i9l/3qbo0+SpJnM3cD0O3ptONPxFNuA7/uRda28KZliuMk6pWm6ZTI+Zdg
iIbvt04BUcbvmcgzkNRcnbRx4aq8ijg6E6pL6xAci3I9QqvoMlcCxdNiKeyonjETSgOs6eYSn3mQ
XzXBzuvPJBkAvaeg6Q7blSZIdBG1Oo48ZU8SZ8bsCvNbhiIM4uaTp8lmo74OS6G2gk+LcwH/NNhW
VT5Uz5HRe7wu9L9CnKcxpHPAYC4kJTABCMc+ShZGl8uJG/4n2q9OhVDiaYjz9IdZxyKlOTHSufYA
lWc9bXwuhMpuFwB280k4oIr02lxPWeUe/ZLp30lIFTsSVfYBdDthF9Bpt8kCCXm4cHD/02WL0GAD
JvUX5Kl18VvY0YY+68hvXlJc7F8wlK8dlLjS8ZP1HMyFaZLMus6l2660Iv+3LBOEhB9PNPqeKpfx
babcIiOJoXftuCjkgXLi8Bp/qJlam4fOe5LrUs4rp+zi4DqiVxH5uFl6Fc6V+bMy1NaH3GQrwU+1
EGM/m/xDtbYYkyCM7thppPaOAGzwFt+zoX/sSuU0qi7MZHGwArZK0dUQhahn0+8+fL4VDDp0Fl2/
OYNuHeBA1nD25y0o28vXlFnNvykbHu98CzqQ0J1Y7frs9i5m5aMeXHwqk5VX1YZ2BwitQsoMENNt
2QKDVmQkqaGn9WTz1Re0QaTAmYyt36XqlF3T7W2+jZM52zRVmTLbbnsff8xoO/XBcQeZHRuHsGqB
lrde5zt0HaRoikifF9XKyW3hQP97KVVVXV8CoBQDeplq7YDTHRuIRtsznkvzp+rzBw3oWZFLOTG/
KEzI0a20N2qz/8kvFOsn91smv6Cg1sjtg6HtnA3clawBxTiwtDPOPPxXrm4D1nAJRMltnIRZwEZ2
qhPKVNZA52Z9Ho2yHwUh+uM2XuDCT3VRhsdSNxVpXzsDGp1zSQQ6jybZoAU5a9rH0umfAT77Ej1C
1enOlB2KoAK5ecrKl4gHvoJ4CDtV9LW0LKgLY/2TJDNkWRSWW9Ath0IcyjkBAtQXaN8VcoOBYC3V
hKHDSC4YRAI/4QhNxCi6QRoaCInjUKx1I0Vee7LyFtxJgCdYZUr4Hqo8tJg2BY73W6BfjwM65ftO
8Fp1fNG+B/xHA1wOTxqlz44QX0QxXOo0LbhxWQe5asaI5GhKx5fkk7MKwdF8gjcW7pcR4LUhwbY+
BknbWrPaCt+cRPQROVbgSVT2+5qzrJNmXJPfsIFhUB7/RmKyKs9Ci7XmyREeVhU4u9VuMP3VWXBz
RgurKFzKCQZ8AGUdjX5kfIH/FcbypYRS/hchndM/LeHO7u/0IceRR4kszPWskoxNb1+DeihLaTht
ZQa30BZo4Vw6QNg+nYXhbJf8nkDuIvlLrHDYuK3lvQneb74p+XeUwky+Hj+g50tIpraXdXB/PkwL
FhwysZmKsInsCvPclOAeFobxeibgRmR6Du33UU10wncmlTaYZCpvNs1X5Iyw5cYS+1vM1FWXo2ax
UelyZl+r90ZQvb8jQlHPijB34lMAt5J6VVO/w+B3zy0RqhSm2QuNTr4x3a+Lj1RtrIFWFjleEyWV
otId5OkvCLBU5GX8pEBLPqNiEm0qjyTOj94FC178Tn90XjoplVxm1SkjBC+asiYa9S0n/JZhA00F
FJkQRgLpgbAcS20ZCDB9FhUFOOZC27Coo6JdmNDBSLy6jo7d7SrpNqeEerE2SpsSMXbatqAfnqcR
YBgoI/hBCVeTyfHX9xiruBVlF80tgCdBX1WvAccXRDiUUNDXqEbapQBY0fvTHbf/fY9P9HMoCStj
VfhjPS4vC+LCRS/5pmdbWAJ6W9WzKZr9Ml3zF9WISuP92W39O8iBUTgq7BgtnwD5nnEoj/pylxb4
e82FFOcX58g94hjP0/MWNooPbSUYYv3CBKdrbUC2etinntmdFGiVVxVgaH5b85KfvjsuRync0BGc
zLGy4x/sQzJB7Obl7aZbJ1c4WMJyKX7T+OWhXKIU9sRBMo5ZRj3U2IciNPlqF15LJMgNxfAQyOrO
97YvFtyG7SWhULaHF88KQYGlLhPI0KZ4g/8VowP9rE4KFojY6/57qWPl54MrKjkHYG1UNs7Su0vg
2swh8vPpbhnj7RrnPIdIevg9+SFclFcq8CE7Tj4dpgh5RQnp0rPbLSV/YAEKzV4qj8KxOdZu8fw7
SPD+k+igEPaU41UswHntNGZh58E2f7Lz/qO9UAf5CtPTWJlmlrR4ob3dm4g9r7jgm2BEVr6gq1i9
fOgqRImE7l5Y9J5fSOIKNyupEJ0VfYDghHnk/H+lqq/XwVVrefR9UvbTd/NOY/Eu1pJMJL4hEtVH
bllHQssId1QsTz4fDESncfxuSwJ8qj4vI8Cl7XxDEn5xYTsbDIBNSuyFukutF5WlxPtrKgMu0OyG
50TB3xw1wIxYcyqBTMQ7bMS761d7SvHOF1GSK/QwFYbRr9KcNEA8lVBUScT5hvyAFyB7M3uW4d5M
6Q30Guz2jjW7riH6jbeda379yJDPQtoneTp986tI4bXVXVyvRJFDJRLckT+g6UUXIePho0xLo29v
L5dzunR3YQ8rTWBw3MLGzDmDRKWhs1r7jfCQnz/SgtYy8lrN3xBD+lSifEci55fbrGWtFVJROkF4
ShY504wXeNGCsXlYbzLYnH/N9h5cjeeaw9bgZ0PdgERy/eXM7gEtn9ssvs0GprdqLLTh1G1mnEnQ
XabsE9tEx2sgy7mgl7S8yrDFMy6P5IQ2v8CSXH0y/1vLNq4PZKJmIE3Qr0DgfHYhoiQLA4RbJMzV
fGNNSvJ3XJUphYZwUSr0iVJeQvgWjF+5Z64lzlddUVOQz2H9tiuvFfdbghngRLCmq0S2K190qvIF
ZFIGHLPqjA7YgWI8/F3CglcxJJQcHp+t1KkXMYDHmjdGYZr34UAqyCW+1TdW7Z0AJxYhIvWIsTAb
/HkhDnHaUQu3lx4xrBmP3lUNtdX3Pr/HBKStWu8fKpt7Vp7KKlkftggN4ABn/CCoYjlwcz3yDeNN
hJQMpLICGfc7x+yvwmlUEMzorLP9Kicd2rrfns8wfr9VQAGnsz7eLK5gUjB9Thzolch2oARSAreL
eheg/3pYv/iwEu+Bh6Rem0jyCEkbbPuL300E+yeQ1blblCCBNgAcWKWWoraJzS2zh2BQ6XDohN4T
JILRbnyrNv0vGZ/Z44h917i0YdwJI9z+sRoL3kcBQ2LIM1tzVeV+qnLaCnpvFd3UfwfKWG3PJrtc
Oscfft3H7grtxnFF3uDI+wN/Z5Jd2Vrz2mBsLFuxgYhdlouKMBB6ppjzezlk2JrKqRT3sCOZhYrc
K0geo8qCZmO8PbTYVRZHa/XuN2Z0A5oiD/+t7opzCR2wKb0PXYFZ1URAfLPBJ29ICK/BikI27PlT
tVuSpCDIlFMS9opWu6Q75LtkoT8gb8NeejlomNczoyGu9jjdhAtZQixmVA95QBlp0arozoMQxXS3
c3LrMJt/ZzxnKndmbKuT3LLJ2x3NisTegmQ2tzNYWVpLxK0CruhMLKAl3P/V96Y8ZZ1aSEIkYaSK
l1OgWGRUi3DWCWDT8wDegxXxOgw1DzxHUvgLIiVGvaZb9lQQ+oMX121DxlWjBvM/vunPrUS3ik3p
S8S+WvZUAHWwW9k7CzpKjCqdQht/OMC1fmz/OxtDBSgmho4IYwztcbq+eZyDtfnfjLmI+vtqmWHp
1xIOru+6t2ux0/MmEBfxxsriZxX3+eCMazUDO30Xw3HxDZj2U182nesLOej2gUfXRpKUQw7Jl09f
MbikNX7oYxNBlqkjSbcYnqP3TMZbbOcoWu6KaiTA4vOTttWVLlc/J4vV9LBDBQeRhIzSMj86tnyb
G7FGEyiM1v++FXK6d0UZlZOAC8GblirXvsp7kg+sLov4WHHOeMKHmrY7CzZl3U8Gr9YwlcqiIO8S
4GZKbReqF8oIGOmehARI+9qh8Rd4l3C+G4DPXFWogM3iLrBm0gVhL96b2MgDBvt3n/VwbpWew89c
3UhHBlLft/ULHrbPG++FG4GxeFRIPQnvy7lRrUxYn0dUEh/6dkbhcerBFy2w2TSLxWSVQdoi/04L
IzzVlLYrPSrWG3ZzQ/+EJlLNCHtUBvScuq02YMDo6WTYpQdghgwVVXqXhTGXtOwUR9U5cgLmKeEW
UkrgsAD9rU+vP4+lMcK1HerZGTPwRSWUC6nG26mo+e3BrqmCvGL2o4+oK597nv3Rzd3zXo9fhAWB
qFyLcuiHZQS+F5at/GmJalpDyXgYIBtMHFhRGkyrT0Hfm5XMPtKbrblO/MRrZqOeb6x5SwNnmu5z
qm8FoVsZYmAp5c792W0sP3T4Dohg0DunvaH57mGS1JWnUbEAmjiL6/VT9rU/bd/+Ky1BIOWDqQuu
ATVAAZNN/xg3gcpmwJ35faVAB77MfrR6HneJiNaXmryUnDt9Xjgxw+ihO3UvYyj/SNoHMK1qKtFr
qPhLEjSUI3zvbanIx5v+ovNNYFWzzHuNRD7ib4nHgpI5JGiLWiQxfKzrBXc/jq+kd23aOXpStbpw
3V9HmktWIz+U8WpEnr0Ws+URPd2MHdwrvBwUgj8RXknjPymtOAocnhCi1bSlbfG1wxm9EDhX6y+A
Wzajh/4pOR1/JQDYd9aURekVw1Y2b+xxnWKXQGn/CqCtBgy1gI55aB5EkOk+mOwEkI5N/vYedewS
6fYuVtN4l0hId7stcFvCqzTmMeqdTcMopbyUPquEE0ADvG3CZUK/mzV18XhDTYc9vd9CGNqRdQ6Q
5vSUZ7bpruR5XEhwVnBXeKl0dDjd8OzxTObU3Hq+BuiEuUp0yq0R7b2Wb6Y1ELx5jBfmNLMCw45k
qtvKn7bJx3YQElsNtAA0DQIaJJcHGz11XR7Ym1oCibkRSGxpGDeaF1r2bdBe4MFuduKEvw9ywUnL
7X0+Ek68Y+mPMg/R/XpbqfqosEsgtqEWH2LZVTr/IQH3/0GaqCNgI1aiOxPBKP3RrKJHGTcFohjG
KTQift3lsM8Xn0CkbwM0pog5uQQSr9ZGSHZu1n865Jmj0F7XsB/7KMCKoZIvGvLGHGLqJDfnTFsZ
+covUx4hC3GfJrV4pb9B2L7l0CbtLg5EuTLaJgOYGOFb5jCFilE7GVR8BFMTeYDJ8PbOLPwwqRTT
ZhfaMTAqu9YU7OMI5u0wPwxA4+fbDjMEZknymahafo3NbsvbLWVkXO9WAKsHbsoRzeS6qgQA/mgz
rBzlT/LNgAoU5effyVE1H8mmdFAX3n+eQAjdHCYRDtVsAsFbTWVD1HDaCT1vk1iIqxCwBO5Zatsw
PIG3uDfhIWt5GJSACgD/+DdguRBLf+mkK9wwGn0kALyWdp2r4oUzuzexh0QAeOkn1OxKivH3ot2f
0NlcBcTnENAWjRcdXerLmHBh5+9ow2Ilqu8+JrGIzxS4chCrcZVVICOawK+K/sRkgx2+1MxZKtU+
OGopO9vfLsn7taooplGgJWTenG0+9jgrrwpHIMWYCw7ayuHJwInBFpQUvewtAG5C5/thAMNAa1iV
1pvri3ifn9ZnsIOuGhYekosoQalcURDN2BBNYfp7jMR5nUqIqUO5MWcED4Z26Oz5qp8UMS7qXU04
oGdh4QqK56aM0F4rQ1YrFAGb+URwv2ZX8LcbcC2xmgXAuhQ1WjPlQvPIfBZGo2OKVetLLO8wWf/g
VXfAh/NGRAK4HfkNiIUnTYgDCzdxuo4lXMwvxIjFc/IaPzVjtlg/jiby/vkfm0bGEEtD2U+qDCA+
6NaDpDCrx0JPPA1yJlgCmRz8UC8Xy+vNHzVUoGthpcGP+I/QzHJdZ36ha6RdKiUdyNUDHP74q2vD
AMvRnWqB9DVk0NJ1vwceb+h974gstL6swq91llkB2dr1qEpjV+d6SYYPQ+sGpD27MBZoY/LJOKdl
WCZH1TW+MHf4bAWWR28cYYuS0PArsVfU00QcU0pUfjaC9VLeNjFZBI2zlElpTlx6mA6gHP8W5iqJ
uB8N27Z+QqCApreBda85huwIhAR042YUqJEmN2ye7bxz09IXwjzGgk9TRAp9CCtPw3ka08IRnUD3
J8C70DGFoE8EzaUGsv4sqLsYViR/picN5GmFuRcuJ6GAHgmNjj9P3sm74+pwqWj3piVeNOUKchPC
xcOj2NPkyu1QIs+US27GyP+VxTaYy517wLFh9r3DO/1XFAoPMg+jmM0pVnCokGIryyE6JcDCFG7H
L8gbgQmKsNIRStz+6VuoFDB0gSVCfbrIo8PH8BpcI/XzUy/GrfzeivWc5ZNNu25mOrDneWOBvU7c
FGpm+/kIeNJh2N7f8ARr50seNyhU/Rg0l1y0ELwTzKKdBayI8o4PWNMQ8G20G43gp+ZRt6ZamR+G
ucmBpYEqlmiPBBQ24VTJpzGpvJfKsVzUB+fNlpi1jRJefJClLrP610wC6OmYa7Txuzgs7C4hV75L
tHU5PGNqfxo/vBZHPMrjQmXcdyFd4hjI1dgRG7vCaSPKAkxAK9VQ9PF+rFh+VLOs4AxhkZnrSM21
9y0Rral5MOGp/n/Fa5h/oiZkxG60dnIvNNJj1qNX9OrybALX5v368qVjZSXKUCiHX5+YXkLFXKul
Ef7+8glXHpnCw3Za5l1SLuPwocoSfw+YbzY6L6TEF83UWKsIf07/dUl+++jtFCoO6gj/xtAmSDwc
hDNOIThxbg/n+7iy4pG+3xGZrNB8Onbmr8oZIyVy9CqZamNpXR6Q+CqF4S5RzJwyamRGCNYB8ZN6
2iKlcUEKRWfYBz+F+WJItrePmcTdgqWdiB9CeUAgDb1h+JDiNAfFYUww0Y23ddubawT3weGT6C6o
mYzNuV0i9GKFfDz/KpJVjftNSmkM/2FD9CTOHHwaHkv+Qw4VE4ypmIE6Vy2V2kEbLZJIoFp5zWnk
yNajLuuKe2Yovb0SFo6CzKIX9Vb7st1k/Xfsdpuu5twUI/79EUu8sETmejw+I1zCP+U988s4Qesj
LqyqqPVOrOkNxqwRIedI+GO34T/YKDQ7HjWmFcemxSgd/eqD5N4pQLMLTHeMlxcGHn53Sr5a9eNv
Zbnd+LWosQhoSxAwAiBBZ19U4GjIQ5fVbBEl5bJXPhHWY8eo1dBKSZnQ3YGofSs7Opr/dDdWx2vz
11Osusw1h6jqxZzILcuglCMlfHbBLOyUxYlaQL4rIj4ETQQhgtBNlYegoHw14cgb6iVYfTuyRxXB
3THohBOO588W+0PupzsoAayRYOaUkdmTK/3YLPRiSl8iHr8iaGXFfRoNVCvNy0TTCpA56+8YMsc3
0PlYdSdVB6rE7/6Fb0/miBmlV314wTfYjGhQgnXGlpauI+ZifpY0vkmQ7OdXlwbprR5zda9boKMf
+GNziy/elxsn4E0Jbnl554DiRBAv87r51ePgyZ4Ff0M2fLF+BL3TEZcXfX+H1G3k/ElXT7UI3NJn
+v4WbIU6NtjvLr4mTRaWu5Y+yE7lg/qYcWhLQPPzZPFdwKuivIzoHG+u7tEHk4DFDl/j3Egv/O1J
EnrOPo87OkgYlPP1dFpjLD9eSet50SOwq7HviaP9fLXoVGn0AdoXb5I9zukX55zuXCc2FSs4QY3k
gG9MbxKNehPkd8pr4cDwUn3jB4/ffy1nqFqZNKcpxtMua9rUP5zVL55roVGvEIgi23JsdlBrxkiO
fWeVE4hJ4C2TgKaPiHsCan29IIBT7vIDaxO8KyUzl0+U7ORcIFzzSSt+Pe/rsM9WvYzVhpYyi6jq
+GLwCSr2ORtWm13mPCn/+gNMsN8uPeKvWv8atHxtCdoLcHVdDcLk3brcpzEfqZEKYDLkBdmQefsB
WpbmXhiwCxG4RYWNlBKdej89dFpGJyk4weS4m/pMHI8fXtHlHTvySXhS7AgjmyLDx9XCWDY+ZYzq
FfWEHpmIGOWpMgAqzyJTxL1bcFiD8scp/SMR9HPA5jkdumzWRBe4Zcd7hf6rXGCR69/uNOJah5ww
Gw/z8EDBLn/ODqVdfexlc/5NAWbIxkN1RPRleZ7g57i2HGGrloMpk3Zh3fgfLusy6qkmMPh7g/Vx
bzLECSns16yRD4Aa46yrQwk3uhfy0ulFbr5lvEpAUtVpJUGPOoEdtUdmhRxz+DjA6zY643EAE0a5
zic3o2iRnuJhjdiPKg7hOwVgwkjQe99nkoKmYX1yNttRVyX0ldJwz+yD64klaqUpyzoubiFdbtF5
wr+uj5AQ5YpcNpw6hnRh8qV5RVaFcvlzkC4m1vitWDiIxXptyuS9UTIzdy4HGzol3BxEz81FRsAy
yf81U9B+O8t92IgeuDpy3tmkdV1hUIluvfR3FcmPDCmtHR02EOlhHXiEnxRLR68M6HQxy967Qpnc
Y8p7WjyyXQQKmqEAIa8tD5i3H1DjHO0FJRI5ucoWdhTp6F6ktx3MDFldrD79160BC6XX9xbqFNOy
EXmdNLpOzkhxNFrvVWAn06jfnOJGFuSAd1fwQEylNT1Sn4eYxqvP0xUKKNcjQkp+9pIvePmuFled
yLKuoa+q93B5zVjQtRYeYIf2tSrTKXA1vQ+m3a2YfiCRAl93RHEYMxgJH8zxu6rEDLUaCzjS7CWO
CBM5zo6zbeqXgUuYwk77ML7F7VPlFUeDiftkl7p80fIcwpkiGWZhhDvTdgD1Joj8Bu45ZMsG5zIt
4752f6K1lCdNCfvyA2GOoQ0ONq4ER23BvY62wNhxsJ1toihRi5+/yJFr15+D95YE7nEJtEMg6CZF
LpjMOMq+7OxAePQzrKmUXJ5UNoo4gLQT5rY7ZXv4X8j/5RgjCBF2F0AMFt1AT/I/Yqv9D7yhEXww
zwrwb9AfNaNPVVzf7EtPhoEsgVPYg0oQIbMEELijv8ckWkLqXDVYeRbkkdBIJJCqIcGjMlUIAl9b
aQVxCX8f6t86L5ty9/5SZ98VmHB7WrbyHJujwijtbaW7mz5c97tjYRuR1zy6oDw60Renhu6LytF6
xIF/cjKZS+pxrd3wWx22Om4U3rR5qglulAN608hFPuzRrFyl6eUTIg+72OEyGFnImhREttjE/pg+
3v1332si7AJrambDgUqxaiDojEyxhCh8b+BPozKszLfTyNF/ZMYSPe4MwbYGWTcDcr6e1lRqZTmW
2vavw3sAdmBGrJ7YG+H5YMfM1OsQ/ujMKDMLJOK2t0vZOffK4MQnqmmUqzElNvoJTH/mSWxBgzbJ
YCsTea+ZE9kcg83XOwbX2A/IW2Lv2mRA+PnhvX6PNTg+XSBITCFv5fH3Ag4Ek9Pu3gNJLaiTRSYB
TVuxlceWHzvj0uiajG674v0C4/wHPoQYJpAQ5oitM9hMYSTHAKwgXa1lJrayQMhPR8iofphMiwqP
Ht4CTTmYRCSS23h8O5J8X483V2y4Fpa32pDSpkhpyz8fp90InHfdy9y3ArvLw3oTr/duj8m3LzMg
cmVzVXdmldxjGgFqp/qitoU+lPLbno58F+tc1pvJb1z8Oj75YXlKAMhfgk/Wq128c9kmdYlbfGW2
bXLLYDPJS9Z/TvRw5DVgAIH+urZBMyg0CNeqMYzTZsDWDt+NsHpWgsm2ATkJsFXfa6lSMzH5RUs2
NJqe0mWE8xqIymt1GoPj5x5bsNv3siywwc8FA3R0hYyaS7wW/jUzXcz/D/M4Ylr6VPqM4ggzIyTv
rfm9ufc37Tu7yPiVrxX4y3HTkgcipxqFc4LjgByNzJHIUm1clRvFHmvsBORc3hkIt6IOoG9wW849
PdrHFsT4hRkEd/3R5+qXLztUY6v6TX1kWgFKe4hkG49AvAjqkiV3k52vwpByrhJF5plEOZKDIIGx
308IvUjYvpZcjtP3qKZ+cx2tPvidPG09pd5FLnuCagk8S/P5RFxMQVa/xOffdkT+VWFJMZtpRoyZ
MOAMhj3wx+7uRKrNwlZilLz1rA/qcI+6eaKfxiD+YVOTxfpPwFATOyKMWF4n2jASkrQkuVd8kRWe
r9pxWLDWwRVzd1JtzJckO/ETPkMOnKWGFyVvoSf3P7QJc0HJHisvMkZY1TcOfQdnjmCppxY0cU/R
RgqcAtD2eqRnnNRcp3K8dzwsldpYuvmDhk0DNJaxknXAf+R3x2ZFdwBtKFeZqH6E02NF9UrH1FIQ
wbjcXO5ZnXkCL2lSxu5Ja/N8xCE3iKilRDKw/mg0Wqgyv7o6M+5ERDIXxIoAaBDcNe+f7zTLIjjj
dXp8NcGAwCGBV00cAYYkmjNs3IqOekFs0qjVBYlApxldoqh5KyISaICyWXndu7mktX13P38gN3sM
AXSoOmWc1m6tSnnRQ1pxJsyx1vgrB42r0igpP3mchrOBkiV14Nz1t0J7MATpn4RWHclLwQdw+nop
hkrw6jM0IBb95HE0f3aOBNvArlOhT1zFUhYwtcXa6KUiKroF1mb6W64RpmClEW95eVL13r0n1Yuc
Avq5tKObJ75h+fvNcxV3edI3Vc0lUyVsf1r3KanqhkZJgWQwEuW6zYd9Mo5uNoT/w2mGfVvWT6O4
4WVzI1Sd8mcWhYsHcHW2gQwjLBZpJmiK9u1llGdf0yUwFDr8J3Sgc+m9df+E26iAi9FiR6iEW2Bz
a4SPQj1u01TfTO0nUap2Ry0b0RGAAT7ex4JaddAw1GlfbCB18OzuF+QyuMkgm1SJFOY9ymY7q0+g
I3YpcsCwDDUSG5QEvtJM8UYRgQNuu1dLFh+agchyVhrq4/nAUxZci8A+CCeJ5/WIWSOjnYbtuBMJ
WM4z87eHc/Qji/qYNZFeuef9oCsDJ+WoQO4uXnOzmXkFbUJd6OV7h7W1y43xARFzzlZW+rs05bfX
eNg6wN5lLdsgaIv/ixrqQYpgWEy/g8OK9PwNLZQRu61sLpINoD95nrDDloc4GNQ+uA72oANFJ5Eg
bewEEIrL0WrOFlMbXbLeHC5fM3G7QIu7i1uMfjcL8Tb+prZUTF/rSd3SdKtvPYKMR7DR8Jdu60pV
Oi/EcuMZusoC/RMa4dvRXz+Tb83h01zRuo2X6+LfEAOeoxiF8lAVBPz93bX7UMwJyiju+DhKnOuZ
eW1wjZ39P1J26l1IfM7xzSPnpDkZKAtB520hF+Mj0VEUnciR/A64Mi4EB6if0tDRlG/iJwksw++u
OqvSKQC9Bv5aDhNqLhew6Q42ZV+VR9LYjhlCgjLFwPzTUZI3vfOlb3W1oPrFKp5YUZTFVHF+o9p+
ocHt6DrQCFyd+F1rYyVQrIzNuUEQ4Tms2LrScc+7sdZPpoXK+GfKet2g6Of/MemgFrUGi9eukGSR
FjT+gbtAstZJByYFgAnock4mwJyn0opvlvzRK9ah3jbdSLvGL2HBFWhmyB+gdhZUNlhzD+9qmgNt
+bWtBMzhIYRQhFMDp1CYlh04aZaYn91eBWLFv3kyhGEgC/5hK7LcnqkkYxWfEmgzoyS+M4Tb7Osn
qlbsFXovpsQwx0qkoSKEYeA2sgL75YiNabpxcvbFLGIz2xqzlYvta3MkABSFc2It3tTBLbzAZMMM
iw3/9SfngT+JcbseULGEjxooZXxe0glzrW02CFpW0eCmhoPNMhSfajpR1fxLI3KAUlRWMlB71vEN
BWJUDa1JnxavpYOKbdH1+HEC/2KY6CPJHJ2vgfTmDmxNSigseWfPLXvGQwkx8SwjBc6zxLiDhnmA
9B8Tz1bSuancCzpogZPVK4rBijtVLLUf/XYvVODF+r1jRi1Di2XGI4ZOq8uwhaloTa2l4Y3LSuNs
DCEmpo89eJSUxV4q1aUDWtIKJMURiJzktUHS+x8OrPdbOgGqikdycvx8YTSEHdinnQaq1LtR9ROV
Z9sHwhR8AbbkBGBwmXTRFr/fmSYkqgTwTNX/E5MJPIVOhomTSi+vR3TbMy8Ny/dpi1iVq0BOZBLo
B8a+6F7XehY1EIkZPaaQatnGE+0aK8IvDQDrVA8e0yT1Wi2Mhaiv2oUPl6j5W90q/bG371y37x/e
Yf7YUxhxBb01ONisueF+FoOWS831J9yeGWhGgqmxqH21/kYKfKp81u2H5HpeTkgyRXhBQ6GPK/pt
EP3ZZdyXrFZtO2pebwg51twjifQfQ9rIPhZMujx5mQWqVW3xggSgoQFj6dmMS/cbN9KeSTG3iqRh
RfAlaLFKlDnkxjJHBuMRhBK+D6nEv+6S7PS9NEqDew6JbSM63gudy/Epeo/1ow2SSSh/zWdS5Elv
95rqUFSAzb66vwMStGheWwvFsschBqvbEtui/h4sG04d+Fqgd2s9/Ar0aXwRjRZYevh/zuuFzRGq
729PhkRjsXhq38/uF/gEORdBL58sxxKlbd178AzOm6UDa2HcUgdXmQuVTyUSs3lsDwapHhL15ygP
RTIgdLwBW9aGjOPMRUasVtBs8/cJSJwR1NsB0R4L3Gk7odbJ9FTBs88HnAg9wab1cE4M5SIJXMnl
GPVkHnHPuGX9kvVwDTL0QtuaC5NMsiZ8E/oZ3rGxZxCBEbxnlXO505K4RGuXEA0bZbtLfEI57PNd
6Q7PquS8Ii3yQJtzQ9wJSG/A6cARwhBQEXFCnZS3/sx8q1W3xyGzZE4pdOZHLAnXOrryydPUICA1
w1e17GmMIUbB6Cl1wIydCGodAagMgNFRcBUtkZ9fljj+1BcW3YHxldQLiXuXgcjMv3pwnQpI6W8e
AK0h7Wnk3S30arIvTXmVk00jXrxGpsoT7GqgbJbm7VDYnt7QS/kt8ujCUBogkkW4x4AnXVeAUSc1
AFZJLL65fl57ANmbGm1JW02v9wmLdxfqyoZzBVbNFXlCs1zGudqS2uqPNjcxUCibUjqLOdjYAbFY
+MD/vaLHUBUOmbwSW0Jly5AUyluGQVmN2kXPat9cfgQWFw9mw8dGPgjscc0hKVchEUF1z6O+q4Zl
CwIaQgKKHf779xfOeLmJCVoM9ABuxIh/sgRGxqj/6vAdeHyWCSskmGv1ffDN4I8hr24/Nssh2Y9z
TI6FbKIk6JSIy88nq3xRWnw46TcUWZcBUnXgYS+Ypfa23oZ72wead5OtlK+FFz7IR551BpSh5W+D
Bs6ZjgXE/V3lb0heD/nY+qxKaKtqmKVoNoeUo565SV8bux1Gv+C7O6QiKEqpXf2t9suINdT6elrB
1kshK3Bhv7n+KPDVkTiclQLg5NzO5k4Un5sA0aG82SsBz+/FSDdiMR66KshyVWIrsTnA2jlHf4n7
wZKyk3FFEakjTc4aut5PgmAROG0NK0kZvOcRPiDlXWd5jmZPhQ2RS3ZBi5ezeJL0/lxyFhY47Brz
gPl9QiL/9Lr7nBnVD/MuDkE7I+E9X0iGOv01E23GRjnnvx/WIWFMUzXvh2tSH0fbWkuQutl8IOai
LwOwm2A+XEvvj7zEiIDmEBZFP19BL9dbXhPpcX96DFY88xNwDZWN9r8D/dOpLhDejRkbQOfn53im
QmWHmw2aG/46rXV3MOlG02rA+JJpC+vGnFpYud3CsI9BgqF/TYENG4HOYY2BD1idTpv3vOBC8A3l
tleorPI554ASZlIQaF6CytlY6pAn81wJ6mEAcybNivWzk6oPdakDnUdERu+naGaCjE68bJzSSOeN
sisL/G2QApl69/tn7g08auMEBhaMtL+JtQzAb1z4CZUC4sn6OFb3L7m3EUqphZo3PQnBZaLlCFUw
2SxQe3HDAMhPuYuIYRBEgNvz6ronFOaNaGDITO9oQ1mU6+79o9Wnnnx9VazOJQPUpyGuIYAVvlp9
knoZKP5QdJOjnb3YctjWbsyxCFb2ydTHEPoh75oDf2fhjp1cBMAO8wI7c75wYjjjONrJY2RBf5hF
vY6cjcZgeUW25E4Qlu6UuSkDhDuh8sN0omi7nW24MEUwo3nqdAVWAiobhMbRtuPhFSiKSUfkxit6
TQV/lBNa4zakP9crjqXiAQ8wiWlH9x6fRzg3eFMxHV6j2KOj4Ml41BVYHBpy1sDtbYnMPA4d6poo
jVvhGtK841KjwOQAoHIDSMzL6InanDTv+V87TT0wWq5PSkUcGcltSrnOiRdc5V9ZPUbFEE42HSDZ
ucbJuOhuhonWOaiTPf5YkgxZETKLMCu9eTcoqKih6adsxoGuiYaVeue411sk2UQWrMtN6XVJEWIN
heCr7iLsCvh7tIOUory8ZUTAPZ8PeB0iy7kOh/Rtxt2Xq148vz4VZV4u9Fjjo6k1N6gLhuU3++Sa
dzVEhaxCcFyVjs1yKc6nSbVoX87avGw30BFKWVZskfNAHOA48B1L2slMvE6WYrtcrlMfpypk1KE0
wtJaRnmhdDg09vWXtbBoBGmMZCd0jhBAIqyxn9OS6SsiOhqTkAxK74Ojofkv3vEAdWdHpfKQp7+i
vdZaikF1QWvQimlA8wJC0HC8JCPsj/4o/9LOBZfvMP0xGy/Q+jsAp9HJNZyP2dZPo8BMr2YlYSia
QwSogAJvx22Bh75qjTNvmZIyXA4QQrLXuVFiZ91BFWx4ela/aZqZeUl9P0Y4vy2LNA2gFh9B7nBE
sdZKvoM87s3GKceKpYPIEikLZRtY7GpakFv4+TSv1nXA99CxpWkt4hjrOrEKFxEPWIRvVNv4bVv8
2bss9dVGqbLbib31djN6JdymhPH6iCx0DC1zWneRBJNWqINK8/12drmfI6rv4FNIK3xc08ehuHzG
NL6Zus/sO1nex2wROScJ2ottYXVmDwatV4vTOi9jsfbrJtLZYPctpuVKyW7yzgoZ17aTtJGuLHli
JvhwuERLj4G8NR1y+MXfqWnukO4o8N+MQshjojPuCTVo1tR3vy52F8kvlMC1rvwVrLBhh1RGP6kk
HGjUTornzjyP0Ui8VkzGRORu5+PXk2xqQh4lVpftXmAsODwl1p35P2vs1uB8Nxqt/Bj9UA3kwovt
N/sA35LnXezuZqIE25r9PAWQ8brlqt8V0jW7khlxwAWkKtD/HmJw+43WZrqU9u0lnJnubXbxfQpr
r0mVCTtT0L1OqIL2/mG2nXDkd/m/WvZSigYqRtXCVwPhVfPbRARgnKNwHmP67yw1Vi/YSsoFx5Wp
pivc3rJddX4tx5uRy6NiFHUsaGLfMmSuT+Rdby+UsFC+R9P1sOeAyp9wh5KwjR2aTXKwRzBsTUeS
cuaX2qNb9OrhfyTUraw34VJlvTz15FInRl/UuFGd99YDlCLFUIevBFybtg9KJ4loEfVEEyrGJKZM
lyq5vWbfha22qSeXCv953/oCJmS5nhQgLTVj+xl+06L/p6Zszs14+bVZHYdqNdxR59WxV+l6WF5y
AiBI7mqs1BRHRY1LZei/6JhAv/fW2VzKCG0MO2lnyNP1DvGO/LSu0wJfDZDuqkWiHGI2jxbKjlOI
3KJvqai9IaMJ08RlthL0lxaV5IsDak+JJCBV1CKqZ32jo37ta0dcmVsbkuksb8zbdFmfaCPLonmH
fnUfzfXi8wedbhvSDnVk5+99txiFmwwUmsE+6wHcRcsiOCJP+vQem44kpjZ7YsrcV4L7o4Hu01Sb
ftYRcguA/Nj8bYWMwWA0wuimznBBk+/+AA7uctXfj7oXi6Gzju4sxeBKmC++reIq7xmL8dFFbeUz
Au5YXU99ES7TensXYA/wgf//O/50OX5WcEeKhZA20xadfffS1KcTU5kZlHao9U5YfnCJzJaQMZ1l
vAm6d8t3Qe5YVVQOA2Ui56oLj5pLZUOEuZv/y296W53SEvcRpwEymZxaZ9e55Bn9fCqhWqE5bfKE
yKp16PyPZOJapRj7AWL9cNxdCugpOw8TckO4R3tilQsWMGSE7nDYpUU4Fx1SiovmFUq6/NOkNorn
scS43TFSKVtC+v1P0BEeERVnBSk+H6U1Pp6jJ+Af+V1Pi6GFuw3FcJ3kP/NY+KFJk8pALqyAGgPQ
0Tn8JnK4sERZ0OTGUdIRYlx5AouaqTlMTtAImGEyMYWB+fh9zw0wf5za5OSReXw+vhbSpSBJUlVr
EjDophp4k0Ri12m5MfKjXBNrNwyaP/8xGdg0oEAVhU9DXUE6yVsOib08nNh1vAAUashNrj9dpQ1E
nzYxWkIvaZeO/IW6m08wCBF178FFEXEkM7mUDFAME2Mx5+avUUD+ZFdaonho5HeV786uzi4Ca2kE
isDz8Gg3pSRCMW7vLDf/9ILCUh9WjAdj4f/ALrJnZB4al0CcJWH9rxZRcao1dH26AK4DOgbqG9dL
/PBxLiBWNp2SqTLV136OWmhWeRQC4Qhh5griVj/5w4a63vhzNpCxIfqRBnC0LyNP5CtTylHmrWlB
2FTAZThLy73+3OPHFr7U4huZ+OrMFrxmWHawas6hyR8whVwTheUxxf+H+IPNqXWkKe+T+k78PGdo
wwq9pL4v92N/gwdH7F3y3XQnfkauDgbO6o0TEinitO5ETuKgSj7VXVFzl7nFk/amKCL0ebFn7mvS
rWZnBveYfcOJocTJTrzMd7AqHAx5Ma8FlmU5nyt3oIyl4UmzApZWWJZfeUkBW9KcuKn8YqqxIzuA
9xIzrAHGK6VFWd4vZc8MTB4Rz4yGoZZ/DaekRIjNqNa+JNL+BxX4FspNfFmB8CDTcgAVbgVsSjCu
qKHqnHpwEV1yBzHIY+XmwCh2pzi+Uob+eYAS8oJ3+5ScjjuEwIaCMi/GvvBvR/d53rKX6r4vaFi9
qSg33srspJdPOJf1YgnGI9O3HfonzNfmkq/fIGpnjo5cLYFfxpFCAjaxOj7GDhRbs18rNhRnUox/
CqPJQS9FdVRQ0sz/Zrg8kdXYMqOwVNcujQPmNZXxUZAfi77WWroshdncPkctlAJwGP9UijYFNbCy
x2ZSKu4WfBP0IvF1yRjWzRXhe70xL3i8hziprvHnxdhm9OZ2sHFt57uxNw3jtT6/iR+cfz+JkS/M
ikA4FECYV6Yg3+5THyRcptZHR3wmFgrE8muX4gYHi6XexaTC5+MlPZX1x1zvMI2YfA9Iu3G6QySy
+MD4fx+pa7BfbaAv4ZOU4avDZdIjO2EfMpIJu3Oaeyhz0PEpUrZsuWzbXB7PxrG4xdb/tNCcUUq/
JxQFntHQ/roYqlKXne6VmNuV7flYmkh9yMG6BcrNYiDuoEyacgQ/dedgEeo5AeRO9nm5TTzy7bzL
SgiKZ9ndeSTT2E6fAoyY7OOx+PLyaiDElZXqJ12HNWYtELkLEz5Yld9UUVbCGB59LBmVmT01KSN+
waE1FCbiPh0Zo47/uWtjCB8Mu6XubHtgEPMluaQMynKZiV4DymtJ1D/+Nw2e7QfCaXF5ZaLx8SyL
r18tETAAZEUWokGMty8zf9cfi9rye0RfhPU7s7rXgYt7DWGTuh2KZcUDYza1bJakuWUuf9MSwww6
mFx6ASspKrhEHdSpnJ8SGLxPTC05dWo46OFFCbhDRi+fFqCbVR/Ke3nt52BqCKRh4UDtLG1/hhwV
Z3uZmWg78hyjDJQPNBYsDoE1Rljs4341VdxAflIMzO87e5Xm1x8EZgtH3lTaszUuNxXZgGnEyE7q
sm7SYmlYlUqF1ozy0gKxico7rcnqBMvJFf67wiIVl21I3F+GaYDJGiYZMfCfHQ2sZQ7Bz5gmt8fU
IRsMkFQXesRxI7bUY8hGIcG2uCkrHx47ws+Dwk4cIFlrWxw9HaS8BI1+cOALrrqluIbY7+mprw+s
pOn3G8dM2zivj5+zIMft2XFjcBISa3rZAg9cGjwH5QeiLAH9UX/dizSww/XJc8vv8OzrsHjdLw+t
hfd0Mhqv+ML88drvpVlxET+2snfa7ItIjvbxY2XmRiRfMc0nMlOTwd1jXtx32//kFWrz54lbMzRB
1VdWx1HCTpEANhlPzDpxvE0TKnlS8ZEcPZ/vOxbBGTrrqEIAkqjZ620+W+9VQWdBug/5rTjokwym
O0xGT+1cHdMcfM28JIzMXTbZzIfUf6S/KYRNVejrMmokH6FDBYiT7ffz17OG5LljJjrWXjJYNydQ
OfXEpuBbswqmqGdiorRUskWSZlV2WSRqkWMvxrNepvM4ar7XfB1WPvyMzuVs6wAZX4u9dSfL+GVY
sDNveEhwQiJwIg0uGo9Jz78seMKIFfvoJM85PGi3O2ZGTa54laOzB169GdpRtP0bIx7UOdEOL4CJ
KfkhXbrl3KBO7zV3rA/z888IqszIsmNDlLU4jdfvDs6lbWwUc6I12pKpPrq0ZWdG38MjW44P1EL8
yjykzkWd/qhF53WX2ZGyDHc0a471XiIKT5qpp7cv/LC7AqdvMXGKPzGnZny1o21T0y9dovKkRbE8
MHErZ3UO+PkR76IOT/2u5SuRZ6zEcomJP5GGty/gdhKdVcjcph8TiwlpaRf1X2NyNt8AkvT1GlgA
nWncKUcLK7O/C/mgT3bmi+tsSvQTb7XJr/ckiyg2ek8tFGPuKiNrRu5+tEuWKJvvi0v3UFVJxeou
gevY5babffaeZcVgoxtfY1ly2TSoO3RO/NArSPK9uvOghxmm4MkyKr3dPrt2ij6EhDZAap72VljM
LykDYokhelWp+D/pcvl+KpEWceN3ddnc7szWBcUqUrO82VivHO4qc7XdXmnB8420R+1JcDLJ5Mnp
4mV3k4faLoAuVp2+J2kbOhuDf4fBkGSe4MkErv5EHiYrNL4kL0/nLrtZlYkkevlu6qbd/Rbc9rI3
V0LYvenmKCC/IhvClZ5HW5pn1c7jtuz0RakHwJ+5nclFxWRX87Wz25XA3Z5HmcrFmQzuRYV971Pw
6lQNIm/BwiBi16X0OkVdx978sIzEvWtFD3GtDY3jSMPcFxdDioP9Q0RuZEOnI3lqMjuVk0AK7Kes
Cw/8kYTvSDej3LpdIMc2FZ15pPpLz/hOcTJAZVEPGquK0+TWaMwsVZ6Q/IaCf04aw0lqfkX3BagY
RdHGTPdK5rfL7kt9fOeQG4pwHlDFbXTnUVSB69pSnzg29lZ3x54fboykLGHcHU0Lyh5jwOS9X1lv
iESfMxQvgXOiXw23haQJb6eoNLj3n30c3FGg11Ki4KztYYMsdjloRZGUyookbumANKin9ZtBclu0
Yg6LevQIZ2bxoTqWJkbBtZovtZtjWL4zsy0UCkdwNjUHdBgKbdoMnqJpfw5oDewsPhRI0ltXYmpN
jtflUMTUZhEW5J8rUBxBtbu6tGbTqlxRZ32lhBKEtEnFiGjUIyeZIKfScx4tpqYSfUHsJOW069eP
uORGgsAdTRDdZYa3+9NbwJMaCzhNjonzkQoxm4O6iuYDgzNCXdskr43eHdWl7reffzghHhvnx2D4
12rc9wFr/tylvBP5CBmN/95VmVZ6fkhLwRm3JXqCq39hepng5oLW7NcvMJVBxd9DOjKev8qDwfIp
Rn8Qoh0mpPYG49npBpGbml9HmGA7r7spGM9CB7yRkI8sluyeHNHidJj6O2ijfFPiN6aa8w/u0dW4
cEYLgN/SYwoI0WVEIWhCmi5cEHxiPlKfv1RRdmcmrFCiO2QlsUp5KW/EF6D0nnJyEMLPrs5SMShh
K2RX+j0Ow1qBvW6g1RoKmOVj0LpGmT0DgzlVoMKi9AV4qDy1GmirZpWRd6HeLm9oBryTbIQehBVr
4xDHoCrkWwWE3ay2kpiGhPPHK1SA6WIoarmZ0D+NabfZZvlgTYg2w/ksjU0hcNxPdqW2irTjI+Rp
bvw31RAYK8xFo9qbVonxv7ZfG4SkjmKhWytJ1TB8GbID6n8RXk8ueQEQIDB66R/m3NESq5jJ0jGO
XnYxmsbExZl/2zjxNCxR8g0gszqQ4z4lhciaGyA+EtWEmch5ChskfWj5kmoNrU8tujuWinANqfrR
/7PuMauVkJ0v52MO1q7P+Lrs7iYA0P02+dCrgS0KHGJuwO8s5kU1V9DGQVuMT54NjGMhoSZqUSLC
sI7MJGbNJkyQAJi6PiWmtUTgyvh7VTYhG3TtRnzf/pI+M3i86DTVuCB9CyKMOHrDPtOGUDNBG7uV
H7il7gmyGAWhlgHp1a5uvNMeuW8/pikYDu9nNkDTBzQnyCUah6sqs0t3tox2+laAX6tfXowsXSR9
Whe/z5fDNIjQNKZAq6XSKKCfgRaUZvwv0ZLjqIbZCdRf/Bvc/DYOaP3DHDeLfp2eEF7cDrgSCDCZ
XSu5uffa1bv+mOfTgOFAd/ybxTL3Y2Cv8FcBUup864o3aGqKL81MhglPm+YfGcV3q4QLDk1beiNj
kv0ggMC8cF9fo5DZpsVTtfdyjSXdu9b/t+fEbVVBmZQxWW8b7eFPgKBD5rheX0KxGab736eFw4Ma
FHmyddzk6aeQTBNi2qAU13B8JAkKSIeuRpdM9AmwkeMnHshttq6H6KcgqjFqRWlkuPOftn2wemW2
T6F17dzvy1ity8EqpVp6bGmYsgPhqz/aabuji7LdLE9MtSnxlQYni0FGRfufDAUbs/YoRC40LMMZ
kK0CAjMyOEK4wUy23tT7R5joLwGfEo8rVfaDiNjRdr3rnxCyNU5vYx2VBypobL0SW+iQDKTzfGjP
fGUOMe/I+2t/3+ooNxzQ8BVF5R2zNUDe38p6KMXMjAilQK+za85OvGGm3AlRXBlKLjZW2hlyqN8K
gUwtWL2kC1TwdSnA1GNSO230Mr5ft3NI6vfCPqW1FuOkLTPS0MgG/IUdEvplILabyzR0jkjBYaEI
CU8nCVrlp/hrYxGP8GdKwBlcu/snrlSLWWNJTm9ck77VTAB/SdVJZx5JIQy6V35Xj8A1YEW3nrlN
kq9j0ggodsqh2AjKl2nZ1wmJU0hVTjOOGkI8DkCJRUD3DjvCgVLgq/Xj05kfnWDj3MFWipOBqpur
AvEAjSbRaWRiJW2KdKTrYVXPV1t2O6yCCp/bYFmLC8y49ECfVlvqQsf7d6odKjvFw4vRqUfyiEv4
KEdHbLtndipueZZISPH+AwLsZtH95pRwPPSGNOis32qyLmh7Lb2QJ3MI4Y9SinY/l6MUo++ygN6z
kEP9Go2dsGYiz5EDF5PPnL7iMAMQ0mstDZZu71aTFvTjLPLGdqh7i5XzOdtzWGJATyDx6qCMxaXu
UHdyCRq1asc+vtpBa+q5LM7rPCisY7tDUviSvfxcc5phgZtV86O5llFH/B10gtAn7fcUoMVrs7nX
6RFPawcTudmLEgXJF3O3swBYczICWfOzl8HHX2XQjDcTDhje9Rj7YRp1WuaMQoUZBxgE7QsAtYb7
dU2IxP7q2a13npBDyLD6oOazLupKe9Xvnsx8NqDpx7IqFiFIQ376ChF8uKFeqXIvq6wju3R9YV23
agIluqoYIaJBnnkEeO4KaiTpTCsLSxfBRltmpycwehBdlsfAqynCVel4S9UdoqaaHyfAZcX7FlRH
94nDqc7UK1jdv7n/Mwqeaklz4MJ8gFmMRxRDDt7tJRDqscsnB4kCPIyX2JLo5ZEX9OqNrBLsR0sB
Ati4eQ/J1GHImrdIi7jhw1YFYLHMqtDQo9v9qEzo6cMTv/1LjrWJzXsm9/cFqugch0idlNzGMgrF
sqrnm4+CmXsX5wtwm2MbBqQg5ahtJqqncakRFDCm3KWleUxLlBFEHUT6TBPSMu2+IllvQp/k+f7o
APRyxgCizhNDfeJDnsjsiOIgAPNHYKw6pnm/Yofb0ye20Mb48++sYFkHMem2ZEze7ELEGg8SxW8P
A3pqx30XyT637uSfMdctrHaV2ltcINKp80ltlfJPslrGR227/S22/9BPXwq6uwNz8Mab1TMcSRaZ
NMibHrAxtOZVWQuD00pBzCPwsfLNgeo+O3orQd1mvmhaGFdOuGOsgA8GzjBOAY5HjOQkqw1gteAB
r2Piw2X6VzG6P2jjqCVlbZwDdfNHJW6bxggRG4o4LTAwHXJi+9O64afL3mtfyFcgmzcjt8qWVIWO
bdB7bHlTYDAdA6ZvVupN3T4vydCZ3/8jp6sK3jXHkLgoOu65+4UC1vROD+T+uNDypymRpAYDfUDK
zCS5VZdEBiOtGOHc7CE+d5RvOUBTpWdnIB9wX3XJumTq/i31irisYKLXBfWup33/tHTawB87kVv8
Q37wgljJhDFzimmg1gXM3VX1cUpDjlNhM1jzFTAeEiF7jBd8AV+nEoxVfOAPlHCIKUxCkOqteZTX
o93zj8lG/eheXhRz4jAEEhgQMyIYXwmxAgNuFM347Pdw/X5s4QLvQGoMn9L48jlmae+hlpde7l0t
S8EHnO2n61oq2AdowKUR2fXaNElK8TMhXf3vpcHdYvkIg0jFgS9XeppJwe+RfOUEUoQBT4gO+4pf
z6ueBthsC1X0jrfTAjKMXUtzpRR3XILwtcdPsFdt6F0aEaats5U0yswj6z3wr458OySFyYIXK6BO
QHV0aDCH+H30nqdTSzsnQzkZP7wCpEWNm9aj3NHewtWK0vrMTirSdCa8vZYi7t+pAWLKEcsfTRdE
ag27qfiNLqH2DXUSAa/RonZn4mFgr/K7xcc+hI9cDQeLIYt1HFz/xhERiG1DBpcAGB9qCp01QJh0
87FYXgLEDTqrummk129vHVDSmjIMZ0+jbBXP9loj918coNZ1VKLAtK9waR1IN1I5MR3gil5SA/9L
7/1RRpoOIeFmVP1k8Jkc517AXOHjxgZ6GJ9aeIjZ7smxCJfpK3wCDfz5C9MrCScyGuJ10yGxFqFD
vfK8NUdSx1sRk3wr2IpUUKOwXG5p83ghosFvSDkmGWM2XFATqC0om3qMQ9Rgc0oVWSIMZM+J7ZmG
s1rvqvjOotskww/IEKXWtsBiD5WpXbzh8/B6Er/40eyzpTMugu84MSj+mN5BMa9E3zd+rlTw4Fn8
i18/PiAsvaFKsKcQCe7Z9Esjjx9sKQU9OFBV0VPTtjbkbaEaxjw8sCUCC4R8pl5cokobAveMt9YE
jJbxLTDyUUxGsIRoqi0IlR3ouVqmPLcyuJRsqxBafTXVPJyuBfq6A5K7KJvd7o2qoNnjVwrZQNbX
xYmi2i2Hpt2amq4nucKg5u7syPmypkybe1rdBc2F6uYVhpKjUU3WTG6Oi7eYfV4b2ZTPUBgvCpwu
vWP4aexxdOZ79hTUznwG1A3o5OgNCuwAkV5T2wfKSnhZUB5MzpwrxsjToZAH9m9Hwen74Nhh9iWu
tW66LTwIabQQY6qfR10an/utfJW4e5Hy9HoDMpYXCc/jCMnw/OAK4FEQQV7wLCBnfa0uC32ATshP
ucX6l7j9DB1alpJP+Hwxf9sAat0rbc3s9NoWe8elxuU3IuQVtR5Wb0699HuMeXNN5lHFbh65s1RM
7AecZ6EKUuQ04I4cu/Z6RzA34SUBj/asp6dPX9qpc7ksk0DraOy2yoqb9cP5j7p2FOGPcqq2XsYW
F+GhUiZOykjXsuJ7/h0TSqJtcnbVwgtgdsACVQ3OPtffsJLbJAP79VZIe+kiOYwN3qr8LGI5/kIr
UU8gpgHBOzkLGBRU3Gw1BIW520q1JZtsZtflN6bK+gNTXU/Szv4nBUp0Ay6+WtxE0qN/lvT7XMlN
A2tcGYhI9PgXs3YJdO62y+MVPDBXtTxmM/+h9o3z1L4thp4brdtNCuy/qd6CMv1clMS1NYBZuPKE
kpAlOMwIo2cmLU2NccfhQhAhNUJcSultrPklgmIsxhOJQYsu+TgZTRA+MvpsMC12xpKURMXfS5ys
gzV4drrJNHxGQzvpjSRIQr9+Ebpe+AYd/Z484TqRPWFzojlFNxR8etLKY8xE+gwfWaaEhowtQwLa
3pCnIrV/tDQX4m/XbcWJo7uTdOUjKVj3wJFjbZdR3wyyO5KwaWuflos/4xrHSE5njjSx/34e1bs3
EW2owRNPCwhk0k+6G+/v2adSh2xqZGWb9fCU0Bde4vEXLygLn1JYdPEX3W/3TUjI3wiTpsxB5d+N
gRk/KWCA0msU26stwC4/whfQrql1nZOyGWP3mDjuXZWR18lyGYuSPRH+oAzLMHyOSXLCE/LuSvIa
OC/rVNTU2cKSvcolCkD8jZ8ymPFHKB6kFNDz7Ap1+SSPUBJuuyr6ZxJBoD3RY9+eNl/Q/C/IYwp8
kTcwyoF0GjygqJ7svaCjaQ84KbYO52ps0Exx9yMGkB5nvfJDNN84Qyn/99iWzvK+7qK0VfHA56wX
vW9j7EAZxNoFoin0TYIEjOoFq3Fz8KIhDApQIUySk+qON8okuDQUHPJ+ryVDEwh6rwcHqisS2TdM
9axII7wtPwB8Q+u/qN66Dbu8OuJK4smv8G3tj/y/YZIbTNMOHKGdVIQHAfM6TIiWr8Jhb4ZN283K
7CgYTHfgta64MkNQfGcEA4lvpUczMJeEi6AmEFeLwUrXxsj982EAvse9eDe+z1PLWZvImErIBN8x
hO2/Rg459dDYjn3McyZCSMiVylVOyeLhkELi3vWrlv6LMOb9vXcdhAQRIJzxQl3m29NNkukfelNU
3YbWCpf9DcFndd1I+mfkL5fDLjTPxcaIdDKC2HrV2HklXKe7NblZKIy4uz6krrOAaIxH6mzg9RMb
AGOnwvw+KlBR1C4+bi9XNXrO1CAw+d84UK9VlhjsCjb+AAygB/tBM8EXMSwZoHlpB2qCZKRmuEiU
uMnR5Gna9qxLvsJNtKpFv96Nr6zGTr/UGD+9xaa00mpi0rvagjdNai6i2YJuSrjJBrzSpP1zu94V
bDTPkEB2mEzqPOAJvAbgd0gn1w3ZuQyLGDF9EQlUOT+/22Oi1fRMvruRwSVCMYsAywdCvyWbzaYr
o2s0DWpOXbU1haMdX+UPqVIaiIbU0nkhOFD1u7ALxkJUeCC3EsCghEUzRvYLU8BbIYfmzOIuHxnY
+1THyLlHdCtQVMPHeKVI/bW+JSa/7EynX/9Hu5zpoKRub7cdgMiEv1c1UE1AA2PcHrNA8t0VAhC5
SnnPwuSNgEWb6nk+NOmHkLSsJj27HnlV0U/DtuETu6Dkb4sv854PpgVYRnD3Mtar8xGqmVi1F75h
QCXTmIB/0aEz5r0mftOVvnp4uHRthh5PVYovIvtspGWbygFLSW6JoX3V2uGJMMhWqT8GuCZ41cCT
+OQblC6pKnjVwlNzZxGSxO1cRYf0TSsWYlERobvlANsa6AsMQWHhWrVxPXztcD0rpHc8rOYiMlF4
YcjKcND9LwZh1mChkx7x+rmYI5tvuJ9GD4QRve0oTsGVK+LH+YzaSg4wO0ZE1TO3afpHQlAH24qU
h7m0zbr5osvohVvJ1iovMv0xcNp3vlpyrHJDBF8sZ6pgHsLFbPLAdCuB6mrHBcQaOCsbyEP4RMfI
LunnzefOS43Jx/Y2QRlpFf79d9dyN16e+taWNWihPRHydV9MBFIN4lTxyQyaPLUfkO7eirVATKV9
pcsmJSbkLAvYUBJ430/KTiWu3WIhUH+j+VpXvWl004kTfdLDE7N24pdWkw3k029ku13xGEojGr2G
jf++SsdRVZWduvaelSqun5ku1uf84pAemrpzt2+UIrjhfu6v3IZ3caKsrKNP3sHFe0fU5AxV1Vuu
9kOiVlQO9q4Bt4IBxtfesLBGQqoxfLCym/RCWNxAAZ5tQdg/E0AWBn2vFjrogRXPGhSAmd6VzHTk
xa04zaH0lQA1eNqZdtr7N5WcwlAfFw9jzJFgVk4UvSauq/UaEZn7jcSjDFk6FiMOxhV1F4DHnXzf
rOpE3SzcojncwHaFHaN4rCGLkPKPUrjo6lX/8Ne81lhfn95nFcgCDcxv090LWwz5AS95tCyCqlMy
r4txOg3MFyG2zRCUopCs6TE9G7pBc68xFu8kOArZwyeMZNf4hu1V/RAbLl/41aCNMISks5BjPori
IAXTiHYbO5SnGqhPsWa5vdLjrhf+QJ1f6D5roWvh5x3EjefCZT6azWcw+e/sbW6wMtiVdZURzVjj
vdci7Im8DRCQ3VbMR0Q2d8GfkdRT+s8lH+PFJd7GD7rK7RMl5B6fJj+Ea38Q1mvtqvXJHDY1IAY6
aUWg2SsFfgmfHrUJZEtO3evU1ftf6p4/flDl0SKGLLAFGY/EkPcHfBNGQQngHoMsRkJrQq4ZBhLu
aeHkm2A2iOvReJmlEtkYGQl/XUP15Gu5TTISQejWbFpuyPCZzCf5L7b+1OlC+v1MdgHbw1HjNaNT
mO3Tdr0fXxliU9vFu+68MnNSx0B+dgfKi51ZCGWuTFhpbHUdJtqDtf29A3PawJDKIobrXp/IX+1v
feqaGh81BrzlEy1pOGCpREFSHRBeqQ7gZRmmeLa0vocVYeiRZhbKiij8d4/EoVaFf/40+g3HDMt2
OCu/Q/fuqwWDqCCxd2844IubrQOQs34ovcWmIUg9CNnTkRLbWV23kFlzcyVlndFdp5nXKgWiMBkw
pxqcdVO6QkP6NE1IDjqZla1ryRD/gH0I/yZU1hqClXYJmViBQCqzCwFvDD4kkZJblRGdKP9vtXwf
r4rPNV3D7jFFdKv1dVPwxpYImFilGeGkUZ6zZhmJa18RCOBSpXUolJnXifnrcNhfFf95rnyHVnIJ
Z/s+88138APxGNtRCsCdDpTY6hCxm5p36lewvqgq0yGyYqhc9wx3ycGneVvq/qVvYWi3N1HP/qm0
BocIuqaNPULj43kHwAD/YhMZanm6dlz4txld/SaDMc+2pBsy46DN1xIRtjkYl6MTKsH2PxtKGr7s
RqB3x8jxU9CZ3pIzx/WPKylfHAvtNkbRx0vtWiAXnjK3N3ZeTO/k5zsDzrOHkY22T+z4NdhCzwdo
bwHHFXnO1/O+fRIUzg5t039kfHtTr07H5TzFEIgWjQprJO6OQQSlmQhsd8xi+BntXJAiLqsHBNxf
m6tlKlccX7Fel9a0m/PhEjjRy5W33EnFuBCwtb0PLmUwpdS1gI51wAkyV7giMn4acg2npT8gJkFI
x0rH4uTP98nWVbuGh/Obj/PvpELjZdk9dKgsj0WGHFy2iMULynl1B15RgUSP1hfQWmAAmGmmyxTm
Vs5wzYBor0ulroJHxgP3eGDlGHvj7IW2qaw1HbskhwY+1Hcze+wYMm1h6tZ+dUkBB/36yMegs9/r
WE3jG9tZXLK9FEHaUYPmcka4bGocsWodfJQ4WX/8VxXIq6lzq/pdddyE8GM1mZ4g9vvNqjzUEQxc
vEXnKgpKkRTdMe/Jkne//lW+/QpRgKRTv7h1BwPyXH3aCEnqVyHobTTzuYfdTRaIItvBgt4JR5U2
Vpg6IU2RzhzYrh4j+HJtgR/1Et6xBDOxGJ1tR293sxis/2jT6jV2K5+EsHRiNBtgaPSOstd9EODq
w0r8UEbkNXkWw38WlwQBravY7D5lKTRCkm3vc3INF71Dl83iYdaEF4iP7MOuoV4CMcWgjddGxMhD
B4qggihee+gE1hFncyMQJ4O7ed7K0xZPoEYOguuLSf+5Hcb5F/62/cRw3UAajHlepOXg3o3naS97
hIPO/JQsrqRrAVBaJcG2nYCgcF/HBfcvJsoa9g+mjy5UM5BjkkAR60vjOA0l5JiQ04OOrMMM0Cko
tbE4BF8RxtDMacXDb2RSIKeqcF0hTF77tMBH6TZNmDpPJ8D9MdmfmrL7B14YzxonOWDATnyiTUuG
zuCczKchKQpOeX95evHDvowodcIXkoCu6gIh8CE/PUoDEBJjRGLkKjtMGOsLyZdD3LaSaFMW3EnF
93kdFLjGAhxNCwhO4JgL/Bwa1Q4Qkn/Pc+n1rk1zVjHg3eS50o8HrpPB799gMsp/HUG0LFwU2Vpc
LzZLIMbnagj16vBfd+kFzAC2tOpuvs4gfq5Cl6s4+folIwqu5AFlccX3AYCO2+zGHNeNyQ5z/Gke
jxEznkVvJWRywsrZPrjHazhkFq4OGaE9ivCs4pWFwpaL9HiJbP+w1sxef50vpTb4dSbOdqw5W6V5
afFPQDvZ4x+tBNFhlSq0pxuOVauzkKd4ZoHOsPV1in7UOJdm+Ighz+IgKJGlN3um39AZ9Y6kzcpp
8K3SC+RVAVFjRkSqjGspK7Jrege3z8NVn8Fx5cieKQnK2UO1m3IZzlcjq7oHfIVOGDUxQOqKaf7U
RYUjy/IkpSlSdmlkKYpEz/GEAqxbtD2Z4ChJfiF89z33rhiJn1XYTPvDXvPIEpT5HkzkzpYRaai9
8BptOg/ktO5u0MrXjmuiQfH/YBUuBmXgG7OCO4TX/Fk7M8X+wPq0WFUqp4IxPBDBD0TVdTsETwkb
+kUBN2uDjs0bGJOwE7u4ZilCPv+j8iKghoz8INwB7SvegqVABNgk/LuoCVceIYPKTTWcrXwmiclI
dVnkfafMGO6CAfHoUCE+EnKNf7NMH2j0TGB+6qddSasDHFUK92/Dte06AkFmoVUjUsFHsw0sfmnZ
42xsnESxo2KqjzDYgIQvyDh3GGs2gf625OERbBcEq6YcGF60iXUrnlXG5OCR5nIygkMZH/dwGPtP
psjZcqMImpdQmkXn6tOyaot2Tcm0ezfHqLlCUyij7ZsPbRWhiMKSLW6tlvuduKXydaR25aoGv2+J
8QaiwgeZVKpP8oh2eCmLcW8pubF6yxnHCHH+GoXuUJdxhIfw6OclJxP+jIhKFDqAxIVKBIMN1zd/
hHyJ9YYMzkP3Nb7SqOcGNdiojVDwWEa6ZAOjzOJIcy0PYTb+AS9pnH0TVkq6bnD1HRa2T4EZeqSz
BOCg6/jmVZYzJQ+B/MqtmMEGU6GQgRmxminkrkAMHWjTDixp/I/gD43mDymFeLx1xQ4fdsd4MrGi
wmNBsLNb8vNXN2dIA2yTxS6EGv+Dhy5TLQFcvRU1x0y/jL8FQjmMjXvvhAk7kIrNTkKO81hnY8FX
oyKR8a5yWhPW/RjuFPFKyjzOlmGsRPwC6dTbnIDRLa6kQezoXQuW/vOtQL2YnCn6YeUTmtXvUvNX
3MJrUK/qDZpRE9BQRSTeDHxAFMk5cK6RSxJZ3N4MWFgMHG8xDGshSXKbPQlRIMiukULHn5YQPUKP
jLrmBqzytsxBBTWHNb1fJ6/BBRyoBXm6sTqLPvh+viK7VSJQRfJCX45Dhq0DxG/XP1rqw8cR9v1D
qTmmFQH/L7ufNbFykYYrTr8Atwq+xmJJcAdjF+8iD+cZs4fNzexJTTeOj36u5CKIonVm0cvC8YeX
CeH1uXZrKc4jycce0HFDR2t+JxhGkyYxI96Hsnuyu44AmESDHWj88CDNnnDgtHyU0C6BUBKxbfIY
i74oF2jbVXAXCV8vlTR4u92TfcRlQ4OXUyEkwgXMT2S4QDNIZSkPyUBQyCXjAuDPcPmJdXYfWIqL
gEy+3+dZtgJr5Go2o7biIy+YZ/P84Wr7m2vrw6wxwcQxmS8yPfFVG0wol1mvytWNKxBj2y7Y1NJg
uImKed7TPD6bfGfHB+Hah1cJ664+J1EZuPOMqe4t+VY5mQduJfKRqVetuWYppeJEDpPoiH8fzGY1
xPz6cBR3Jw2tqS8zIGCBsNgyRGRRCSSCx813X+O3/toS725nL7RndFzo2/wEzgsEhKVyXOueP8wk
cMSmfx8PtEyuzTNAdpLZTixDTH76mq2465FYoZEDWOkoYqBTX3N2PAtYbcNzTnVpEKKOHxxe6km8
HRDLdZePOmVkZuv5VKfoOAePBEDHSTVA5R7Jy09UNYF+ucOyqKsg4Z1EO7Ewsv00TFXjvfapZpPU
tdzsNCzGJP8sY/vukWkqV1otuAlQsozN75EFTlDx3NHSnmnpIOsxM6En4L36tvsYE40l3sQzESlg
O3cvWW1QebAZ3JmbTA/c5JNvxxW5jPMd+iUNcbAoI31kJurZAImeU4N0gf5BQzJUhiwjeMM6iGL9
CMBWzYMtjHfRhQNiC8HDHFjMoox3Km4Ttl1zITizk1o8Kulwn4Dkj/OYjpyVk/orQSAMXXHaO411
Jv2ScgclSTCZI1c+UgiRNF3YgxIL/8ZfMl2b9MZ6WFYkAmoMnRu2BhTBb2jMr+kS+CrY07b6FAGh
gyuXN9c7IIc3YuMpvxKhEEtQqWvCTJzxgXW89xTrMb4qC/KnC8ks238mzHjTTjzBr6mhQGDkTU3R
rO060rOav66Tpupbc32u7WByMcc8yFq4Qp8J6oWFAwzG0r9So3C1t1h0NHmYVWaHhEtspzYadw9D
3LedpQRV3+cTgRp43KZW/Co/sD1Me+l9MFiOYknH9nIEToL6zfFl/aYO5TEAEvBEX3vWIIY1EW/z
UUMnjQY1Ugi4mrwPkMpZWKvEtxHPzN1mFjzJSzDG0jUrU6Euh7sJzndC4/pdo9W+sgn/FsMmYzeo
B+TKUJYvLc4R9ZS2B3p4KWESBaynrFaugTJ6m2SJlL/FMArrJegAo0yK6UivONpVMVHsyfBp7aSm
nJtuusDz/0nweTpM1XD+FbtOQAqHOA/zHetAA+e/ctH56ZA12eyIbxnQfAtpMKBgnOE89igeBf5Q
vvGESXzu226wCk4TUe2RPU0tL/JpSJs5YDSW6uNCAtI/H1v5ROdn87ATyM/l/dDHWXlDlIrZNvaU
nYC1ZmgIK0qO+bXWSDgUcKoBWDU0SW0X11qwabyi5u2qrBsLMnLGgFL1E5j20Xza9o1PCcFRAV9S
vQEEpTBTedL9UCTkSMbzyUPsI41+AYroVkHT9qt3nfNMBa8CfdXcM0A1iDF0h9WMwCXqByaSJ9pf
+73Kbk21HRRmRFC73Hu0wfde4s3k80yzMLYCHip2Gi17R+9Jq/F2W2k91gADmW8wjq1QA+U+eAg4
I5WbEPiUFPNViuhLAjoluySfhqGrV2R9jLvHgxb3VP3S1kq36sCiWHZKaGnmGkSnXfKyrdTYyWFM
4Gb6AE3o2y6Dh79NO/bL98Rjx+HQD33KJO3AR/Dt1e3jN6Om6j1oIZAABKaSktWw+lsjcJzlzi22
AfPKQLvsOe/omNm6Y45CeaVOFHSzKbkCPnss30mZFGjLYYs1B9i+xp4ZHK2W78amiL1pqyShieep
CMALnjuoSlbLz23l8NsydzH5vBawvbaemqBxWjFiBUCrEDhj4AuiOqpZL+Qz2cIkX2/hWX4wLB0i
GvGhQS73tfuZm9yFqBiQ1HJGyExBzu794IyZW5pu/EIVsm3vN01BSlrH0iOGiZxXGMKys0haQY4l
kuHc1GY0pJIB0o7g9ZTGnkfP16ih87Qd1SwAu3fIvNRLLx6RislwGll9mham5iYZkMghA0fpWgJU
ObgmPNssM3h6iLyNY1v+wX2T29Vo+BV798q5AqNJmlu7giukE90wqFR/0dGZd9VAaHh2oytOpSnc
QIqTjTRKbg3ylQgxEQ8M1CuimpuBKTeGWdIHof+wc0TDApMCLi4aOlDe64e5bO1qphyKqebp3eO0
qvQgc0gCWB9xW9xD0U57p4AL2LpnduGgOAo78CMm13iwbDdvwU86CMLkgCWwCYO6xBqwPlJJOQwq
5KRenVYRiBkl5uHou4D4yLk3ZYUry2QYFOWSY41DhKFHBAmNkiZbJQYAorkEOMzPesSvE17cNVVK
qN5C/txOjc0Y5oG/98f54OIf02941s5dvVjx9SIfIIwaY4i6gCCPIyTPBzXDMCbQN1PZNbDAy1r3
KulxOly1K75kw9D5RIZSCssxGZBG78nkRM7FsA0DH7WnRCfa6pKLwNn4B4/ESCMl+yqPxBxcmORP
VGaMuZ5d+LOnPakdxQGrM2FXUwVXNwtd2NfJeVqr4Dxdaz6Jw3Y0LhRPI/70ob+90dJ0c//9VkvG
XBeLoAQg6kHXO7DPeHGmximoFFUk7lEed4nzXpG+MTYVpDHdyzB7oPNxg0zj9aLZGMVbA0fSWOnx
GsmX4DdrWcQ5Txcr+cNvoE10UR+45sgDWctat8ib3609bHat1lSKSwIqOoaA0ftX7f5sKm/D0mAV
eCTUM6i/knFxL4dN9bYLfmYGPGROklLSVT1tBqDhMiluod8rGeP2LUh0+HQl6BYVsTLyLd2Fea36
5gjruCvxBEDz5w7nq7etY0DFjZ/Rjr/B3S26NYWf4mrA2cu50ZP44EUXy8LHS4qFdHhh/hzOR9sU
7++D3si6af5jLCCbn3IbuWZfAzCVhQttUaTD/nUzqOnZ+gc8s1qomd8PxVszQG56I9Pe2tZ3+RTy
Xdqt4zECByXRgRsnE17GTLY6OyqCUNgnwAzqEVoQwZPqIag7ue01Xa6uZ7aBe6PLyPnCsVNcJQiy
hvWeqvOfx28CbDJBTZQPrlrC+3FpcGwQ8DfIUfYDX9g7cDQXul/WbE0gqCDNVy5PlhVh7xYTLzeh
YjoSMiHeejWv6ArjGiksOoWvwzS6Dty9pxNElNCyauvgbk37eLPzXJCV5+yx4hVwBAZ82o22vkKv
28qz7r0cGjKJn0TE9FRghSEXiilnxt1aCrWpsNzVyfk3CGxP+M2zc2/9zXoXlbQqDOTel3lH2otS
j6vHGlMP013M63mPhjovwLUuvW7EtOBdLKHKEvXUjzDn1hKlL1GRBTwEWjr8uA+RVXI2paUNR/Xe
rYqlR/5fFEK5Y6ojjNjWPkN7v9ZXx1QQ0miZ/6PYcGNpjThxT7QjkXTnYCR3xCC5x7JWEN2/XrOG
bUndhKNGxNiWhhc0IRTrhXbBkCXlGqEz1enuKIWG7j57PgicQHqjiLDuYDboMVHylg94KO7ZoTf4
p2PtBtl0Jb+2jsUkh7K8q/qkiZ5mF8436eL6GGuyxM9F48i1Ru9ZgFwG2D7Vf8PbLkFZaRGFqfy4
fVoabzxHPrNbbyxeUy4Kupma0CpREjCtdPGWk1rvcjQMoWppiqwM7CpSyyQx+FXH1kEv5+NVfVBA
ZsRfx5A8+mEi8uFqbzVyIpmvtUMaKndkN3/IVQvW3J4UKl4dpuk3hj6xor/s19EHqXdkREsmieAd
IwBAx7IWUd3udiL50hXke3mX6/Cb18/PvdfnK/4gu7MhC7bYSFkod3rzAT/OBjvr1JaXPXzjBml7
anzNByaTOYvGOrOQ4GPRZ7tecWvh015zOO4jtFarBPkQvbvpfZAOtkvSNAw90R8oBxBuUTg4agMR
2Z9FBg1W6KOhVV7+zre/ThgaZWpnlOQYcWIeCeK9k+aLeCkFDp/5oPwEkO3YXT23T4Zk6pMIQErx
TuJeaR3YNt6xv6Ictmw0dfqqjGHuHC75cfSOHCiK7gY5lKoOZsXk2o0imJJ1wRVkdHW7SZjRmdP7
SN8f9eXRLGQYo4Q2w43b4CEiX19H3clLGbOFoEYwquz53yxirHIgCt+/pJEj0vYdUIjxghpw0pav
/lXKHxW1EWr716k+CJ1PqukqPgx9VpMKmbZQfTh98vZE8m0Q2g5uJPitVkZ3rygz5VzERKnFM7TW
jTrQcXoA5yg3r+kXksDX0s/NHcl90QeooRGYVbLrYiU1Y3S/IJu0HVwGgDyJKOAaEYv4l9EMolKo
s9pYxSytEC4aIrOMsNziUsW9AsxtLGRYcGtDUziCgAc4km4FliQALld3f23H+POotyi3wtdofdx6
/aMsGpvQ98u+5GdsXHMHk+Befm1Io9CsxbpyMVqQ7obNnWIDp5RoS2EQIyahQJet3BthZxGEQR5t
yDEG/8vRoKPs/1r4ZI/CnUJevvhAsAwlHXDlglv/fds56DrLB/4r3jAknYqOkLBpRiPcE37Ow0a9
wH1uxo4mrKK6mX3ua88hzK1tE9cZAtlHzl0cv/YWgVyml8RzHyWrD2JbjSiU3Sfq0f/BCGZiEIj1
8xBDl2HHYxypNh4qYnMDFSnPECMkCXsLTUDf/MbobJWq+Oajpdf/vfZCNJ3YcLuCaFuyBpE0jT6i
gnXudXf9WBODkgmCDqaZZde1TIG/K1jgwWdCgFaKe41ahcgnqEkUY1FWJNEJqhNflz6W3e874djh
95b8rFYQBNo//79Q7RfChnysmFZ3c5Ur8t8bdSmmrr+PxKwU3HBOFe4GzliYdiY86tfvGXAWq55I
KZVOMpmfGG61UomxyEYiLmNern0BiYm/uGIqsiZlEAlkGr2y1XBcxKQJiPUuDM5KDUwctMNPW4So
rgYI6oFua+lRTYKgQbyseSITdf36Gz6ESQhQci8f7cgJhK5MzNUyssXi/b8ywEngCAvVnftVM7nk
heNvSTZM3Z3qRT9RHGGn1tCJ/GL0ouV5kxAAUCOIT/tiXgUTWkgiHfo/ex/HbsL6B/83yZfUXgIK
a05S82gTv7sCBN6eddPvmKHaxCzUSCCMEfKcxcFGPoBMWoi/t+IJRorNKQb38M1tMmvFkIsf2TpJ
jeZtnH6Q2rzrKCCqg5zcQP6UglH155srPM2tQLZzt0vKpMCiegAwakqWG/Z8BY+drYhl1K8Rg5U7
lwfbIhz6SK6Pdierciu89DpLCxhp4rlAeLfmxeBQYJVbRC8BkEm4e+K8LvCLGGO+X5fDu1xn3PDF
jomvTgSO+VaZPkHSe+BDTrVJTuir6gno2gxmO/m6Z8SsMB56y2ad98lTtjKSpos6TnKCGPMVVZdP
c7JTJM0YEwCr0ABPDJvqzdOu69tzVd9r6IgY1puHqybX54sOyGgYccqAeApLY/PCYAHl35klCF8J
dXCpRMFuhMe2R6+ucCeORYt4tp07G12aDezi3dr8ylk2WzjYqQ393sDzAEPB1XsTd+1KwgJmY7w2
6HGkOP+E+3jUC9YetvDPL62RZdSq4OgTGaG2bl8IYZd4TzQO1b/u0KF9b5x7IARlkdCtNi2Bzrxe
VKGjnKxeulfwRSVXtUxO0nQgEXWIflVLQVKmliDcEoVqlJckAQSD5+/Z0MhH269SdbxMwX/5pNtH
Lthun6ZQsbnbWXOZhRlU51h06gxJltHW4f3f/tj45bO6TWPVsvhlmqLShwqzN8kCwLyxTJxEN51W
WAhgbNCfTyQWVsLoY2/sCigTFnTWQvU5YkfYyhQJlStol3bxXYF/xdgdufp4z+9Swjl/qNyykam0
MRdcB0rsO/syi38WTxwRxfelVgXAd+3ZvuoMH6LWPbxqS0LsRxsJnyb0vlcBPqQOoiCzSie3Ndfu
QrYimXQfTH2Juj0At2SkQ8VufhLNyW/F4GdVOol4HBR1woQ3GFhY1ZnTvqmbR8WV+vCGUIxNdfKT
f29qPa7xM1tnig5/gvimUpN6Aywqni0V2ItCGhT4I6ExUyxjXaGJXtu38HuK1R48gj+0067Ee5lg
21Oo4GJgYdiGj/rMOfHfZuARfmTlvC7GOPL8lC5OM9pO8whWcKSEQxGHUO1ZmdXx9Hylj+uTQx9H
elCH/QqFk89RJ71ezhq32aI9FwmVYr/DyK2uenItftPgQdoY0aERSAgJzydeevoQHNb84t08GQI7
51SLFWfyiTbvbHXbe9TjZC17Gr1p5uI6UYZfVB6KJ7j20IO1EmtGerJsZ91pwM5fltYR+WCtRtGW
e1BOJKv++qBXFC89brcwHwsE5oicTgrI9ckwWLPCXIlFVTtak6MnIrjMABcYqQzlEz9pLs3vPNDR
f+KS4bIrhTLOStcUerRA9/88CIk/e4WcuxsUblKqlGyh0nxlkjvOD0a49hQuFnUJi+UMImSjIh7c
jG4Iif82CfVWwBeMPkKqp6cnMqE8UKkHVt7Y2JuQFYfz7NkDTPNx9pOh6d18THod+be3gUMEGl7j
RF0DoOHcA7KDtIBprbkBpuKPS47LiqbVCTWu5Lxd+EbsFCif51w7itNkaeDNyRF/tDqnOBjgOlYV
tnznEpvRUUqfYF5MHIRTDMx1BLCthgRxfrojncMVVneQu6SGhr2Afz2PDSgbQBqesrMCJNqZ1eGT
PbZrnmbob6wmuzRImeNkk2mr6IrjY11XVvQOVWHgAK0dMDqloMXfR2mEXu2MSydlH1klNS6HQihV
obGcKRu6mZHpJEecqqxI5HO+NFHWuAR1C1jLSXnVUxFgWoKRBXMc7AGCZ9qkNDMgj3JS5LHm5FM5
R32YuPb/X+tAB1OiNjH2bmXloI20qMeAKCVvaKEfcqGjG73KlFIxBHEdbIn9DuYej9F2cICGhClh
DkJ1ZJpvmzDDF+niNoEyLU3r6o2tSB3CbBDVUIdKOMS4bbc3SEa5jKIYBNR3j9f07QcNyW7cbkWq
5RWrBt+8ULds/eud/H0cZaEXTzMvJFAIl7lkxASNRkIvlU0uf3gf6FBmpTdtZri7oLoO527glQBf
MG1JEGbAAtc/VuNmVaLrvj9qyERJ8a1vsoovsabAYuqpTQZ1aPtFohG29CVWmHsV8yBlRKq+R7B/
cDARnUVi9hy2oE1Op7hXXeabPQbsIs1SAJDEx4SGvtnGS+z4fLloJDk+5qlm5akEoeQUP2PNv/n7
S+To3yBYyqVpo9XrNu+eJVZs9GhNGsGI06YvGDVco3JZE5vJYiOj9Vls2Q321HHouf4F4wiVsQ3j
Ia7+MjSkOUcCY+vC9y6ev5p9bpMlkqiQXaGcofI+e6sQznYnz8fC/FHjucrRKdq9zGr3ZHY6peop
Vz+dQosXhcPTiTV20Wk4F0Z8t1AYt6nIvPHZlxIN5cfh9Ezu0VXS/Mi6Zg/z/GRXQNjlOueYoM/r
Lg+Y99tJrASEMgxMEPb5rL2u8XMgS7VY5d7UzLVSAH7vhq5rmZpnviwhInbl1vvxMvoXNkAQOrsz
kurLJzaVQdnPgwgLFwSxRwFyRjuljeEBXYpJ0B61uzIrAuHdL4fEZ8OW7TIhX/X8Otqr9dphQgqW
DSXrpoYoaHQTb/jiro3fhbW0kXQWcni6aNDsQNpneC9IEjY2ca4y0OAOFRER8eGcZx9VUOM1+Ge4
ms1qAKNkNVY54uMTzhiUgbcu43+zgxkY3jIcS9fsmjKGtNQq9akc5W0mgrofAHJdaxbYPDVwkwAx
fGQIyEE7NsZ8mGvhP10EcP6VshDS6Hemv5KvzJtF5smpGp7OsCM9GFcmyW96c2nKbCX49VJwHuaB
cNvGc59DP6vY94fZoNkqsfdQjLpHsubzaSmMZk7mIxvJ/+88XeoJ6FYFp/thm7g1BtDQEYONSW/8
1wTWzuaS11ZHVRKbCaZB+HkdNn1KfHct3XJ5ZzODwQZH/Z0ZLIq/Luu/VM/e6qjVhNaLJPy0vOUS
5PmtvYEFH2wO7lSq66Z48H4CnfMStGWlF2NTlKhRJjuVcPRiwB++bJhn2eQpJDR7BauEnkrWAbKn
n/DUAEyg5v78HUGSeJUwv9WgAMTvZDcwBoNh6QVD2DCkb5phl2dn7B09MOi2Tzm6owsTPOv5oFIo
vSNQrxISvAw3nfVqKHUI4VAT6eqBfXK4hSVun0poPnNOFkxe8jt1EDKEmGalDX9bwMRHo+VYM+4h
jtDjtdEbx9z3IKVRS1D5XSbeszCoeJ+QnCHLrod+Ngz8ebJHEP5HbRPjpFdKBnT7sy/9toa5M3Vq
FG+7Bb95Wu/5q00zC+aF0tHR0Zo5QLnvn8/OKeFsM4A9NwM1ytEJ13Tq3/7YNztVnnmnb+LckJVa
1ood3sgXm7X/RSgqY8yZfZ1DAjIbJQl+q1/OPe5DrTfMJ33lvN6zBYxZYkv1Pf1onz+93GHWeFAs
V+l0h6P6FvwvzynSJhaUi/pmnrV+je5h2OuWjGisMXj3GAoTeB01N7rssBhz2pBCgz0DK2B3+SJy
8vONkUWq5FqQK3xkJYP8bdrCl3qLkjqMK2b1lifN+brlqhavcxlwpqGd4Oo6VBoyzydHWIqWqIjj
NZ9tOUx7LbcQN/d9wgFYhtk6aKzrHs17p4+3WSbD86FZdwTwNWf+Qkk4p9I1qLsMnMf9btKIEsQQ
uyRUsdBEC3y/llD1Nd+DYe6lkNT02G5syB8IjE/gH8mAQA5wa0/I/sa4ri9pkxrsXK7m+q+LHuAi
p72ww1K+R3pkcK5FJgHv7TqtQ+1N77byzucXHHEWyG4rvHInL512AvWQhHipWGEqLq1STzX4TQ0v
V6z4blSTvifryqsMYtPGKFrpPKf3i/vNnC9rf70wdmRxq1mt/92S44gJ/HVqSfhPfzZdGkNomgVP
dY5gS8+CKE/B7lkX7XnH8zuLnLCjZqlESsLsZbzV+dpkv+EGfOXDBC5HKtrQX8Y+coSCsAVx6v0l
ePQF0fY2oCkWOxfwhYz+3JV+Gp8IQ7el1aFYESX0tHXmT88uvhfY1NeFrfjBB/VoO/uJblNmqW66
XC7/eAyObMdG8yMAgPjheBRPEoLALaa4Bskhnu1rt/fdxLgBPOZhVMXZRCoYfuj3RA8PXDN3d99h
uL2PdbGILWWkD94HQhAw9w+u2DGXrXGxsNvZUt8V9WEFUq++4h192iaNkKCAr6YNlLldix/PT3Vy
ORtnhe1fLi2TGcZf66/yrkUMMG6kgB4V12qoIKbvfo2uRS87pA9x7wBycRwvzWC8fbSkLeGjvRS5
jjV7us+kRvh0q1hfE6eA2PHIQzbOEC1GJFOTMRF71OLcugeeVnHIpzSY2syZ5AWPVWXqn/Ic7K+P
W1M2FIWtHlcxmbBzDKS7r9HZJFjygfGuVMOyaBn6bw5AcMFh6f5RURbHTyXYb7WWTKlayzX+6heD
3SmWDBW9fwz77T1cWuwDtaT9fR77jFaLo5GUr0mwET1ty3dYUZlE5FJB8pNAA4rxueQpjlIn0EA4
GOs1gSntils31aPrw0HdLsYwGb1GiuwMg4khwKMclNfyukxMz0E0PFqVw5M9mgoM5T9xwj4Dgzbp
dBHc8//9x/c5IyLV5Rlj9BfOyfLD6y5HGPywuMW5Inwh/cs6i/8HVRyLTCNq10Msobs1uaTgxWlL
H3d6PRdMTPODHvZNwvLr3Og2AODWydh2hM+cPT3BNGPzdlXNioHzLFhlnAYROfQ+kWFsUZEY66PG
agMf8CJ5Z1lqk2CWN4vYIRlC2bjLD6XZxAuKiaGFnMHHJnXneuyGBbUgpGaDCdSoGdBtnhhgRpPR
0b9QKFT2wT6L/5a4tSs/KhBRCtiqedQ9maqQsKtHz0BYwa51lL94ZZf6AzIssmkAh44ZbY1STth1
UMrGzFBkmHhlEwX3dRaSDmUpdQXoSIPHk4m+6G+T9sDZPnOFD55D0E2Lx3ZdztVzVCnk4q111ZbW
PEbJnINU3C+9dZ5mjR6e/pM1mkC07swkIcOEJnUypKhBPHwwVlilRRKrJpZMdGJxTRmVk5zEe1Q+
ABiXru7dUmPc6WdgoUdDJyxtJVFiFPdj2VZqKOaaMV6UJtgImT1jhjufAg1HF3n3HgoNrDPHL+cg
SHCKXs81uamZQaFL9Q+xzXmSQ/l6er0o79HNW+XhgJcWalKgTVTJ/7femz+8bckExTtcPV7MLiaM
TN7zUhT0MSHLkptURxw90PBswUdaIVPOxteQcGWUlz6CxWC0TOE7Bn+dM5WNL3bY8I0P76NmNG85
sBgxIjuocoIttkJcXdMMJAFC04JUoXnPMW7XG6qoDk6FFVzYMHGmEHAaDYydzuBwZLXjb2W6lfNw
k7VBqWihZ0iv5NIHb8e/ctnqS55JpdFPjE1GIidvATOPc876Jxn9jKRB9mkZdrezAejcL1epuSPP
2XrvQrvihCATJ/vZLvG/Z4y8xmAWJiQ2W+HwVi4XtsTvzRp0WpSRS31EqCgKd0MLph6evIaBu+fV
OQRPMmbTVc9lFkim2HhV8Jz9JSUGz+u6Fw0NcAOqK4GBaHiYBIzllXPa7GXM71YAJ+bvd4QZIcrn
5uMbGSaREH6j+fMHWYoqxqmo+zzg3j6KM76pgstp9N6q6GgvdM/dLj8Zxip9WY8l5y7GscNYQgwG
v0AnAzyVCt5njLlLVs9tFQiSRW3gzDCb81SZ3SdjL+nRwK6JIdzvLtVE2zFqo2SLRgyI1eXu0l4J
infAjwCGPqJKzM/21RVgrJnG9jyYFK8b/K/XQcrtHVIiLBhgv45H1y5eqdnTIbgCcKHsTsIyqxwZ
PgII5m/0wsSyfuulg7W4pzamoArFJ2538P8QsuiJFXIcEXFRTqeKbtq8InsrbBBPA9EfyXgHJCku
PYsLW8z1ia0IhFSE9mL71p/nqOXHLxFhqrpASvNF/oARSLOhQeeMc3NsOExoleg43hN3JLQks/ZS
tjGWXOTyJUyJQhsTg+jl8OmnA8dzL1TG0Pwh+Of+lDXnO5+jS5MRYPalt41TgVmINuxFO8jT9a0g
EH5IqSiLFVoKXmitXD5WDZuTxKQuQBfl02D911RW2OyldTdef1CQjCjT9/q3ua7xp9DXg+2Zw49i
l3JGF5+ZgwMY21zkdUEI916lR6PICfruzhrScvGUp9WW3QGooDs2lSwCXw1Dn4urRZxcjFa4fEqX
FvVVRUnMwJvpmFOF97jvfxwpRHjdEmVDefH/E3oYDRdP1g633uU2pHTmqa6HbO6SdGr7wrHacfcB
XvzWlaHp81/Eo7nfOZ0vFtMeaH+zXZnquWCR+jgby545+eWqPVeUBgWBJwlBkhwa364irC/4TztU
wY9pqXtO9hqqnGqTTFqdG9z7uR9ZciMSK2GHYZebVX/jXhn/P9eW4w5K0xV15EB5wq+pljsEYkUm
BdggEqJmK5Nlf+9dKdXjstY/fBkSkEOq78v0w07zolP3c+ywHwq40A6QfryPk7xGKEe/YySpRNIw
w+9M+O1u/zyreM1giLNzdgLS1nAuz0z74gxj4kuzNGuL5JRu2u6wNLvP1j8/nNUPFqZ3BPkEUw1B
ch4iEquC1HGkLuhg7l/hsb3moSu1hJJxTc6XYfXNfi6+lVhiCbwA3yskTLm2tbs9Z/E5iOSpXLrx
iMaj5E9JzAxcgAQZWehF/CGiLxfvxGjtL5zZW2AhN49tI8C3bK7Lu9svE/TGgKqxFevm928dTDXW
9bqvbT5d6/mjPAiNI8mhcpY9LsL3TaLjZqtfGGQ8tGlkEoIfLig3UNHdBdgIkKB200jMTqGH/5jC
istxmxA6UShsiUe58gdJok8QRy/5P/yvoSjOqkKJrwD+QXAM9Sln7le9h04xFVE+0M14CpMbcdmR
0Mo2mGCFYWl5vsTv7NvNE7UP7u1KKJW1yn5v0Bqo6EBXH4K06sTmM1vIxsNEBWID4Iwen2hp2/IM
pQWTAo3XxNwyjuJD5z7Vp5y2F/Q/PiRCgHzhympLmb+w2Rm5bXTUv976P4kw97Zt9polh0hcgjxx
tgdFX23HvP+DKAG6Ep0Vc6EEyh4E/53eTSLYlCzTTJ+jkDS91c9a0XFOEsn1d2x1bOrVSAF2Ip4I
exc03XUlp7XHUKYwR0MkWNfyFypRGtcCioCv2xyjJey4JYQEaIH+9NvWZC+G63vWfY3BWEhPiDIQ
s5Qs/2RS8daMvz0YeYT0uoEq6ENXdK430WL7YVSGLILLw5SoLvaWaHTs8PKZtfa1OmBefY9vlmZ8
jS95iXH0spOqArZarztpE9oIpWkT8ybU6x1S3AAGLxZfzn3L6OoWjCPMuVWk/ZAOWAHxtoAIfU2p
4wO859ZMidSH0hWz+IHat8hpfxYB7tVj3Q2i5yd1L5l9BO7Qf+GlXmO4//kR3Dq58IxF9hPK0CZs
XDIx6PV9lQo/qYGfBCYT3dnEnKFXiTZailab8SbpoRLZoljqucZpdnHQsVQEWx7kGB50cx+ZC9kq
GFnooGlI8U/octqzF+afwETAoeV3/rsSmzpmjp52WpurmacTl3i6xKj2nOCdztebu+DiK4oRw0xQ
kJw5hIhInJx9Cg+3w6mdN/fpE7VHDqO4GzRmwCVqPpb058liT50c1/YTLt2+/wYVEqVvrB0ZMtdC
UERKfn2y2lxzvpoblTDtmZWmKEA7DyxpgKy0KJGtfk9EEdfT/rMmUlMsjRpUaZ7Vq6R+hLwEQ/Nv
3XJfP4MV5J1TLqzyYezB+SXmPHQ72ZITzedHZ4Ft8wA+W2gck48xAQg33ifiY8I8AWYFOT0hgNib
UfsxDY7gvKZ9B5dHFtoaCSXvUuWYSD9YbammFlqhvl2FsqNk87Wy6qiMi9NyjqSoE3z9JFLQZ/+u
uvCXMoj/MprE6XBynFle54MJqfWcIaVnZfR7nFRWWSmGJSiM9aLNg2NCcobsEE79BVnQRjsXTmcF
WC6kC5WDXJ3gcFqwrnx/8cksrb5TPtld9X8PRTm2FiLICnr3Fz+TB+2oBqsR0a+qh+T6tARLMYrg
dGU54j3ahrw5uL4psBxO+ll0n2fCx8RDDsXiXeg9w8w8uHn6+mETw92t8iDVf+Zi4IQAlW+J1k7j
QRlK61AvOl1KQBPmRkr+LjGqb25bjvMTKYx1ehEZwhJ+YvH261IQDfIAwL9V0gdAyhY2fGcufe1I
nhujvedP/XmCH22yXn/hXoxMoBVqCVla09DSbDP7qLnSsw7HrzBZDIxtRC9XOdsx87tx0AfRy2ee
/0BXrU1LxIFZBOCBmDAe3o47ucLtkXM1uTdD6KnFAVb2xUvUUwykpait0I37dOEcesqaU4LQFeE4
ScubhYtng5sxjnLHWFHku466otqdDpdBqYEJdDiuBrzjttu30tltS9buPgqhLpaItSgvOTeWiHzF
1750mmDyeTIcAaMLYjHL6tZsrQZZT1clza2f6pS1Qu7VulMtJyd6Q69dG0+mGVCPIefpjaUwkD+o
3317+H/GcAQteI0Apf5jzv05abH+i/MwI0z65SIWqrxw28rArEOMhn0i8RHCdMle4w68sDCz8x0o
DYnuIBm/7HP9RmekbfbKNERSkq3lO8nfWXXeVBMnd4b8rERTaWeCRmB345D2NvZqZjs9cEhTeYBR
jF5gxoWNdBetuiYYMhyp1SJxrwfZ3iEO9VFOLTE4K1yLEtkLuIgiDt87pkd1IUkxpQXMl8YdXFyw
/M3HRQhFKOtCtEAwlcOexbtE1WX341QUUZ7WY57TGO20VJ8I1QPpwEZ6V4bJkVI3o5rmDKgq+OG7
aug9ni3rk/sCsgtyL+sC0wKtS+Na2EnDlMToSQYknMBqWXNpIhtENV43hUTolzhkqvwNT07tghVD
MDxaiJ7CoBDALbWYxRyEZUleVFBVg8KmFni6exGIL4TbDmDz1i5CGsgrpbZP1lWiVzQDikn6oCVi
nTlo3nqOoDnX6qrQkYddSenM80qFptZg3t5AInXGl1urrCVzOfXz0Cu+o2wat0TEfxqyIVoTVutJ
UPa74j13x9L/UyRvV+O1v06wdJ8D90BGx5Uv6Uxd+/C+1zy0SOGu5xvHYYyRXo+uT01EXRnc9YXr
JM/jKmmKNMYStF/D7IOCUqU+A+6pRRTi1wledl/n6szPWCvTJQ5NYdveGTvEbnE4JO2i14wrfXXW
NP1ztgCJe9x0K64xUVR3j6EvI5wUFcbZFiQsC8PVwBpySKzcOSsSCOtPpOZw+YfqvFaIBTHK6a0Z
dxj8K4CD5ga6WDPFj/sSPC5DsBlFhe+kXV2GlRKS4kLuyUvgq8SdUM3AUBTdK0FtV+VLPivyYCy2
/T+1Ejxw9TWM75H9Y3/GkzVtgFA5ehG6CN1q1G6oSjZUwOH5xp2ENIVIL0f8aky6VGpXMAszw9OV
YHe1Ngwe+V+vNpQQ1wcWNtGVIKnRYdehxHC9j4KfpBOEP1zYD3m5wEBQeKbhaMtnnjizpiDpMwa7
n2YGP+EaqQ9Iztcgv4D33kN2DLLUkoLAzvY2oIpWfPYvnpb+QsilWdQiB8seczYOouOECMBTzEnv
6rzoNIeusPHIJEXXqdTk4Fp3augrCdugVZJf4/7F3x54AGbQi/pXHpMRYvh1ze3ONdcz+u1OGm1o
92oK9MYRYzTiBv3QvsS+OLmlNeUsRivoiBrhuIravq6xdUHj/8hhPZZ9Rt/Ww7mgngvmALgwIJxo
3+NozJa+JuTKrpf4ni9TwH0X4zDcTVzMs31/4fd2t0FRTl5ytg0X+Z3BOXjv8AGNHciCNG6FQ9Tr
FtIaibmLfvJAPZ6bp+goc8CH4R/EEAjdQdGDamNs1f6YjnKL12b9EqTp2ZDKjUCLI7Ga6rM1i/pz
qQzwbekaoUMRRghDykL8K7rLDOgfne3eRIt9exP1NeffBsztNPnzc5koNkyk/9HETTJgS5nJ+K3v
qO3KjuOzuMC0X7/UFYi67wFYTWd/zvqq41cYJBE6mZ44kuuDTmX8M9ZXo7eY1ob18eIYqLWAZJpl
YU6CnbF8LUU7XOkWbQHmsc1c1jZdO07ooJkH5sx+OeJEn9P6XK3hxk4DlagHqI8bDtNa7Ez08g3x
lkd/a2ARm7dLjhb+bLrxZ0LfbEhuDbJFGD4L0GW4PBvha/4TIPotTl9atcXf9OFQpm1n9g0Wgef+
8vJB/KwCkAUXZ2L1uGEUv0CuWC7go8TxHvADlMNBZEGAGHY2mEM47IFN+Ag77Q4mWVCUWP2kR+yL
tQmJ8BxHoOLsMDEDhvgP2TcBfv7SN3rSiJs1KMgfnz9JuwPNx4ZgtrWtAqJNyFOaqYXd3hh7PcBP
uVRQt0WTBplT3QS2PiyLeX1/TMZgzcpIm+RwXykGzLCCsbFO0a0QdLv8puV6s8WarZCyemQq3vFS
gC7VL0cAAM7d8nUVo+0jcnDjiNVDt6Bj+yDb8ncbHG4xoiD45uc2qSAGynNB/OtMskXqk/3p46Pf
c+mCizZ0WHY9z3lLSQFp9jnp6SLGFW3borjPvJjnYYAt0WAVul9bzjaf+lOt68hOxCF+IwbrIHLv
08IpFPH2Lg02Cef54Akdh5hh4YqCgHPs7qCJPiyBFe4y6a7VIB92D505tTP7m97teB83mX6rGOR8
8qC3CPGmbdulluMjCv5rg56xuwfX00Y41+lYKOEpDlOT60P+CkIxxH4v4Fd12Ubuj35qBh2fPEbp
c2mPJP6ZRVOD/9s5r6uXkxQKLUg0lsCObvIhc9IgznKDmsGcy7nDhFWOwXe4MHvX3yFLJRkj4vcN
q0+YqO7BC+cSECsF5Hr7HOTg7I5i9jrJXAGiAJIHYAsgM6GyJv2ZU11jRna8Oo235FC0k8Y2Boxt
yYDliguw3laedS8zRyqxyJelkmeFmeKVitXRLnduqxVfRlJCbgA/Vw5qNhcdUK+kiVxipwz9svkz
KlOgr2x+SNQojjkeM1AB27KySn3JaduNyKbt7mhukckJU9f/+cTHJ24lH+Rt2Ims7Rw4ONO7EM/E
pD9K7LGpzZVPM6J09foVEhpqylVD3gipU8OyFvbREVzZ41jz00SBaAtzBkk3kCMBf54YqSrJyvUD
7QU73XLULb//wsesyJ/GYT0SmLLAz05R5vILOoZTk5jmBMfkkiO9HK0tJh81Uyl/uhYKMuAIMW3c
JIUQ2Fmmwncn0sqa4RJLpw9P4EFsKLqHGf4mTqt+VUZd3U7caAwwRCJlLZpnIiGlz7Cw/IGsbs0w
zBO2ABDKE2hftmkjoWr+KBBl/oEmkwrACt/CxfuOUvp+a0BKRIgfoJRDrQ9wugvKHAOVKlxL+ah9
pKQvLfzlLp19cQfN0cX7bHz+Zu0vJpFRLl4SVRHqJzb9nmxSdPJwQZ0LwJuY/0U4QWAYrnuE2MpL
YBDfex1/g/6W1Pqk/FWWlccEUHXs5ljVGIO/5+AAik8pFQW2OFsY5Jm+bxTUn0jbvzRDwotv50fx
pvKc+jlYBbjkhDWPK0c/iQ8Rq2B0rqbuUJRcpsdk4p6vFoLK30JZckmzQRlo5xNMCXz3Ew4bESy9
rOdcUkI+kHmtofKgAz6GGfNDOTAm1gd8fHTag2lGxQNoYPhKJr/HbumpNMPCKbOLvI0PbrqpJ7/5
pJxdSQMHFiiYjPTo/BLA462a8UksAepryW6zHP+aJV9Z0zqIWfHYDIgA8pu7/W7jeLMw8XF/NmPK
33arCoU65mWGx7j2IXvUvIyAIRQHDx1B+GmQuSmYUdOczKfOW04b8UFRzszkPfOrf1gdtsmAXMm6
Zb6UIIhyJUQCirD9c9Tri8FI7k9x0vXPL/HTzjymiBoCieWuVPjKpLpx5B8IXs7EqSvMZ80V7LWq
tt6g2E2LzriJecIaNq01r3csZ7ju837/2W2PJfq3YmOudGIf9hSFfVTW7m/JCRi0Y64wwnUP9jPD
paxLEv5TwSG7KJXGYqnCGdBkNbdtkQf2sLeO6fLV7Vu6bpZZZZfm+StDtQTQcnT1PMfIPadwrcfD
Jzj/pMTbpcSTefuMP45p3q6J3aoVESp1dYeEe42t6l+zp8S5a49WDvMplJ1MKVX3BBfosBt134Pd
HGvfxlK5RYx+2RWXlXVUHT6GOCGTu8ipXlm1xVo5jrXnTDuJxPK/DPrKqaQ4H+/sD/9OjXXVSiJ1
pRUl7qRLDzo4jROQOhUugWXmX4cVqOWjhJxs3N4ucesR1uoQHKgiX8EBfe23MaPT5Fx0FeTfQi5e
yw0zDBofn8o/A6lhzoZw7GTM39HcNAjjyugHxkswzPoIqvw3NIMYNWD3DrNTLxkLMGiDjngTS69j
+1iSroWKkfF62Y4UdshdgoHMBaKQxZFDPHdELl+bYhFz1aFLlkUaQVTC3s59LdWEj5rSPPKmYgaj
o/T0jonta4PmjnVpAJfdFEMqnikYPsKCae9PysiR2qr0CiDuASl+KaaE7xLAJiFFDf1HhnjmuXdh
R/geTaCTJ6t/fG2A+Fnr5b7IqkntLxjUFbYro+D96yaHsZUHaKrgIYiDdW8cUmSJHSGQ0rOvI9zc
W25Z2qQmKlDUKJdy8A9HJs3fR3919baH7Q/mhee4cfReXf+rjSvUnFjxaTb0thxJNqi/wI4AqqU0
81nweujS5zpVtz62V27MSkHPboP7ieaznR++wmPr0XjpaqBHk/lA2Z8l+8MtL55s0MxKfilE6Yjt
dmMiyFgFLYM0VhS6YHXMaxb6dvL59ZWqMRAZi1QC/TCZkcx4qSm9GlWZnb0BSlHH/y2C6rQvRg0P
dy5tkFeNjH405a9Lb8sGzCrTrDNMzoBIM+u+8GnIlMnx4C8SIrfzYsf5cUF//bsLC/IzhvWRZlpv
HaolgqjlR5TAp+GBeIfiQLaV/MYp7C+nkdCgd6d4JJDQ3vW2DBdxB0oPL23mrbYBZtLacBgmqjAY
V6BiyGVKiF72Gm6KZoBuuRsQv6rLJ3SMAHYHjo4yPHv2QCEItPlV+n2B74tehIF88JlHD419tx9T
W4Dmuo4Fhpw0sBdu0AP/2ugJgNlhWG8x3MoU+pCTFEX0Kd86fpVtGCndtvBG4LZuCIKj38cl2swx
cdcKQOwn5noSc0fA6L+t/Wj70PXoUESFMSew13A6nzNqTUyqhXHLl3Duw097KVi1Rsc1BdLRZswZ
67h7RiSgHaUt1b+H1QfL+MrYvV+W8IdtPi0Ecr7XRsdoD1q2btmeM6bRlze9EfZG9bJU0fPgLYmI
Y+Th5KZoVOWtAiDllX65wc/km4dqzTWWbvaUHrCzAA/jO0zMLLSEPYb63C6UVYTfyY3wDKefAF3g
DiMLzTi6KQ02nJ5Jr9Sbwb+uffIQZSkzcaxZ+zgcU1ldJmj2RgVcA+8PBfGhMRTINTxw3IeNAmcb
8LeeeaGExtJOgVG/gIRv+eqqASGbT963Nz9zrgIF1WRZ1H13lUBti4PQAMa/twq2teKG73nhwhCk
IP6Lovldw+zKRJOz7yYa19exTcLmjOp1390H4a2oxcGw63P1vZSU1zlwZj0+HY/DHRXvdUSr8i39
XhTQAozVYZ5SwBrLyTNbzsOJjNpsGAhVFRqqQ+OOVV9anZlhXmC4Fy0HTHyMGXUcpOl/SadrHw+2
DR1ge9z3JiSwAm2qFsTZTMfwDEJnBdkD9vub3Rr3VIawVU6FFty5RfHaz6dyVjGHDZrNKIa2DyGT
EKYnsbgsedtSCKAD+FQ6frzw+Edx47uUC+CgoJx97cRi/1mpCLpvYgJLrEPOS+ObUh9Fa3PCMS4W
nXjHG8suUyvSNdtKYpH9duiAWl22KlJN2yxbAVQh7d2oEdGSeZ9kUCsrg7lkR7K1FlOM6rVG3mco
mptqNBhGk2H0z17MvLCPERPqRXRe79U3pHXKzRTbhMEkZFsCnXpdNd06PHUM8MSUQibMT6Eq0lq+
ADqeD5PxLiyejRbU/EJ3n1oUT3PtcIhgSoeUdaEZk7E1Q2lv9XXD/1slXPmbyFzEzbfRZ11Kpcgf
Up6hz8cT3xHKbaySHwzbEZIYZXVkNqgJs/mrUk3TriQKo4Wkpg4fMJN3uupLQnRmUhogniKg2Hnx
v4908QcmGIJpKit/pvaD9Am+S7CAmRRC6bda4dRzhUD2d7APEF0G01p8GmrsXqnc6J1n/koeDW4q
p6tLBmWySTN5hO683ZgbIpWSQJi+1nJb5cV7vdNgY2kxe8lkwoSmedFaoajbFONAauS/fqd7Auvi
5mtnWvwzkcoKwe4Qm58cCI80vAG2B9qnM8MTlYkqQu2yZ1Ryq5Rw6IsmyLellRllX7y1eZ6F7xcI
lsN3tL/yt2JTgq2qczGA37eFzuQ96D7p0KUbkP3TaLJESE77Z195A8ermQNtAqPaSAnaneXaIyhe
SVH7aYj7PmqsRy9xi2fS2g0J85DMN6wKtrWumwbsrj8qBwFJVUZXs/MpkvG49kJP54/cL8ymIv2+
lwmF8ufFxittEZ18A/k/zIuOT2oitmvD/j2JFyxzPkMvyN7rkUJaG2dqIciTfwLBbFoAfHn447WN
qzJvZY27rSA4LjR8VBrCFq+Bc848FgN2WDkksbGTbArU8L5JjoB6hvMzIjTQcWtpRegdp86fmsO6
tjCSleH7veNkBXFlhNGko3Gi9aqr/+/xfCznxz2OT4KNCdpVYYFCSjvz07/jrzRN0ixrvhx3cdCe
7qXcmbZ+WOuZC8w3Bx+58DKnmeO8cPe/MJ11MAck6TmFKJ+OGJ5JMB8WaUiOJ/592r8Yyt0setT6
b2jrBQdlVYhDlz2PY3CBnGbqAF8ob44dXEAxddhaWwsuwj/YJYyWqLZdLGvUfFS0Eay34eMscCfH
XW0a1JcOvy3HG6jHnR66EsHR+P9EcNNaHrDiVG5kJZOSTWXZfefcpdjgq+wHyrS/Kt/tkRFoE1Be
6o8RWw3kIxYgdJnPIPEqaA0AHBsdbwZK+f/JQTnfnI61nlpId45XoK5QUvh+cX13VwHlbcRgLrv+
0k9B/32Z5F3nqTE5aIFY7eBMkOSwdZ7WCX8EY/imwQgidJieO8ADTIuayh+4zyYdI8Heklc7LFUS
o5iz+dSb85ZwDCKg8MGVz0N1hnRZGWdy2EzDyMs012EMhOu6j6R4kFPdDUDRT4P4/FeI83ZVO3Nj
NZP3946z408Kk95qMnaV9/yw/mvB14YUyuvGAhUVXL5RmhJ0Jmh82jdbdtfZOIdBDFKS2QpI5q3a
F08ybtrXK6ww/Jr9WnkK0SIvUNLHHFsdzBt3nTY80qy6J7SPwiJvZMoJb5JJiZti8vMcS4LkwyEx
RhzS+45IYloUHYH1yeU/GlqD2ByzAujpUbdIPlLt/cuS4ov7mwgBGcq6WEh8R+PlNb5OnA1MeYQY
dlcCwIFNqXTqbJpDBuIboa0Ha9aGYGiCytoCzVh+jSivKpC8hzT95USsVYjGzud/jfXAgPUjTR+R
+hRkhXizHwx/kEcfroaByWNahhOeeDp3MfSUyaDkXPWJyG0b3Cf7HXMGSYYUecgEHRhKh7Y86XeN
GKnEO0nmIZtC1+L5t0D377BfkYanJL3/D89FouD43nIXS25crOJ0Int625LoFSHA2naOh308AHaC
9m0zxlsEvu6xhrHs7Nt3DmBt1FNb7o4NIDR2B89c6Kypk0KHm/ZOI7uM+mCD3rS4TCmUpMAoeOun
AeI8wtJID0RPWWcufqjWBFiwTxeCvg/2nQkW2oeG8g6xLTDV4dn1aqmSEs6RTvUsShRcBrquSIOB
dJeNtxupkdnzzMxGbxaeqrBo2p8tz7JhbEEEur0nlOky3iGUoakAPLEVeykFE3F+bV0mSW31qykM
qLDPkfZWYP6VLv2Je38EWHhSw8jBSIWEKuvntzgC/DZBCpomULy+eE4oTL4AwghMhNtLbopr5IcP
hes4744R7l3grF7vXjWZIESWIf+ZJwVhSBJ8MXCeN4xSlIwBv6TYjiQ84Qav0snEPt6hauAB3roq
VDqKJPNQrk1i7WCZCJXQ+jmiAa1rBnrCFc9wK+y3uOPWAIHCYPhP44NVT4J0uP+5PIwxKXrUvEBk
C6QAOveVdyU09ws9coZ5/PhuJKg12vr1MQF5qJ3gxcIofPe8KGsGPF599X3bewfSr5+JZc0TA42D
GMo11HLCz8lblMi2jBKQHWoXO60r1lVfEa/Wv9l8F7elsj5jX6A1MQgrG/ocsmjqYbQRHxYGkzxI
yLbbaxDIhwSxgfDyyvewMbFnPxvGNZbmmEXvkvYw0ZNs2t0utIdl+7QmgaH/i6VXQ9SgNOFVFk2L
6SUA70Tvleki97VYFp0e4msGTnBFBr7x2C5+L9PTN8HJWe2q5936okMY+OR1dEEDX8/v0uQjZUkH
cEslEkvC1AOgFUeL9H+q31PeU7ae79KMODFmj1FO1za39ePo3vlj5SOmea1sivVghj4XZ7hJCs4s
pGdbjy9VcuEwjtGZRQv9gShf9MYWrkJ/dgT8puYcFLARdFJQfrrysd7nOz5EqixLlEYiFKX1a5xC
BDHkJfJ1opYYXrOS8yKwl+W77bnAJlIIJTQymlOQ7n0p2sZIW+InVhFHDeQu9i989C7QsJr5E/ZY
6yaYXIIOQXXa6WW9/2is2gcLV6bpkXhOi/GoejvFyUzEf8c99j79DAFN/IQnnS1smmCUbB1Tyf9i
/la318RBIq/ST7xyedP4U5XMkbWfI+54cSqa9a8AuC6PSMva4VZM1Isl7WITlYVIAzK94UYLAARw
yylLCEchscUrjx4/YVSR2klFE9UeK9t++GWj2jGTaVG9cnEjR6PPI0KVDFUcPaUu0wnX83qD0oCA
eUaeXS4O326IBCuVF/IM8azobzzHAZ2lQyvBxRskqMtqb1yyKoOv3op++HaN9G2gXTKax5HYIdM/
OM4me5uIU5QEyQYn9LEf7HUzU8tKturdSpXNhSgptbDWU/TqJZhdAHm01eCXUQh32bjrPA2Y/s8z
Mb/8qWsA+BpS9lC7VHNnNJFMB/sZ8kmmUbYf7/ypH7GxvOE1m5rOlXAOzJDu2mMR+18ualP8KF2v
hWQOudTd7Jgvj8fLIEX04QtZG8Ghdm60K+n5nX8/G0NI1Jvn02POCNedtBewp0/uvuZQT1w5RFkR
i4QbOOXa2vblvFUUMbx1oLw1qQnzFsLUFfEwsqxBV3BT0+fe//anILx0VvTSuG64ol2jXdAw2f1+
fwbD6vqOx4wBI9EWiGPk/3hgXLDM62hK6+7shI3Xzd1UA/qm5mpzGDIkfPmGa8a4SK9LQI8YMW5e
vsdcqm31wenE7jRDYqNB/7FfqpNP/PrnjuFjCX544X7tMY0HgLkpYqcwb5k354ugw1bFkPn1pAEX
/CtxajcLdiP/yDhaOMTxyi/GEro5+SuaKh08LJjAlte8+3b6FOOjbGSYG3M9QVw6f1Si90VPWh1n
LQjy4nSmOLuKi8X8hM2q+66z2yZ9t4Fsoyd8F3SEkLIdMd/aaLotuC06vqYvX0PNykQn0DvRjL3p
TkVC2iQ3w0TT0JP9n3cjHaf4G1v3ynXz5qXKJN7sbgm3GBmgDfqWfwq6etPZhgMTbX89BcK2T1h0
lO4W1401rQzuHHCtAIcI0jHzApI3JiXpY/PWpmOouGjTnsyK6r6JuuP4QJxqyFQ2C1o9fZ+Dovb0
RLh/gsKUAcq6VR9YrcoGjbL/MiZifADqaCU0mHrHHMidcCwLCg4ViuNK3MT5E6lnGi0w9L+jyjqv
KKDqrQv0t6B5rk8pfuwA4VTWkvXeW4DEWf9TMix6OWkyC3mEIGiFIYLWQMnMhuiDYeoaXn0P5FuG
lE6FulhDAzz8TD9YWrcE/g1yks0081cnZsyv+BRN5f4gAWyP+Z5ZlGVBJETcPtlDYHd/zMR9BPnP
vJjUTiRsKEstJ4lItg2SyKdmgANpvnsoywHdAL0eo1jBqIE85TUNvYmgqxVj+9wae+Yx9PY+/Kds
yotVZOiY6mw3Wt1+EZ2FEGQZw1KIIgPGO3Mro5dmj3K8iQmIhH3/KSYjwToIKgo4VMAQ+7e+EKVJ
/EU9Kf7h0uSc/AsFZ7pN/7YHNMMxfXyUqC8GdRORlFgx7TCf1oqKQieXyLQhBZoxKFz+N7fo8/l7
0kpgCX+NDjN5lqELosnefk+MwmfySaoG0kZ5Okj7OksEzwp/TUnl81i6gvFE9O8uQLIRvdqPGioe
rMdgYTe+XAmlc81Wevk3G6456JSe+H33gM0bUEiTO7VlqC/XUlMoeIdygZXRLxMXBt8YOr3JOUOn
L/8vndzfMqTeqPb+u9xeDW7x221vtpKN8IwzSfhqBghJBYcxJ3HdVshOdx7HIRVfFDgnds2X06jp
+MzNRRUXouOr3ctpRVh1MpR2yjP1Vi6KK0n8gnqHMpCCP33njRBXvZ1iiksXAxhvxOGZl89yAB7z
m7PRpaFmuPF9n0getQ0QAQU5FT7EVWcZx3UVvfdCJpOdeEU56zz2ICWZrftZidUeGzy8DN+YvI0B
IBBaD32KSq4oSCAtQ4u+/L33B+od5y0cZpuBFRPGcCTcL5q5kzaIhrOOYor06LLGm6L6fCGdKq9Y
Iu2LEWhpNtzDKoCwquMtUcrvJ7nfEg1Cg1o07N0snyeXYFHHwPD2XyXg5ZQq/tRh5YFGcszGBrSb
cWvMggfVHnP2xHOwt33Px79V+LxiMr1Ihv3mffM33FsB/29VDfzB2DfEt/C5gQQKw9c5txPtVgc0
LWbFVP24r4zAlZIVR6GUgZhG6y6xwOKFVQAoeg5yljwbKII6JPg2JHPObdhI8rTFdsuFX3DXrrcI
rp0Mh1IuvM/DXLYtkfMkoA15RAHRh69w4CAqoCgpxJaokU0NqhlTgFW7YfhW28pde3HgNUBEYvyp
L0+aywdNxN0UJme95N2148gfEn+62c14lnoYuAOlaXVhIGcA21avI7XsK4TpCfsq5uHgKH/mTfSh
a+70ZVCUqqpgN+Yb38E8YoNx0WC9pFrHqczeXuEGURnUQQO94sCYF3XxPezEPl1NJMXgzRa8XCwC
oB6s/yCokQ3d2+h6jm6CNwa+KqV4AHLDdGgR8ec31fJeKo7xtk+iXxl5bSruWm0KsgX/YRq7tLNd
CvriZHJFFAv6sUmAJnXC0Ea0bObdN9Sig5jRhTBGrJ5Mbo/+JDMt/Kc43hI4rX414IUYmZ3bvavY
gTjUcdBKM9ZcR+FhA5HTIHSQmHCIuD4vf2ZkyVe+hZbiyqsFagATnYimK4GPcMcEhHkQIyq1IFLM
4lB2ykUqQaaGnVooKwrvuhZgmBxS8g4Kk6IeqaUK4tZ/NMf+YwKq2zmw0WDyb2H1mX+kWyX+K2xk
jnVEvMY2QmcFL1ZieXofDgEy0+BphaBoY8SR4QtkujuOPjh6Q8Af92rFT0bdWdpr9NoIgVWjSatO
Pi9TooPn0PnyFTBBtwuog+nfpcszbGmswzn+bw5K843pIhw7IGMjLx6WoHodusQq8xnfxHlrnqEt
aZO7QOqJPJB07O8a//646SbnBFZNu6kkPXGN8ZwGxaYfQKSV2WP6lWjJK0pzqoUdRxvhQtOD0VzI
Pdadx74gaGSFJF1eF8DFl1vnVp0lyJzPoyv9w+LqLpQP/75WSyY3QcwMgRBa2DevMuStjQj5Ku/m
XMNt7Nr4W1XBqIwdk0o+/eSWrDhRGY4taCIC+W7052aw4KbPmnul3Z/WecHccWouUxqAhwY5f9sN
qCZUyQn/hMAXMi85S/Hx/jOtjt82F/nx+4mYAWGJVKeent8EhOGn52jKgqvNjoZ9f7fwgAfV4ohG
+F+kQ7ma4MssSPLRxkvf3hR1O0BpEquqIFN8OuI1FDQMRBE4wCU3KhrhD6TOcMkgfzy+kQGYRgqK
mD2cAeCWYaQEPz8qgVutfQSsXN+yoFvKnqXamwaRUEFfbN2l9vqMwSZxhzxxCDjrz1BDvA/U5LOz
FHg8VuYHUPmC09CqtWTpgY4axa+qtttZLsL66OAnal4DORDjvApiyCmYXpbpfkIGaf3xkrnHknKw
gWjd/UnvHNeCT9B14NZKQ9SfWuJWgixkfPBGh2jGcAlOmOXjDmC8r6TNIB4trdzWakRkWFjwGqad
RnRQnl7auus4z9zXX8eAsxA3NB3IP8OVeL6FmW+AYXw+TAlEvAZnnVFDkRXCYPlmX6ZQnaWnJ6Aw
JKemAybjeF+gnY48HuJwxMSpfNPt+J2NUyDxePaUf7CNUGSXaTva38AZpCaigwA4bLJafHdywizP
a0CQgTLO1Gj6zEepr+iCuerr9NIglBAoPT1PSiF7+9BMI91Kvq8nHitb9Wgxg6AkorQyQbAcmG7o
cgehq/zkhpVfbiHYDr+pi2xP7CAsMsIDAlD7e869NLwtSqg4CnuQJxSrxPewdF20gz5EZhirKNG9
pruYl68mk4ME75upHb1csp2bS6cbbNkg8gzK4BcOBCnHk0o/6wx3mmmJaEjnDuOopFUM9MjjwHt2
oDmKooZf1OxTRhr4vqatZnsfLGXekS+qv1XdYMXNQPQSTcGIc97KZvidaKgtu+QzqKp5Urv2dvfq
aSZuqLqQ9Pz4yIY6GEw7n0bgG18GonaaO4fu/gDXIj8/BTStweK6xpF9K3T8KPhZzjYPhyKXvONZ
s2ElZzCIKO/wtRX0AIuoSMUhhpQrPh1sa1IfGIhuglrDG/DDrI4Y4Vs3JCCKsWD1DX6QsDAmVqMV
Sz2Ei9MtEF2QYzr5acFATMWkFOnIIwuTvNvUXdaOabJ0aElNxN/GcvIiMggvKQJ2I+dQ77WUbRQZ
X++QIR0jAWTA3AJAXoZFbw1gl/SSa/VPsNp1boBbfn/90abj6Q7/imunp+sD4cR2qUPPsUmioEFe
LlFQUr3tWImsQjRnjrQCJVw+1lNxniXOwLueLXPc+S05pvYuOTt7Odm6MBxDzQm5nOQNdqrwYA9S
PnIIsRxqN1a1xRx5QfDZTejh1+mwSDOlVDkPgvC25dF+rCrdRlOTrCs2hIKHI/bA7qyQsQJVwrXg
9DOdozxb1FdJxidEJq3mo0nGRAkLOO747OOJpb4rtLOn8MluzFoWoCuuZau6DoLCGWGLc0SOsVi5
RWMTLXFh/6xudKwdpSi9Wk/LekoWnZKYFCFN6ycHrCzVHD3h9Wrb05KKJwJkrGZUa9N4DXVtiFn+
RdeWC8eRuf/uFieGhVs+P1EqvONeG0rrZRforsCjdBp70KQFLvRV5EKZL7vuFhGk8PBaRr+c4ZUr
savptKUAb0Hln2ut+R6tjfSTHdU+DHdbSlyMbsyeBEmHmOd4cNwFYQnaXOeyF911THkyEoj4RXeZ
ZycNLv1TxlBmi1bY8cGwSff+/v9H6rG1pGT5o2fbr2sJ+3iXqOq+n+Pc7t+qrZlvC45OP5JJg5+D
fr1sPPsQBXKBEAJJL2KFQbWZFb9M297NTrJXKYJ3TnIqKkA/BYjjZggUKlc5Zbt7XEmCjnbpToGq
r6XTOWGCblesbEY8xxvWyU+prw6ttGjXIXGX9U2RyZzO8IY4tF6FFYgwrPkc/O5pcw0eBRE4XVjy
nH3DJDjEteO0dV97zVhA1vbod2YCmEQta/LQg7B7zNtBItQFIlmtHGoNbDsOtzo3HM39bjl+eKdQ
+H2MgbfaCwNhryla0zuiGZuHaIJ/wAdUzFkFRLecA1w3GlOJr8/mKKf5uECWr4MIYXv/AZ5zl6to
Pnh6PEwhUe/SUd+dcZ+6Fn74kCZ9XuypGIiPmXZC5sm7Sslh3OFKIEdI6E4gDaCpoKm2+8QtHALM
0xWe8lpZRkPTfsWWZSiJ6eucuzTvQXEYgDNMkya/LF9HaFY7LWFONhseOdIcUNQmSfWN/zCdYTBB
cT4L1NlJomK2is6+RBrEPCNhBLCmuoFhBKpbbz3xLAgGqmB5wu/DcMH7azIUnDSF1p36bw4zF/hV
DVSESUgkYeRxjyrY3WkoWRjUeyWTMyvbCnRbGoYPbW2BUUUMY8ATdV/OIPqDJQf4q9/DVnf+fHEZ
b6J662DaBKujCYR5LQggKL7Gm26Yy1VuhiE3J+wdBg3rKqS2ynUocmpjCVspW2KAb2dQAz8sG9HP
vtdNI1lf9RKVfwXWxUQ/tes0Yh89xxkwBVWSAdxe8q73W9nlvfNJU25AHhpXHgI153MCK3wIAszf
gZ/VfqFFaiIxSEHY5fySc5cmiZh5AAuia9NYShg/UokYY/A2C0Oy6PYb3Lkj9/hsseR8kCt08uEx
7DAzkc6hlQ3bKO5RJ3o7tXWEMBFU5+EVPeF94orYrdXwEYBR2waE2TZvxvrJUokOn/x0fXqBvnDT
e9nQLYrk5E4vrNWiWwfnuBu8mU0fOvb+nDaNYXIeE7wJqj5KKJPwNwyZVGLLk0eJi2QG3S7JskC4
OxotQCaysPyft2/LdlTaIiQI3jlhPGNghMzL5Ber8t6bRaU0Y2gAoTRagz1VdUZkPe/kz3ufXxOY
o49GSPO/bffVKgnwFFmMJh7/jOlr26VSHfX1oo+br0vrdS25lOAV6T+YAaC75zZXHrtNPwKvsZlE
NfddU36QX4mmYcOiiPsPynPOl0PucERL9kXQU1gQcnmt6elu2f8qEpp/twB5Y49r5Kqkce1eBE0a
UAhLxxyBIHZfMN6lk4/Tw4PhnBvYtK5xn+lE4PhYHf0xQ3h0WJ7vS0hR+qaZF/oswJO1LQxUqcMB
WTtgVUSJAHZ7bLavLR6PjcDvomFq7F3pnw9gpQwHbuRQ2wWmVf2nS8wc0jNse8w3tQknsFfaY8oO
2Vyx3X4fwW6vVCtiITnjOqwcX8A4y9fh4RX+KKbfCW555UpaTGGNX9LBbknWJjVA+1vuzRWW51L+
MmZix7VCDgsIFlYKw7HqUaQGYdDesixAk+QJqHozJWbvDBWCwYL/2/2bomtULL9KGnBhPa3N3wEE
2X/2TdEdyNFzbM4u+ipOEgBNDpvJza45fWjIcU3LKSSnfdP/oWZtrBhTwtTl3qcUzZg1AUJwezY8
VnWIFeDHozotu11iEW7MyCfgMPpW6Mvvp4wwAT4w1GO160Gf82bbA18WUfTvd7PlFG3xhDGx3zzK
uyBmWkza5xYEVNZZBuYgcMRdpqJGAqPapOb+/8fxFnJNwP7phpsrsPN/PFIchIRCM1G5IbyBJbbc
we+pn3vr5mprL/7l1Bwkuo00BniS8/22QvrGe7TqwAj/mtyHqxazRk1T44GE+YcStPdNMoUFlqcV
mjGepv7k6CtJMj6zqAAQBM29Ny4G5a3wkHosTqWhilg+6UClnEsezggeK3hE9mbcGzAK9xvO91Xu
19EuQBOSIcOVdnyDqXVz22tWuW8w/337Nde8uXQg8/A3P+UBFKX/FKz2m2mJ8HBCkv+/oGDYij2A
8wFvcFahoxMDI70TzYRPT2MuflfZZulpNl9antxAVszI5tB/4CygLxO6kIWu+R8DAzGrjrW5bXpL
fKeOhZTPhEuNe+i/OfmvC6SsoYQxYVfq6oC+LY5KgDFC94K1geyN+3dRoNi7y8iuVyyvYl3BjB7y
QferAT0A3tnlnCiHo63gJxV5bpznGOKUvy8i9ubPR3XkvvtcRlVDH54Sx6Xef9AxjY05Tiqi42oD
+MP07MV1M4yqiEEwSQvuRJdb+7my8Fe7x6h1SzSAnxRm+81nOHQlt5eorgxPSVmnwjTFn9H3hLJ0
fXVHYhmJZXPOFmR0rRkDVeyh/Hj+VmCMoNkVKZ4cnhGr6qvEquCCdO1x+6QK6wBU+IvCB32cWoaF
gbnO4avQGAxOpZDPGNOiijOGTSYT6LeYdnQDhdTdwau1PdYL25Zt/YJ+xOlntqQjakdVMDnayGMb
bfyNuta2dEiqLdPcIk7/4kCXhPubCuZRx1tAZiY2AP5OcUMuVZCDMRnwGzt7PQBdSAvnOHJnZKN+
kn8Z+V6Ey3hJRHzSoJQlr1XNJml4qmuapXWzoPI75odw2udYnOqolQP9smiAnqlTf1bnS2LbbqZb
X1amqyNDMZWRva461h+0N/kHIspoTJfmIjRVCBDr+0TpQt6P8EypGPJCEJ5dv/oAX2n4Ujq7DvMR
ANk5aSOol6qMjjdgZxMArGoBdCwnZ0Xdg+JixVqwfJ/J03PnaAfv311L4OkH7k50v/C5/3pdtuBA
Ydc3w5zBvxuM88/817/QkPxzs6Xd5MYahQz1ebE5a2NTM/Q+KwlpEpCMFQTNf8AFoIlCbDLUCurR
X3vGI852Y1LsRYWANeWO1/s8UYWSuedR5TycNqILlGSrMUZxcS2ow7hCJhPLRA2b2wOLYbmPCUaV
HONA0hH5UHa4Rc7ybCCXvXQBohhb3UblLyrglTKHcqn97trSUfZMXGhkPV1pcCY/Ns9Om3rbooES
kVJnZAMbhyjFgSXdWJZNm7ciws5/kNMxnKTqZ+mOs8x+grMGqFVOGrLJ5I9BdHJc/Knn8TGkWMKP
MKJWfrZRcQ+jYtK4q79nMe9SUpCGIid2tJdh+z51d3eephmwmfZwjELHKiDcTYAEaA5OJtHbkUNg
CZtRIvavrRFPx3EZLoocXroniZHfEYKiPfICdv/f7mHs8aeQb8Hgv/4MXCu9duM1H4Y/ZZDMDiqk
XE382pQlpkJwZjCy5hdDlNW87Fm2vTml1y4nIvO9MTa0h5mx+y01PFUit/7JQpKfum3P8u/tYVZj
jJ1dUV4l5A5iQaW0ZfLLZxCP4VmCbrBulncdRCdOJMP/HIVPdyn3VBUnh9SbK+7lppEBzDNX++iA
uV1EodpKbj03ocPa53j183I/LPb5D2V2x+7OWAeTthlxWa8ga+uVFDWezpUxQXflRwXJw1fVqJJQ
Y34BVhjf0iRiKANOi+WUPa+Fnb91Suv0mqYKYPYtHpRz5ngK9G6Zk4VioMkhGzuBrf6UK3zIwR0L
TgWCtZqgDQQlK2f9WJsxR13LdamArr5waw7YUn5jnngur5nJxXyQ8M71r23xe7h+1kRIgibfYePE
zAyjgy9Vm+kICTNBhk5MdEs+5OOXbAuYmWAIzzv1GbX3tMIZL8+UpHNWll1uq02x2OnfIiZGSf3Z
pHyOFZFyc7pmJ4m9kH/dkYh2ikE0/y3jIYu/iCV0ZIqOO/v7zRPLoIx7IBO7n78BWgL3xzOUi7jg
dMauotPFfNY37JM6DeX6uDFsmzysbe8C0LgKbO1/AitZOT/y2ew7tYV9SXGR2MiO42peXE9f6GBJ
czUloM2gfwvmj4SzAxK1cWvG3sCCHSeaZWhVKP8wUoFZLeuOF35PcHAkt/5sPgbkcYptxcFSg6ur
R6aJVH7kptiS9MYIZd14z6dveqMj/63CC4g52YDeVTGkclZNkSl/TDOBcNCgFSrxAmKznNASLG42
/xkF68M4lwf3eiuF+taqr+2byHee7hzpMozv17fEGn+82X3bQLHS2iJh6M4HB511yOOHH6lJRlhi
Mcs7oFCq6ACUl6JK4Tzm8HGP4hu3hDYO9upa3djKB0qpxWJaId2kp4xAaP0kFo0mZX716EFFST12
AUoeFxGRCQgUFzKtSQDaUzoiDhhkis5U2OzdKx9hTTaZ+OAwdr5l2KnkKROEzLmvAWOxX3DvTLHV
ymqWbA6TFW6ON05+BqULSTaleNxhA/7fr0zUdyds0owSDXnfl2XAuJqGF9BuQY8CDkRJ94yeC0Xb
kJGWxWWgItf1Pf7MdS/uyKP1MNIyzlAyGf4a3z15I2f86ui5GtmHXptiWNLhtp6faYViLxR2MzaS
65lrLMgFE8MpP3s3ZP5fAFy1tFkzYsBhT0Qmq0BgShy/FGPiR9rsqu3q+/E0T54wGfMFHuCl7YAn
e94zcPlEIPW52UkShjSTUKfQMVwGm39V6mpj8X4YM7/Fcu40ogeERYzBNEMQ5O21zv1Qo02qEtfw
7ol9UoxEj8zrYzrgQbE3SgmiLRdsmSgjr1QCVUwBTEn/DcZU3LVgj27D8pKhgSPpjeBZD7P22IFO
KTGJHWL9V7fRHTWvp5N1sEWxoFtOtssYoYWRkLoesTeHhnhGTdAhzUohA9GiTPdBCKXGBnhKuL42
vqeFOpI1ImKZNWkpe/g9yLM4KgEohtp3HgvkqR5fC23PEQp56ofZ/hlaJunEqFHEi94psjLcFnUX
gp6puep4+Nve8vEmrLh9uWY3ombqLVhMJRCgpPxnl2Rl8oXpBLm6Uzcfq8Gvc2FjqP+V3PDejjGB
R56BZOg6FtziTZxXlezw6LbqZIf309qaW8I41MnG5SzvVZFbb1pDfTXWgeXLLdJfmCVkhlv27gqS
G+PAXYwX+E3+dBRVbXEGiOxAl2oxSkbPfNzUWLVYKwsCOwARn3cIeRr8VSumtAZAnq3QXZBd+i6B
Z3dAHoO83P1aDNBw6t/ELrvmWc6g2OUX7WzQ68cPWUI4fLp7NAbUABimfzS9gPL6auEE3XOjm882
efDeYzJCElseCHbHdRG4mo3iXB99VVUHKvKntMPNueTSC3wHCbBiN6r8YRKe6YhDxkqLJuoqe6Xq
zPp7jLtzG9+I4wfgVW+47o6WxVKbOpNLxrV4I0IBIq/+EqSAWmYt3n2Nq2QLmziQbIDku5OUYFaa
Vt97sF2Y2rJ4pEHzqHbTj/d36VPsnc7EgjGVtnlQ1ixHUsrXpWYgJrvU8UjB3Qkom5rwgDwIi1dM
bWkuSU4ibrQgO52+wqxbJdI9OCSLWSVXH5Pvuwvy+4Li9WMLvMIgzBF9v3ReJ8QvzQarXkIs/I2t
b49wG6fzkMCwH/GsXAGy0rcfhDrU+oquBGE15QlAOReZ4AkklZ4mT4cRK6EdIhAvBtBjPCfF8weU
XUvFsUAZEHj0NG2MjdC6R6xve3mIr6DYyhcrOzICXNxSpsR9kXGXs05bK6mvPf+s81dBUpeuBDf1
OuKnWlb4k6KZw7cm7B/83rQNhZY8+7nCLQodhJV4LnYyGVD/X4rXo4PSMgJXtCdiy8DTmdpGhU0N
rYFLaNzHsH34uKo/f1mrNPLmqAhl+byg1bWYe6puDoCh3qzFZHSqa3CCp4RInBEvQIEDNynNHJjf
NhwwHASzFabiwwIX/vRYSE2ExdnasZOHMV5Y8fEqT3N04YwaRynIHVCnOW3nEr+FCJtIrb2T8f24
tGqVEM4zKtLSACYoY4hbDRn8shuV5tIkyzG/dL9hUa377DtieUZRPDD2VJgubW6iztk3TfVVpryJ
EnMAPfOzIpQF4PenRkpmpE8aeJkgJYQLc9PgPjsQNZT1U4FmE0ZNuUF+3H8wwdsJsudg/oGhfqVv
hIp51tkipbJ1iTDH3YruK2BWw/PXZVjDvW9+ve91lhAkgVxS6JjDGqil3YWc7gfQGs41u15v8892
B2/XGBWK03o+wpy6qsSakO14d0c/1t+swj5fpDL39F/BQNK7HN6xNBDPo4f7YKjDSO+alSjLf0BN
ZNlWreZRzzvLsLPvbb2qRH5nK9j2s8QPyOgJHCdVB1/0MnUVrS4Cv4jMEsaWwXJmk7rwItaay5TB
2gCb9WaYYDOTc3jBWYm4Dx5EPNSPEb0pmATTjAZ5N8g3bi7od3gOaUKUYwMdQmpNnzV9wb0qzt7u
9Ycbxdk05kP9FYdgROLrW2AaxgWoS7k2NYl5NUv9Yfa2S20lb373Z1xx5VfGgoDm6O41+i9etac+
ylPR0hur9VckB1T3CVaBxc5JxU6H9xyNgb1A0gawoHlS9MwmOhdtL4EpNLp4rClPtW2hFgjFrdoB
yHXRGj69beI+XLrvN6FrpUWzKMN49+8VMA/mx396K4E7mAm1dy39WBu112QD/ctqk+opzNXZVNu6
7rLgD25JpT2vfDHi3mzrc1zlgqaB/EtfngN7dIfs7OWt98hAxAJcKio2PltJeVckYg7mBqucNw2I
ao1771EAzWWViWWNv4H+HgdxvIZZqWRczI5an+3u9aAQIavjhdce8u8MsysXgHB02N+HL9ShM9TC
88bzS1v1rOJzAh+lJIr5Mtbj/KfgKgXUAtSOI20BroYgRFFKUByAbHULSSrP7tQEeilzBO6y0cwz
njo6gQrNKOzxj8T+YTSf6OdktNW11bXWfJ16coesc6KQTUz8HaObwKx2CgLYZ3yRQoXGu2HbOVFw
aS6XklwqfkCfJrLQPfngUOj1W97HcqR/+RIdxNA7//tEfDkpPRapFtgrgccKkHKPKCru3wEACqUq
dWAq6Gfqon7QQWGMzZWMbhx754eMnvyMUHkswCLBr6P0l/VweMkfr7C+lazjuh6GgDpmjGFnNx2R
57YYNrJ7eenVpRH+F3wqhf2x49Orx4HfkLXGTmNkKfNVbZ3WG5Qa38Dkf28fLfOsbrrGzXgT43gF
fnVfFo1LFTHjWbmYxmkJymla4xVnWV4cHpVoAeBOrf/sSn+iaAkLowitl6giSRvyjYt2wgygOpF8
yQj5vYW/2j2jogehnHHAouoOeAR9uafqX1UzIwVKHjK1cEuYdNR3uzZD2qjUy3Xg/Tf2jfloqCTj
6VHmbZh6r8JWBI1psiM9QkgEElUAYVIP7rranYQ1m+g/E5L5MWvFDM4uv+gWxUSpNFt6vT2ttYTu
TP5036GEfwgjgq905DhD5UPIjEsYy9RE3KfzDStgDtTlyjWmShHuqQIcF0pU/gxmdB5jVwMPiBEj
ntaB1m8ffIFh8+KOEjh3sKYGG2L1jeZZABUesKPQZulgzIShzO9M/U9z0eqn3kzIg69lIx16gY7o
nrD1CyIRPoctMjDPqJRZa1wyMNOAXQcmL1lmIvmKxsJNRZ7QoMsljdcNhMo5TKsVizjo2BIkQF8D
BqHtmX9mjdLHy3Pyka3HFmeS6JZXG04biTPVdMDmS6u6mdrX1mqieBmC4JBNF2iRbWWFbEqxU7ch
znoRUUVz2/F3Q9xmDuDmD4fobGfJRjDWKS42Ov/NDP1BNW1yLAAjDOuio2pGQlgonB7IlM2XDYzs
c+n3cKALmR4gneVyTa8o2IuOk+hkasqoI4kmC8u3RLSP8LWZcJ4O6zOF1MacAbu8LZycFos9F84l
N6Pin06JkKecTLoJQjV/aMo/+A2GW+6ZdOyZTrwAb4mQnxXtuhA2QcIqg7gSjINfkX7KxFdkbKnY
IR/ufnDBqHZHG0ltv1ZOOSB8o3Ps8Qnm3CG9KU5/n8ow6OsSpwJy5OzTXsWwgHpMIJVCk1ShOZ5o
rZco1LRpAVuf3sbqfggH0qOy90pr/Q3yb0oAgzD6KLGzddp9znfyRCnf2/Gtrv8L6aYzaNiAHJhr
lMpPTFmH2OkutgRU97Sy8Ov3rS4pJ01b40X8juM/EyyTHDPj1Z5BHItP++zJPSlNAYbqWS73rStb
wLxhiJk5Bq3+pJx7Wf1URas4Mv8LJ3p2HGD6FXDuus4/qMvgPdMWeHTNYLcpVh07BTb1AVzDU9Jz
mkoXmulTa5JymssPPg88svNfIhZudNyNAYled6dVn4UqvSSYfdjXeXghaXlQXdHTSqWmzeqZZUCs
EnssYNP2H0Jy0znZ3PNRIxgp4ihUPn2l5LlG+yoLnUeb2jMroZac5Ol1Esj0MedeqOWC3sSI6oGh
V9zOGw9PosWY038Gur1HbAnwpuNtvvAM6V954PIr1/wBSlg+XrBROAu9SI8jaiPn7kOMflZcUIAS
NU19QFouBbwaVrj4/lpH2JZcSI06rgJaTg2Gp2sPd+dTUV713v39htZxZnKou854LQIkFBLLJRY1
QCIAh57yf4pf8pInHvH5M81M6lpsEu6U72/zZfLTOdXT31us/WFEu1Mfb9hg+RzNbaZHNwdHZDJm
R+nxHQqGNZ3AIHiRezZh5gZRZRa4e9h+rMFKqXu6y+CFSeJYINOllDxK1DT1dQYl9sd/0iqRIHWC
7WoxVKS4i/StRDmzo46aAeio5wmKTQ7DFwp/Dqh7h6pk6pssPr6afHvVlamA5d5+tt8Klr65AmUE
8Rt77VcCC7U55xho4MzRzCR20gP83fT5eZI3R4p8r00rYFhgYV9Dfo76n5RkKEVjWzTI0HLvpGrd
x6O2FR87sX6sXNDO19gCZyii7r9fcuCMc7QFSAM0/3sq+dmKq4BYRtR1JoIm6PpXHBw5Tudm3Ty9
0et3tnUI78O5um63difFAkrGOfMZKTzga1LqZcMLmuyd69ZwWgeLgiRof3+aIqC1BT6Et3T3+8N8
4WsrbUSUyB7UE6N3HpSJmExJHOZ/8O88g6CrfSTmaaNzDB2KKIVvBBXGHOSlzbP/FzqsioXd8p/w
qmoyxxywxmtz8eJEAtK1SHOey9r90zbcgj7WBmeCUkQcgSu5ivL1coYFvvmDQsP8vEmKolggumGf
xMRagxY+3GixHx66YP82nz6u0DDHIaPSl+vgXwBMvF5fMokbicUpkDwDumpb91D3cNKZNbpc/9Jh
ybhSrKY6eolvIYOVizC4nw5f1Qbw2RKQR85naoEUBsiQ5Muxc89yzNbZZXbBYBRwxUZrVTg2CU9I
fiz/xajvkaFj3FsLeXH/I/JZRFLcpIb0iDySFZe1PFuDWwl9qY9kYkBroKiQOypdHPonNOYGMkfj
rX8cyWwyxOv7HMf/dCfavYLNW+Iv22IhY9nMWiI6lI81BIgBigRq989Onz7W+H6whF9FSQ/rSV6p
X+02rWn4N2VX2d1uXRG322oPyOCZx1BTxKjjtaHPSzxOCUCk2Sf37BpJtQnu0FgaGRhEMmpWhHt8
IMwepTIm/CjRxZlKxhMdi/pqGLz1CDGiRZPYaqqbt5KDFCkNPzpZvP5DUwFoYdLpyZ7FBzYrk2My
3MCLXhZlnv3VkR89cbZZdnnRtnQ8EskteCzL9xt612oCD8pkZ+2JJZ5tW07NotlNeX63MG2eu48A
WnssRu4UY54DQC+pvgUKS6cS6xw7XhydQbiSDl2bK45h6abpvdpKveS6Z4Nod8Y3aWnZuS6rnKlv
Hqskc7viCmRMjqStk75ouxvOcrpRL7mgJjNoU6uWnU/+VgSTxmjFl02kApTFsbzRB5xqx6F74KNW
EwyOj22euPe5xIMCtxpQJ371zmAoOD1/Gk2W81LyHUqbEjhslf6njbK9nnaNDTBjBqdDNoe+TMeO
+lCaj80GFzjPWq4GmNQEg2WPhiou7LYMzmWcvgy8JveumMkX+4sdrGThuCmmvFrwt9BMx/bxYfcQ
a3dLhiNAz55WlBhm0S0APwcG8zaenoyXahXoCaZlF/lzZXzdAJmZ0dIMszPzZQWuDu/9lXiRGMHD
4wT1UNSAnrGWnFvNV30E+4ux0QHeCxy3/bbRfm6PSshJ4xu8mS71vwxFBxiPM5caKmb0NXngctob
cULJI46Wyna92mCmpN6LqNW91kyxP7VzS0aSbQvgLd3AiyuROA4QlaDs3ZmfAnelkokxE8F0gk+L
EnR1SxZ7CRoLXTK4m/7WyxR23LarXlwh+S1ECBwDciMOOnd2qzcdDzWAIk8FMY6CKH4dpOOQNmw4
Gn48j0i9mM/qtqV30ZlTuEYWqlk6HKRrGcNKYkFz3MLH7H0FEioZ55wygoyUKgum24kBcCMiH6OX
o94aTJKFmu+atYWKw/U8q65D/U91fzzuWIPxJhF/DCBpbrkaoiNZLw6S7Zvv5cDnKzX8WNGtOSGD
s5PyOgU+nLCz/ifdIkbaEqgb3C6WaaZ7mzU4//byGafMDMkShZxtCy4oHaQESefnUd8mPb0Z+9//
GpKsWSFn4j5SyRU6LcxVImsdZApe8x6mV2S2qf5tyWzd71U9GpWzQDWOzBbH49LhETOf4Xsrx4+1
8DD1dZFGxjVPtyTJl9p7hE8BAffozhwX5Yg0pIwARXzZaRLEmBo1dALYOOujm44M28bFBvAHB9aq
POlWaoz76xhjF0lhh7E7SmnioB/bcCzIslVpoElWWCtSfmlEgZyX+nRVW4Toecn5X5f9flxDuvgi
+lfFB+55uiDTtipLs18Qv4DBjqPEmuEJTdNP8XxrOz7IQyAw88/+PlfLWS3II1eHSMN17f2L/toF
gkKtFGm9vPfMpB/o2j1i3XQReHfNWdspJnxBygfFh9NBkheYFUMVQwIGuSGP5I4J3F7sezHPXu+o
wasoNdeXd1uVSUU/UR1glxuX53VVDRCYB97owwBAcstQwVeRObcFyVuopvNvbHiIY0YBUr/8PRrq
6v9kvZfT/tc7fmopWm1X50biVX2BoNmYo6uDleSMKl82TfcKUjqRqYzYaYUHvBLe6ybdbHRnPMOm
9GxBqGZdkdeksyfBQsWhYwmUtkjmXS/58Odh+BPxdaC5LgBH/SY8lnfDzRnwe3LJJ4b5twiZBQD6
dAFM1vyjoRfWOhdLj1857jiZOwnxdom5ow9hQQKytmM/DRqi7fMK8lVOoariO/4CcizAvK6VyaRz
B7DJw7IriUsQI7AKcUFyTLu328VoV7eMiTfiUtqYhbRnwogJRg8R4oi/D/SS2wIHOi7BELzCdl6R
7alQmmqlFJk9uyGNWvDftLgLYlLMA8fzcLbNUhFyoBUJHCll0NrI7kobgVlBlnW55NSIZTUlvmNX
WYRt8vRWE+36/FSBTliA91SZC7nRZWNyuScUTZj3ZYlEONqJ3hd9DbYoGcv8H9gsPZxtJIpH/xAz
UyqhB6qmarNE0TFtvZFbCsbn9q1V4V+0JWf1h1QIM2aNHTOl7r0a/tg2x5RvFVkG/lGMHFaaRKFx
jdu6dR9QFRppopP9LpFwaHQ8UVJiwUKftI1v3F30ySr2CN04diyboQVUthkAc07nIhevC1G1WfFE
U0DaX7K9E1MTbXkHpODmmnrp741oTCEHWyp6H4sDbE/XXFmjAEKCzywBdG+ISbFicVaDQqtK4bf0
qOXQXMD7Z2JqMz/9kaLMU8Gcm9qyahY5gdH1PUtnU9tk+lUQW5I8SYuCiav6iLWC0SWfQh9OdYdy
Uyha2MqoAJhFOyeyl2xDpnyDJKaPnGZ2u/UohQsG/SoPotX9Z98JJPBtprweqTCexaJEtiQcwL5y
+AUxmETUxZSkp+AKAzwcfzo1rZYNLpFoGIxzLldHSLGfSXvURI4eZvLKUnF5NTHJ+vUmjAY44XUU
f0CL5IAnFPDOXnIv9jNLOcug63HwLSpKBISzWtat3dI52vFErItJUZpJZDI3Y6QpYu7zfbk5D/V1
NcUbaTFTbtcYmnq+QHUpj3zsyYppkotpmK77VKICYgKJ4BzPYp/XU2l99zJwbKwqVTMO8YlDcas+
hd2KysIHBu5osCkHTQ1ojDSXfdKY36sZhhGsg5lWiVSrRQhZ3N5uvrIH1L4fToMjDqqUOSevNbuG
bLyvq6ddZtCI+Xo2o0yryqsbruOAJKfLdVFfTrCLB5vVdOWjnXt+yJ1aGYHhw/zJ4NF8hiUq0jGm
aqq5QyeGD6pkLuI5lTgtJ14LcBXGWdvKwmMxQcHMvyu1CImoa7MdbOFDfkFTFElP6KS/RsdfIw0v
eY0lgPt11jt/LKiV8kpPILru8+wghZhxgASPX/faSAvokXVtxRY3Dt1Oc3QK9CtiKuVCQ538Ryyt
GQ1IHNcb2uBsLzGWLKWg1LJVqyGOXu/nSSXhU3AyJzghhghq5P+gdx4M08f63CWDkLJRorn/9MqM
5e2utnUASp0PzoacqQvshWnq6xftVCD+ucE/X6MU7mgwJMSsz6NPI/IbeLzuFr4cz0ZzqQjSG454
w1pjqkRgqyjsNvKR9KDxm0FhZcLvyI3SE8Dt08i6l+5vBr0UV85pM+Z74TN68+kF8buD5Pw2gSle
SJ/TBo/6j5na97KCXkQccZz7U8tCuN4DOJYe3jzbjzyxRAsxf8uosc6y2RozPo/nUNaToQKpShpb
iHTtiPyauAylOYRCLCWlop3wJ4pIYl/H69hXNyrHtd5xmRj7LR4lZ+ayF1nwMM8C4+F2Y3vuNpSF
BDXZTsj/Q+BjJ+CHJ1isIj2s4WGUVjh2AoYb3VULuS73CzC2PyGUoWzVFwE76YOf5QzKwn7NvU84
n23heK808H+CtdHoxci9cyOvp6XoTHTJtVMtJFs14k9P6atHxRGzEHCNmGPCKXRGzejvfA5bEa6a
FSYqFF553QQgiFlqz+5SD0MZd52gT8fscM+ZqMs2wDQNrD6nBB5zS6HbG/T7ttCtTWO2vcyUfWNd
ZA4TO635ng6bnj9f6RceCkn4wxXXEhqLeYLG2jhN6hxR/9+IhfMfUZXc6e/SMWxZR8BgSEBWFCt8
a+b/wMnDqeNsNC+zvJYgbOUNkQr68LWXmr6rVxtcQgId9SO4YF2+IA4lrLzcrQm2xj3bDToEcBlA
QdamfD7UEGGbOgGQI9SOshPbTYA+tyo1PjrCnhXtzUWdSzm4UXoiDdMX+dTXz1QljbL7IDqRMYCe
Y1zA8xWoa55C1xOQNNXFxVACnD5jv8xb0xzpVb3gOS/S2hUqziTuOEmckrke5ZBs+uCsbY6swarY
zGY4U+SV0RCShAgmpTdnvenzbwYLGhliMDA1LmtrLufY+MUn76y13eNE9MnGQn7u24dtF8S1FWHh
eS9Q30s0VED9rHhfJF+nqOQvnSyotklkJOpNKj4oX/6wTDAd6l5v7v/5wXyEuF5eNFGWgUyP5wNk
KC1DZLPy/0eSQDfQSAkKtuvXHnmLBBIo6x2BzfbSrqiCxBgLG+nYC6IiFdaRKVocHqbSJoaxxv0X
yNodp1n+bxfZCbgddVfIHMC6KnXab9JzQjhXbQFFL1PDTGl+YTuTXhIpDeOc29HA90GtE0bWMLX6
hZ5j/Fh++3pMbv//17+1Dr0JICTjL/O1nKbGO4kqXynX+bHXXZYPCHgB20M/K6XaFSByxs4Xq4kX
LFE4fmT9s5uGChTqfnt2qrWnEPT7fw0K5HT7JFT4lVB/d/6qKJ3YXoa4op/zOPygCqxi09FazXFh
VJCdPzNipXqEDOYu2Awk3ed4Nn6rZrk9O79OgRHklHINTKVHfBQsOnT32zpRvCHKGSsCHNcYUhZu
hnKAAE+ZiklWaZaXxBgQbd6DGTkLKuAv6a05PlU6d0zESNaj4nzzhT5EXolXiraCWZ5O4BxP+d91
6l2o1alkrnZA/1n7aABBKbOGNIsm7mFwqtq+C1t8WamTvc4sfCjb06uHl5Ji3HqGIUG6y4Rgpsq+
AjmchNl4GClzJlIWo7PA+TjAo/EHgz0InvzQkYFcxWlF9YYPuirXZYaUQ2TU6SpveLfQe93g5dUI
yiyX/rJ3gmtKbypEJ0Qppo0Mnmc7mwWG2KVUPs4rrW3UVzVTuCjo7vaz4wcpK+ogkFay1FjQLabN
Sb0VqRC/SeCuLaAFnEJWEH6neUTKUTplG/Sdv/GR+849GaLdIZoynjbt7AONzhxboJbMeR5jNNUj
mfObYqZAprk3s8H8UDdmubhsos8XM1QSRFammw+76YMLqn7GniXzE+HC/brZL1x4tNiakftKFeem
y/15R4ld7qgiR5wLk/hawsWeN3jrfYsq6RxFIh+jBPunPUO5bakKMDGAlYPS8G3VLUW8jrNlyjNQ
mtOMzNcjL1riQQExVk0kBG3SLvdttt40SDWWzuhtBmsB6p3CJ42q2ZX385zUgtKkzyVWaM3xlfeK
GM5KLMfPZI9OaK5h3HHTEShhkZnBMEi/AM1zTWxemVPmlLlldjUL1TrPXS8ibz/aK2PKeKkhx/WU
Yd1jWFE2JdZj1mzfAkSVz2tcy9onxriNjjCy39OUyZ+5yvMIMm2jv8hSnHhTU5rnoY/q2sjNFfPv
jI+grXfN1ZVSV9BIPjDUIGXulEgLi1pNPU8LU0OmZElUtqaxXEknrQPn4//v7xchld7VeSyvNw5y
K4tcM9M19Itmf0II6SUcGWKKlbaalxsq6aXDs7ZreCjTmg9q8zfg7hi3jnbdTVtqZj6Dn7VvnI6g
r8p8UpQUXvGUpWnz8/wtWNPWrohllcZ4BeeLwkGPH8f0hGmkYlBd2riuwt9Ltuum/suzR8U00Fi5
MdQilxHmb8Uo1kwmOL6QJLdR4XKg7tbJpZJokx1ylbXBOMJ0o6gl2eRt4E1nIP4DFX3UbkQiJFPd
oKQdTe6HX4xEeWzbDX5GAziDXOQtb6AZ6i7IoD85rSCDYxHcDFVFk4ltQfhx81GK1KtTQCHeYKqI
xo/hjMsa4D6TS/r8sSvi3P+qEx1sOvhHwbTejXeeJ0IbjPj2OCgCbknZBbIhuQh8TF8SFAtN3m3d
TdI0r7P+23K8dV0PDPQfgCTn8RNhepW36e1KsE19lClfdkbLJUNpdfNmwjpTgydsUTLIzO/6aGa2
YGt91RZFWVPzejOb8dgrOUty2Jnl4jButIWECTLHN/dSOjkQzicPWNpRx16vI/LkiTSb0bvpyiY3
g1J4TW20yoi9bxJFPqJ1s23KHI2wIjduPUoAlR23iYKA+xZyiirNK1x0tJcUrPaRLpCRqyXv2bCJ
8ThVW2U55NAgBOYJvvnu11AcE9rjj0xsbDlgx9/J5r8qAyyBMwDPagN8kM7p9VSSQ4nDPubT6HeE
3Pk9e7Zfg9EJG4byCKE74VnZXYrgiP6qGk1b6hIWYliWzgHN/Tdo9ia65fuCzDEuz2IiZo1rbuso
7D8hUoYnOJURyiZ5SCj4IqX+4W7boLI8zaahs/VsnsXa9MKaCiEfwg85nr2cV/3H62pL5ojpOFxq
3PUtUEHSMOnBFUrLPWWN1Hf2rp8JJb3yRkRUGmi6ZMmWmMzKn2D1iamiHf5I9ryTjKkpfHNMKyfI
33K3t3WJ8/opwMIccB2IpgDbRv+pPR4rBiGUvXD3ACZO+SPplnGlTwAuGXrK8el6I5hAZCjAfvA0
jXE+3kBvUzpN3q5S77k6NlG9fJflTW+XCAOCpUNTnwFHcrAYhGfncbV7LILuVPJZH3+cDSQf63FT
PY95CeQ2IAEXBwRMnC/n4qknsXUoS+QvSwwbSFFbxJEDJorxlzwbnBzWVTDfPhTiPyZXLuLQpPt5
pHq7U3v6dwpYdtiwr83tOUqhAmlf9VAaYG+Dhws6m2yRrBKWVX2nq4kQHqhLcalL6pfcTOqrcpCn
RjJVcFFIHw8Naft6ISbZCtRIbzOSaBz/m9013gub2NkMl9F2E+6j15agsekkyAD9VVUCNGPut8NH
QNS/LahnaHrT4b9qoEgnRzKmJ0fOMnawCZ1xk0F04RRZxzGODyYdHV4NJuhLToHhMNBQ/cLPEp0r
apN5MQulEs9KSLW3S0t2WDfH6dWVOByG1Ut1Lr27xRmR2YUh5AERugg1nox9g2DfubAMH2tBk5Av
RmirjYMyWsA/Y86UezbROF7eeGX16e19/RT3eJ6XEjZWpEFfop0ykNlOp3Wohvo48SIx7tAaLOD3
Y0nIvOUXvOHHkMEBrMsyHFMiJkJwEZmGpQtmAMvlJuD78mQK0owhSqM4jkHwvKMRPIiBWyDl0jTo
Tto8/nidgJGBqLoC9a7ZCoBxBkqHadeLS7dzaRSIqEXiZHQ08AurQkEeQ8Kvg3L6loOwZtNvxITi
LKhkM6covK8O7CHYdXXKA/5Wzas3z1AMVS0GXFrzgpJTQTYCB+ymO1QSBv91qIhS3u8IM9YY+wGC
uRjbmTeidbtP0w6rAsQh8j9JJhAHZ//ISmVkdVbGt9YXGnRUeNFClD6hJsJGm0KZ/W6pBXAtDsw7
aaPb/v0vdpQOPmy2EC4R4EpTt7RlIdbDexMQ8ttJMRIGP2FJSnVwuoO7EdO0tpmlIueZ93yyYZPw
CsfR9lmX57kLNc4vvawYO2TxhHAKmUrCtIhze6PC2Cr5kHzMu+z/bkPRsszS46P6BRUWsKPWu9FC
JZGw1XMu06NPzQno4j4uL8WJTnNq5avA30/L5JjUsZr9Sh+KCUxObPJdItenzXo01tV5aY1wb6Pg
SXDnL+oXHH6EphegrwUrlE9PEOpEC7ZtZcdOBKHOiSMt0RFdjzDEaPiXTVWkprf+5vXI17jdfpBL
mdKCHcvKilvZKtdSo0HYHEy+c+WuaX/46MYjCdpeeOB583XvgiIuKmGoyy3uE1a+4G3xNupx9Yco
/7cNZrdxsaCpuS+g1kJiH7p/JniKBWiw8LEdOEKj7DFnSYFFBECeTSSesbXE/aChRzU3G2Ux5hda
VR5PWy2NpggO0qcb3DtBMJI2VDKOuiP+R3/2nWXd3t+gQ6mCnRig+tS4o+iA94tlvkl1304jgzmb
C8SJF9dwvXrM/rcnK7idnvt/GCHze7plN/f+mqtSmcc/oza+s7mIrIAXUC9S8PaUogQswzFHzKfZ
l8Z8xYu7vo25ymkPPZ8n02byZ+7mqZHhtEQW8qXaDxeUOhIvhkJo9BkpNXBh1D4EwPiJGt/IOI+W
A87O8S/ucGPIFtM5JJASQM6U8V3i/f1MjXqbf6W9leVyCgHghk4k27aZdlEk5wwEcpb2YcgCLO2Z
YkJIriWWH0tCjFHqLS/x1r0yeZJTGMiswVsB1/pOjsVXBu4au5h4qF3qAi4699z/tUS0tBfUab9H
m4DJwFuFV0bnjM7eBkF9CyizI6EbRrbWKae0xvk8CuL1o/XoDIX0Knw80UMMKPU/TGBkmi7pJrFl
ovQmM2rkCnob5dJ99MIgXhVY7jh7bt5oXg/R4eOwbs1+UEjiWq3ywxIYEvuXwsctnF5iOG7GymTW
juYpjwF5QqB9YpNZCD/2dcmUuMa2nxMYoN8PyhPAF2Uwi6moyey0iouNtHANepAOEjcX0PPiSJaO
6ns2fPhqyPNN3p09tKlTZ6Lke3TFld6wStife+pEUKculyVBGllcMw+ZWORMKa4kEvdtH9cJp3CX
yc0kZxpvoVuDj+DkMxb60qCS5fgrgkCNZeh/sMwwuAimn7i5xx/xFvuaamnIzTK8LkfYJUQympT+
atURrMPqEA3baj/7cmN96HGb0yXlcM7GeMpCTlzKROS43A7mZVgLwnAR9vpqfvtLWU/J1RDr+s90
ODI8vLn2Vj78dLGxZ/kas6yCV85J23bCC62kwGloZlrmGLi9eyQ36U5gSv1wWdql1YGuVsg/XTX5
6OUwPjtZoW8Ak2MuAfXJo/1/XjylA9CFJRzprEWkfe7P6KGQpnzOInh0jh74Ylagk/FWYTg77lyF
iDvTd2AO5xtWgI39Gs+KcJ0QwKWSsA089zse1VGeXx3i+blXgrOBdsZdCOcU4GBRVuxUXJdPSI4b
nFdbsjIdg4lQpxEDW87UWFIF6RBDSX9usS28FMdeXCrtSJtAxG9AtN7E7pP2I3cRnXRn0Ozsc9mx
qSw12cmsNRvWLf+H2gaby9GKTkMtO3LvRv5yD969MCj+TUY1ARFJtfOrFO8maS9b/2xgOsdKuSiv
zLV+vdTo/rW0qYD38CLQ07/2SSy+otA3nyAJFOIDPg8ZZPOGlZikr54ze2HqtHHLL2JA8nALNEXn
m3deSoB03zeEGiDo8JL6jAK/2RxUQDSakBGOQgYYghrUnqc5ScWVLyynLLc1C7hY58Jd3MjZXW0w
fzdm06394lPWiq45UjvYRAcRcmBuHH/xlI+EEn811Ej+AJnL1FQpTMb6pjbfqXBvm1GvrrTgFHft
jCbN8rz5g9DKjKCzmCHOxTkP33mn1fDan+eOEJMnPHb25poKpEmfwbb8HbJX563wkrjgDuqliC9j
nCyaPfC3QBQ4G5fyLjdEH4B2F401uMV7L7r524ZzbCt5Z0OT4Ca9sjj284XLhI7DvEw+IdWFxzFD
BUZd6OZ0hDLvdR78j0oSBJoI1jKoUyk3FnmOu10IdYrcyHtYj+mnQnhtBze2cp4sxeEZJtX6ZMv3
amLW+D5i4eFKkcf2vY88jEg95ctTKZn57XkhXhreAiJyINt8duTsz9MhMtWDwaf1bi1bZQ/P5sEC
nqPmSGu5M6rDZUJjcvQ+VNk+t8XqMKo1BPG7jEQyAa1yKLCdMpWmZjqfZnzbb1WaQyak0hh3hCw3
bqRlzLlJas7lx3mTOSJ5k7UoToiVLXo0MhQGoIa0c7foXCAOV6GBnhGYA18zlWGZ6jv9rEVfU5JT
oW58d2BopFlnBrghdbYn00orBvXVK5G7PzFpH4mGNvK7ayXaHxIdr6PzIN/yo3TRLIYMFioJnmGa
aJtVwGK9Zs/PuNU0o2iaGxj3t9lKucXOsUnfffACvGDrp3UCBw9d9Rd2FobgyJeWLriSbWW4is6M
oPSguGGrvM/gz0REfmUaXDeWikv6YGrDYx0oLS8qd/dJShQCMQebDBWfQv0i9Q0tA4AB20nCTwDI
UtAPHP66KcAlpCC7+hj+JAhkR4g549pStqrW/Cq3ykCvL82xl8xJrmxMk2Fgn8ON9RD56izjnYJg
R3S0JRK43GJ3twLVihyblTqBy+0BEC54HXQobl3ut0Q7w/4fIb1DZ2NsG5L7MZOVWP4IzJAr6ZhE
lbF8Rdr5Ps/SIpbhixP4uZAA2esfdIcAERTWs1ay+lJqAqBJSkTKKe5zaSGIqOT2dbLDt/f3ifj0
NlwNIyWZ4RaHFRFi3+Kx+2bZ5FmleaWAS+xU4eJAC6MUhfBK6L9iSnuuii3l06WZ1ToE4CVl4b77
QTp2wBWedmk2NFxyvH0bkil7Oq2CYKXXLxxqlyqxcAEtNQf88nBOootKWX/ReVF4UaCJQ/XnVJq/
u1NC8x/TeLjlNVVfI/pckDOlBRq0G2Uo5UcgxXkLrm/ZP8EdYOFXIeT7LCmtqtRxNqOeYq/XfEy+
kPBoqobH0yyYM5+7WO1+gdNIixdgk9SxJ8Ehyy+ZwiVugsstaZWprD6d5L9cO26mUXzU5R1CoZQY
xhvkSF/gvpwp1PrjMvpKmuZwSkAWp2kDv9fSEPlcZNeFfi/yio3nuoSK5W4LS1i0W9CWMB2sUbUM
8QT6OL9Wc6H5SHHfyEjjKbFU//BH0xgdlVn5Lju8l+UdOZ5CciEPRfhVuntbmlmk/5d5wNkuF4t7
RKcp6TVGpcQJ7jqzG7jFO5ol+F0006fSp7Sy/mj9zsQtetf5wbNf9nYzFBtqa3v3A/B8E3QLjW3t
u+VCRuOhPXUaTwbzAmtz0gVRFKVxxpiclspNcRIVVEXL4wKEX9GltejrHQgzc45RtNdZ11v+KfMY
5JJdJ3P5RZj5eKxOmkMbwRYMYlzb/OVgguwnzHGqUJZKFxxZ3/QjXlBTspi3br0HzryoouQ9ROur
8pHEOGC4g97WIM9Dj5/sk0/Bemh95s5K9Td/l7k6Z5D02C55VBfIW1IftNqKyNwZzzta8saZB2W7
IVjH8OQse+TzCIUTodnUyRAHdMN72UnZIjATe17jr3lPyW1KKZLoYgCsPR6Lrse9/HP1M5h/D4l5
k7w42WrdeYsSIsWHC/aQqibOCVRwW794bBDIYFNDoVtE6heX/UtOKZ9kSEl/yqj2E0S/3Kjtn+5t
+nWvVIyTM0dTp4SQaXGorEdKkj0cEyvpldz+hqEDCVUNARf200xnfR4kJjBFTmTnl7Yqm+xMXtsm
9oeocNTKMJbYuW9OW3k+IkqFrCbcW6Hy9kiFFWYdHkE4hUKG/o8z4d9OdNvjfw1t/KJoVEWhIJqE
jgsygvj5rO84LHCG1KoMimgPc/GzVE9jqtgGr72CmWGImqR8JmylGitbRW+jVqy9FnGzUwofTpj+
eL4LiNNiwAw+OrYDbL144EPdswNxIE9y20etiuJm+wpOmXZRWXs/d8y7CGAoI/1Gx9+DcOOD8K26
xmocxFjm0Zsvo5oW3CRVt6o8dRE1SnF6I1QbWAPh0NLm/NLJgpB9JlqUixEZyiIj1qK/XjMQaeC+
mMejG3t68mBzGGVY6AvAJI1bmxGDVGJr1wpAu59qMRlZ2dYZGXFzHS9FLbCKJMq4vZGxTT0nWXFd
1VDu3ROW5sDBWC+F2CfPGeu9I04v5IpSJuBjp3B/KzgKyR6lL7yD+zrjgp/miySZ89mkyJNIFbHx
KbnKI+4uMqHFi8soZmQGblx0D3xDXnbdr7pPiSZ3SVgj+guqXDimtPg+glKyQNVlVIcmQUYxAisn
5t2aPyMW15CLYHXcLh3O7zzWob/qdyIF0U77f047+Dd043QNGlaJh86aYL4XtUwq1XcXhwDUI4Tk
J/HjtPOxx4j+Jsppa6mOiwAk2PHEEjQPZt4QbxgXUJ0sFf3r9imfgTf0+hr9gg+wqQYyBjp0Taep
+Irc2VgoAOyhZT+dRhadzpLWtq359Sj5/45vp0h5c2olKE4S0SJClFSNVPIsQsRYatp4ihj23zue
svw/VGhTqw3jc9mo4RYDikv6+gVRLfNT3ZmTM1ROohEbdOFhavhn5rFZBU/RFGw2C5v3gxLv7wOM
bYX7GAVTpuBqRJEMza5KAdQLD7MojUsesIR3T4tGCMVLJpP03VVtgn8Mn3Lur/7sz72ZdvsyPnDI
Oar4qKcD3yF/ASFuWzCUou8tvv9qdquBUNQz4nyrQ+MuJ5Z+Ym3zQ5gvVct3R/W/TgHj+KRPJ0ss
4DQH/GyiOvis0llfmv+lyL4JWD4ajBt78rKl6eN2Aa+qDRBYBY8j3Oz8WoxcJT8Ed8f6VzT2B7Xx
EBDE73VL1JacuGndsnD/i1GRX00X0wcW/ew0s+77gOGL55gp/NhVykQephqWXlNgzjTMZg3aadQK
fa4G7yQTX9Ms+zf9gOHXXdgmJGLkL9Hqaz0MOf5DQXUr8aLEsD5ukVO6Y+mFlcbnQ9AB8eVT0RFT
tvhRnTQWmnF8Ut1bombtNWZVtGd8eq6B66IMc2ngsiGXaJreOaTULPAVqUu1j3FBiQ6ix92oRnQL
pCX/+xm0Zwqk8Zy/NyJ7aKYCDRQBkTiPzbfbA2FhDUVurmxpp8dO8khJM2UYBhfZnRtTdheBU9I4
Czr1E+pNijYqjNThoNcm2+xRuvwQftoJ5dGyTHB8XrQvvcGsqH4M7y48dN6QQfehmFibNyk+ZkQV
jCYsyFzicnB+L1mXi5IXGndd3VT5O/Ud+cY94nvUK2Ltg64r9MV2YjuwhHRQ0ZUr5KO7y7IU1w3v
vKx7vdrdRDqjD8aKzpo5togjBI33zx+LT0zA4W+aQhyEOBn6U8amwCZUGSG2eFgN02leANKHSPVx
U4pGfj+iagjcLDRa59A9hYZB640SDk3/QZCzWxlnJaylUUl4qUizFTCCrlkWDcdREZYZ+H/HWR35
P5dIHZw1ihrXEj9aU6mHhvIUtVcNlkkVXFvpWir5/GF0lftU798RfT07OlwJJIcJ1WxRvbRaekAk
p0RvJ7u/U/xpRBl0G8BgVn6b6xM+ZA4ziOOg6Xqy7e77JMguIzs4rUUM/BNwSGIPF38OiECRE/KM
Hgns9DeHRtXIVUvfWmkRgkHCNUpGlJXz/BwYsznV+zpajLZOf1wXWotlqxfv/UmLUqLG4ni0UUSL
IRGYxSDUNhGdDLKojuEpxVHCQboC0auzwvzhpyjjGsLklWq0fh6YzEW0Ph7ph+Td3dB54OOA2mn6
tpbrqEephFeXSzYPW9AThkwP9rUn1ZJWG+PL0scuLW8gmhWpdSyk2XhVWYYj5UV712iqhpb+KIuX
TaqJUK5OXg0yLOSDMMRSsDywSNpnRPb9ql1XJ+3lFrKQswLtpwyU4KGNwjGCKNO6Nq3w/pHTxfxQ
awUycJx0XauxJgv7NYF2VS8gB7jW87749uyIZdviZnIgvMTfTkPjzzGcSuKBizRQupGEZ6TzAhYL
QVPZm91zlGkHW514VaqJvp7vlaFgYuDOfcwAf+DIewDtSw1KUIZxhG006Nzj73h/awdRZtXiq1ug
HVDp0CblfOmoarPwiTrSxF6xwJpma87wXm2DAzx6GvZjGZ04pv+JColVfz34803DVjZ0w+Pgmyap
IKk191svimlx3wXdZXCDyxxdfk/xz8ojoIE6C7gbPDT7EvoVCeZE8EyShpr7SPqTSt34T93EvPS7
z/0YXi8Lyl2toGY6b6zVNQG86UrQ4ZhXvPV009Xy7opO3IlJscNSQ011pop5dR22/4E0eEpGzGA+
e0778PjJB6wrcVyaGrety4Qjn+x4QufaCKB1IC51v+0LC3nl2QGqSHXwN4rd8q1K4ZW/wQEwNzup
d8/fMndcQcR5//h4uA+x7AwlcqvyLST3NAz5dSnhZXFOh4a6tKsfBcZqoIc8COm8YTLvlu7kVAAv
fOabh99wAjxIGo7BytLlXRQzzH7bJEfplHNld2+uwFGtp/P7xbqT0NoSE4lKjhuKldOn8atLCGhU
GGxWrHp0NMRWgVEEd3edvXYHYvxSio+4zDkWO4hmVy0/xNlJPMWcUdoU/r5AzneNlvUoV080B+I7
tsK1CM2CE6cLheBKrU7Q4bnyK4VAM+W+bwZXgK6Oyu/8OlKOlkN4lF2Xy6XFdyvIMx1ZtzXgKJuq
I7GXHhYj4PELkgdVPTF50qC/H6xCH0yTRLxsJAvAWSliwsYt2ISn27qbMb0fbtCgn1vYSjj/LiVC
WK/fN6eoSnvsyw1YuTiv3eWs17au2w0Jj59sAbbFce3xbFkl2Jfz0CVmqqgZBVzfmvee1V68Svb+
88Uj/IyycD64Wotq6M0nb3q8+M84oBJFLUIpClFeQx5sBr//h7zKjtPJQEg+bf3lgRAQx28vAwp5
Ohb7KrfuuIyF8JZG0LVaRF4Ca42IBlhAPZXofIve5H3iQFzWELBY7wOsBc3uyBtoyA+uBEzV5o0Z
DfSmhTNGPSu32os4A1lXmfkblN89uR62u6vfk7GK5eF+o6+Z0C2D3g/M0PZfV0018O/o5wdoGXrF
J5AE29dqgLMBmp8yCd50kKdxHkEseSy7fe0+mzo4uBe69vhVuDwxmmrN7kN/kxdgy0lM5ZhQd8Lv
pKnmktcWiYLi9Qmzyacts5okB0C0L0Y8rmumg5zxiDKfChu+VAlnDpdCCbTwoQEusBnsaec2jiTh
x/VZrF6SRo6AYhi2Q38kmOOT8iFfD5b2oJ3puKEjux07ET15iSdsibsU5KVYBqF3aL4Cl2pt+QFI
RWCJdwD39zlz1Tqeftnh0A7eefmiMwv1si4YdFXNjecfpDKq2/6H57krPU1gEm/aH/Y413noUl5J
p6bP8eEm4wlHy0sXct20a17Ktbgc0xpfxperRAvY9+95bj8BY+r1XYQ0OLpA4vYITtkMYyDIO1QP
P5v5IhMgClzUtlvH1JpgqYr+gwLje3I7ezLW+u4Lq8zocdFzh8aA3D3FACSXkf1YIWKAZWne5i22
ds7p8YMW1QU21QtKIir1yAvwkM721gvtvClJnUiOBOEsyPqp/SN+0InFttsReYlqys4M9pC0/erd
ndtayGc25TpDBGji7fKde0hwaThUuJxksEfRmNjxqWKnkYahbJmokxcWv5wmNuCT2BjtSNhnusjC
7lyorYYYxqMPxOc9BgGbatFg2K/7GNr2T9pVLGBVtCCuY0Lwg+zlAGW8kK+3oP6FYx+q5J/VXLhC
1jEj7NjxK/tgK9YSifGR11rwNTn2i+gjd86OPpzt87mcpBfAFJNS8q29WYgs/idG9n4YgI0DWSSV
HLu3Uhr7ls6l+OwoWJ8qC5yL1RMtx0Krn/dkOzDqF0M/R6/kHKsuGQV4VFUeDZSSNj1/aLYf70Dz
SHYoiC+izkXgTYffO4/pwjm9vJWQAAZ/ZUmd5aBM00G6I3o7SZJNSgzdwCf3tQwLh7ntywCxc3qr
lhf+k+gQfEfkTKFs3idirjHhhCBli3+QRlq54U2NhpEzh1gOFTvL3XYa2knAqJV262O6ZlyjNtOk
hTZ+0sy4gMyUE7otSekN/alugCHsnZ5sgXH+i7EQaMzRfPVqM0t2sUmIEaw2TbaP92aAHdR+YFMM
r/7oE5fSsLg2S+QbgzIFmHDFRHussLWeOtBnt/77F/NOtPzbOIVeeQoTlx0J6aYq9l7fFdT8TbyU
4zKGEWa8CI5Kc7sijkQXeAx6Ib54jnznfvuHXUxYT9GQXPnPOJ/OxxUcHrLgDTRKzhNjnO1huSzQ
IhTQhvIMNqBYsEIZ3tYQH7pD9HW2Zko85OOV1uAKu+wLjEkQFMpC490/fcXDvFgoondJvsiECab4
26DS7IHk5L/7C7iSYFMQEVOCAlmYFNr6wqFO1NoOxnnQDprXrKz1DT9CMR+dQEhmqX5Z86e+RhJO
0LzdH0F+JSrOMH6gQhtaaMulvu4xR18QQrOLeBJvsXeL2PSG3Y+SYplH2FnwmcWkwp/tCw7x6pqi
ldJQVcjK/sc1qiK9J7s1VchrPkNLdvQDUiO/sPpNdam8STH8vISx9x7mZwPoMW0IfzqPmp7YXMxh
+1In/I3D2GHHASgCAW9Ecu+CtlL9161NAuy/cwrda4B91JygVOAPmZJENNYp/qUznzfPclcfSEDH
WksndaAgjdEdnk+hXsEzBvER1f8tcSWm61Jya3Egp20b/FG1tWDG2IlcxY3wSjeC5z6hBRe2PWi/
ssVu/fCkGfR0fcfET2RY1cJlUn5Sy3fhATmnH2Yc0v0UWXfc95c+xk2KZST2fBtnGHxC+6vFh5i5
cZLYtedNh31qdUpkSGzjnJDwjb/pmMM9fPfSz+niXoroOol4nGvouAGypOQe/Z6lX9gI5Q9FA5JX
jXUcT/ThpQsT3Rhra3vxXzS7Qy0kfgUEJDB2sd8b7CfCwewl/9sbVmtcq4A9M7cmFDknWyIUm+iO
FYpjAQiYEavZekO/HwsptqaG80lwGfLFwC8FiLDHQTj8Mh2uYw3SeZ2YQyh+UtBfepk0aDscsL51
9GChmRcaQGLBWanNfcsrMxXo0+8rj0GejOMG5UF6K82FO9wwwo++kImkgfd+SUc0ziCniQLXrU6u
NtPKV4rEBXYbs4Nl+xb6pBGPR286h6IZu3ccnM3WBZSyjiauDW5ibFFAZ8ZLVjb22jY+mbcrjrvO
BGcF75yGWVVScuL1evwXgV+Uc5cF9bPeD6OxIPaLDDzEMsfNs86/6ayV/PRVDZY3qWLQbMtv/Fyz
EEiM6YKx9X1vvILy2jMp2dqYo5Csg383gVfwLPXE+bauQxfu1MmpDxmSMqKGvzSWHizN9HCMY3Sc
0j2KnyrAghEaz8/233Z5+mekB/db7qId3mrDImNup+vu9XLOtQDBjucqXUysCCK4si8RDSVCl40X
9HcCZD0jPcI4LsDU/ICfrknbsLFKEC2vgcjhPNEL7tKVtN0p4rl/Vxm9bphvic73lv9rIbQBJrTz
i5ZbYFmzlanvTQx1DpFh7qnyS1DhV97KcqNP0FBwWjEcej43deP4rYRSnFjDxgTI+T0cotAZT1lp
fZywkUxoGCkhdnb/ROIFl8E+iyqd7WH3UlH6WKOUPHq23Bxtexdu1MDzBUS1zBgZgpJalndcjGmZ
EbReXRQAKHES+v0zvA2cL40GeMRD8H+bv9RovEH6kuzbQVOkbvddU5WCp+Tjh7d3kxLpWDgSUmCX
OrYQVdDWwx9dMDqUl48nDdHk7x+Um2i9/e2kX66f9TKIIh+ckRVrJXGWNA4LS1T/eS39tZe61pBf
hjISIM/KY4X8KQ6swyrP+2kh72i9JJkJv1MFbzUSCK5z1arin5L2TB3pnlZcLa+QTXwt/wBsJloi
vIhz4oMcVNOcQqCLTUn8SWNDqtKT67ZMFYL/MxExerNQ3CcyH/9QtvBdomIhfFUN8S4rKBGl5t9X
PvAGW33+OStwp47DhKeq1XpwlSPDMR4TTExDMsxMEJSm7sPb6DU9R6qsFKs20dkhzyB0HHiiPGKD
uNKBLm2eZSXZsSeay78AwtQPkSK6nvrlwvjNDu+Zu6nqcTY7+vTX3HFRoes0ERKUB4U06rSkxuXK
rn03mZhabErgh4JGY+B+kuIIAxvi/Mkxmsm+i01rXcNgBzs8+d5zQmarE0VqnZMyLqNwPZqlMC05
nSK0KJG8RKc0gv080goTkOwMBqMimKXGCegO2JBIh0+r8nADhW5gZflMxlJbNm948DH7znmpwusd
69trNGrhvjtE7y0drRieOErHvGNNZ/WqL6pILd08J4oRfldSF3gDkUAN1DCkQg9jvkhhiy98ukc6
xt2KLhkaZz5btZorEDZSkBHxv86CPkO8XFkMIuvVFTWA0tYkzbZUOLMdBQzignqzCxJmazd/QsGh
GIo/I1r2XwlL2jmNPxflAlgUboxv/VH3bwFyI8FJxp0kXueR20rcUTfh8acU1fe4CkG4Et/v1MXF
AwuxAkycI2qXeFbsPkM0qYGYsjkVjywklF1aMgEfDqyzx+9BlAqb98shTtlQVnpyJ/q0YSOXV/2/
1gnEPHFoyT+xpUUCcEmhS0z1bC0KFKFzYFLcZuJaeG7r8uJk0wDnbCnD9aF5c9uaQhthMM2bZFyk
TwxsT5Zk7aaVPy1B3voyW/FaoTMznPVUG5x5UBuOK/9NrMZVF+AbRYxsxL4miy/oqMxTSWFfvUsd
Q5ijsOKLGXHpzqEhJGdpOnutjS2NcQld9vBHi7xb1aiYJwt1XEITGig2kwjK1F6mvdUhu0egWYiZ
5WLLEnsSHPAM6rfVC//okKPXg5iYK16s7u/+is/AdYKIGgOvr7H6rWMGf8Tdl/XLV2/iNi2rzy/D
a5fMmQq4fmv51jrLWLrsRcJchUCtGfmiyvMBVTpGfDExrIBEzNy88+cG4yf3/HL3OusOli0PN0Xt
P7vpSTPGLcpqNRIOvvsbGcwhjxlsMHjV45F2ogNHlCgtbfDSrQRH0l4DMIMgdd7i1gQi0KJh7iHh
Yy/FMmoY7Y+Bm84Ge9S+sFocAW92YI7E6PV8VOIg+QtJ32L7uNKmcyhN//ATUk/AEPkpA1PIL0UB
iEN/cDmdH6enlgm9CWRGmxSPEGkeN3YOPW1q6w5Y68U1vozCU3uM5PpA6AcQtZ6PVZlS5Y+GoF8l
hktxCEVBZSHUhmbvJUOPgfiSR6QwbRO2LYZEwEWcFY5MZyQB2itJzMZXMpKF0bpJ7+fBymDej/dj
zTmJ+xAJMFVue6vJUNgQ+4xvDFsdr6DPajxABc/KRRmeJ8FFhVePLZOoVRxNYNNNKnZ+Q8gv+FOc
q5dFIRYVxIbu45BTB0b7an1RddSGqAdlG3DUOvNYNNqCERhwf733JF250EEdjTLiHxna7c4IB/o8
OTobjKJNzR4oPgjAlQ2JK48WX6ko+RwiVK0oH4gj4bYo7OPGteCxtm375j3FV2XEwdDefYfg2rNC
lZ8G4psPcoujYLd3Kj54r88qR2xm33P+80lsoHKl1IjaueNMVNoOoZtPcFOvAkmBS2Z7wNMfvKX2
TDdGpKdv9K6b//7V9cEVc+iLbMfx4tNOIq/35gmLQpmDtoaTspcXRQcuV2dATRRGtulDcsFayMVl
kZVot48OhyaCaNelhKJIAElcjZaV8lI1I/cNbYcVfMd9Lotup28eEmW6Rv7hdbdEbeTtUswZVTWg
BVgV/wpqs6Dptzz+H0+E+iMXp8vDvCOyJgFqi/Riq1F7ISQfxaSStPHdo8WiDSdX/C0dHl2ldWdP
OodnvtaPNoGPBhFqyZgN+izbKaC2XlPCbS61aFkOOyzhvKou54Rkfe3icSsFDW9p8CSXpaRWZ7z5
XrT382f/b5Wcn6GcZiMYewQWDWi0pEbpebGx4VMRyzpA4EIFQW5dRADY4irAlIovsy/dw4Hfg10z
AdorhFrpFv8AOTCIlCQ68xKfRsY0UjjpZ7efkuAgqituzEvBnNseGYbEKMwmafvkYjhrvRUDeGrf
7bJqcx/nHD1egUp1XUe5kDMMEx5Bm9LiMMnNYlBWwA5gmLbrwjJ3xkO9xPYcc7DmHdQAOC2jo+3h
X32s6VQwMRF6IPIageI2bJ5qglvumaeN40D5azjqmvnIlQLRIiXdUrRbUZ7FJutL4fiVKDdDYWOP
oIP8GP1tICvp7bxikzmIbLp28wrC0JWHyleAOEzjGoneGDJEJW3Nr24xv35JOfOEkvFJFB2gW/bx
OJbasBkGFDbFu8lIW07u6yLkJvMn7F+tasvQKBALgl11Vfc00wh8hl7sXbkd2s6/SwMJY8Wpo5j/
lSdIOV7PGtFZUOM66Bgwqrm4QaKIPVCxl7YFlOxzeKk9JfdL84YEYVW5Y0kZOMWmxh086acidvdK
jHuv+bdIpEI2oCLJ/rdpP8Ow7kaGZuzypQ10bk+Gxx7UGVkYBtaFSXoEwmPlnzn/gBzsXQs1DnqE
jqVuk6AK4NUPJHMUjU1b33mwc5aUr/LPI569H7h9rsmZK+E0wcS4tU5vF+hBuXPiIUNsU7L7j3De
Ox/vsfVo/0UuRcZL+BJnO4d6oOyNlvHW9WWfg5cNJogxkpXBGvuMKh7A+UFp+lB7bh2NdKNzjIe/
eCx6dC6rcfTingq7oAYTYFRlT49OQuKSeBvWHtFB8ZMKmdTRIuNnMjzuN+cgs4jM1Qoz7HVKTcdy
FaXhb11M3iboE9wyKsAogz5ZixrltC6Mzq+aXM5b66Cq39z58dbsFRqC0gGLMeLR3ounUki9ye4/
MqQ2EZ/IohTrQ7pBDmX3XBOfMARcKUaYIb3qBLU2pW5d90iOlbPjj1d+0bEAyLGNs43DnVoJ2uSK
IjbnCfLMECIiaZMTgx7qWxg+r5M+iRKAROKBV8DoUC22gkeXwi7I9xpKmbY6dkT432/WJ3peNjeO
/2Az0KvJZjuPSLQNDG7V4fS9lHTV7rCgMy8d+xq02UFkdFUexBXAJIExrfOef9I6qn2nt0xtntPJ
qcQYGuVg+ctS0nrLWtjM7UgIVLto2mPxJmx8G6NTDtqWwopGLDfI6dQkLcTBBVhhr428yrixSqWt
yL4QFtQ6WVJskuNvjQ0kzxuW+OFpbwRHwhPTLcerhl7AobZjY4vOKTpgeb2ziy/b28gjtqZODWFR
PEmY1MLjK9Ou9Equ0VGR2ANKeCX50gVCL/FGWl07fhzUhhhzA2qhT+l9PwdOqM3tX+moUC7Bxj5h
bYC9YzzrhZZ4GaxPO2oab4YpYSCyxRvJnHehOqZ3WH8+ghnItDUe2WecOVDVx/H1ZNUPIHH1K+h8
FVKR2sbxEUXdEpGOJqCLZsT7pQkSZcCkrS4oTa2Xuilk5785b4B0AKa/AhdwmBfYN+mUzrPdC3lS
hrGSU5Gxy/U4HJEpAeelAUHsrZzoMZAUwUPEINvrtwEvsWOh9V5yRVYDe2gUeTC7zwSjjQHXDgpc
CHy4b5MV0VqEp152yQ63UmLOkSdXD/C9DladnI46Ad1gZcmiEdJp54KUIT1sMHIdHOvMYZS6dToX
pEYwlL+3qqXkpOPFJ1T5gDqvPoP/KbcXzY8rE9SB7v6GVrho6j3qJQA6gIRIhSby/qkxUiESEG66
fTzAIyuyAiZZuPTWRUbR/FoRi8gKW/mwO4W+AmRNaj9upIzVXGxtOWjomHmcGPYyjwhojroGQnlQ
5ZDHokGfKQmCOU1csGYGVaY6YLyxQmx7QiBrXr4aMsshY4SR806uK4eD8bi8ys0CtKp3Eche3QFh
j8BrXMYOnHpakXQq7gvd6HXWrN0NZjBwJBDpCC4cmS2mgEF2Qe+5troQsupJS7gk7xLnehIYyYU6
Lw8klNhcOLMS/FW/r43FI7+Cj5EtuU4d+YN/f1evSsk35V0IxXf234RwcRGYjGJR2gkQKpTYtu61
Zjzs09mgMgTvrauez2S6UQozdLe51B2/GekwRCsL5sP1Vf1UDOxRHCBQPyrY2l+1fJmBZPqETMjf
AODNZubUekGErcpJTDNma72eC0nlqNgMKOivmRRV600rT/iRRTAV+9f2aRGegVSQnPt4jD/3+fUB
wso+Yy38uk+ll2F5HMGI5wzPTfO9s8GU4CWUEWIu3wmftDSyGTU4jnNQnL7nlBEKVQVcgbiPHeOd
uKGfradD88zo24uvl+q64pUUxEY9kPGX4YUdvbt7dtQSfUaqdmyLm+V1CfBpEo2pJcD2QIpyRglb
+Ki6C+3kccnG23WrX1y1dYQsK9j9UNea0kjAR1i4JayIYfhp2kygSNfYQooU8a0tMU4WGZZnnPXu
wkSoHit7kBgC4d+ACopVpCXnGKp3zciQ74ddpYoBkHh8/4X4N7ePr3J3htoRYgVmCtvada+nKCUk
CGFgmYzxINGCrMqfGnkqMx/pRCTQiLYupLWtr/g0BCebKIskIDBAi1g5V8bQSaXwXnbpV80g4/nk
O4p80Q58+oZQk8oW6Lskl2Eas/D/uKFQ6TYMyXd4Yrv7rygIpFOPT9obG8fK4R/cy+Xe3IFBgtBq
zYa2fn9qzuz7jka9YfFEV74O5D1aYZTdDoh4dALaGWVl/CwlbldoR2vrtzqGiYpCgScfzYxDN0YE
wHKWBrorjplTL+Ahcs4ZrzS+wM02izkjwLkagDDBTOBSw0D8IoLw9oi5tf28lSKaTPnk6RwNx8Qb
Golkn9oAK1vr/DhijTZwz6SqFjbC33aYyyYTmhGbiA0ucZWMoTntmh/92wtXQVAYlAYf/8X0DXYZ
2H/oZ9CXmE6vpzOSYzXmWQigNzCX+UZ2UFtz+4Nb1dSrWl0tWz9KpUBuv398bzzHl9IJPRb4PoUu
1f3DN8+sxBRt8C+cpjNGOqdh8y6ydx/jKAMHQ5TzIkUNxP8rwcTZFWaqPfTVYQWEzL5/kzb0Vka3
1bfUz6rHoCh/FjgipyYQsL/XQcHHUWKDGRxv7Ki0HlA6q89js7PrgQPzYrVVM3WzciqqmuPJZcfy
HRabbaT4J3Z1g13N1EUxdR9pZ2WhP2lSH4KLbYMSzUvADxi0ouY2EFKffJEbEidAF0mzYBa9UZ/Z
fPM+jJ7/WQ4QSzhW2FmMxqzduAopY0F3Srcg+yVqtMOfUgVaShvBW3BSI8kTBeNW594k7vUCdtIa
W+7XnL3mLYJIAXmWx6Qi3uHGbtl2/jpBuJYmg8VK9ID3vu4rXy7vgoNy2KKpZD7E6/lq7YxHrza5
RGsbcHT7SOoWUhu0FZrV1+BNjFgoXSG9Qo4c69HVFEZkNOPOQyvJNh6sRQ+DtFsH9KZupkQi9i/E
g8Yi3143uPkORamv+qgEw89bf0C0esDbOqxsB3ZeT5ZkaAyMmqsKdkc32wPsB8/ZuOILAjn3Gzxr
UFEnwMuWAEjq3dI1YutVtvRWTFD2kK1dreC2Ni/kw4xAt0S9C9hi1AooH4JRJG7BPX4DLfhYPZC8
vc9HtgL9L7Ug+Amao0asYM68k6Ra6wFLFDQpR4J+JLPiCfbzLjJjnvpv0A8CvYeLJ1ZH0VtCFWEc
up8jeiSgmugZeRy+nbkeZZk0h4lmD4k2Be/iD5fgGuGaWJnMqJfhRqKs9QVQudh4Yz31oVhEnCGm
GDEpGqd3CHut8bDycpsi3kinxDfuNEr0mDw3GI3mGhvk3vV724/IA6ngSjt+ZgDYzMMZMtzblVju
SebZMb2PZ4uuCTkLDMOd1Y3E5twQwhYP+SiotdioqRAcz7r56p8WrsEasPlTqnaxnznlrKeSZ+Sv
2ijB9GThyY5XbyWT8Tr1d4cQ8mlRLEpW/5xjmwm4EGnKGHfMnrIv0Lw0XdfFOQR+G0TWbZHd8W9q
L+4BEXCq+KURs/FWPefhKHr3f/EIlhveXXn+q46Z2AAHAYnST63KreGKlzW8y6uOam7xF8V320H4
lYW0/ILJZtgDqqj4RvGOvqMj/laxv6lvMFAaS+rCcSksc08umX+Fce/e8fnXxnAQiHjveRcqOBo0
toJhlwq9s2maNsiU2WaCH2zSWzSrQjAVDQmdh8R55ZqUCPDVm5OXISN3LaSVcltp6C93ISUibFet
kFHubOBAw4dvaKK2MweNwz0qVGHAjdvkBolQFPKFof2mHFPirAPjOiuOjIg1fjpRsci+QF4vN/xF
BnGQfiFAVJUOuI4ps2rUXwe81erq8U4ovQ64pspp/3DViApgj6GgZ0K87d7WmN0NzHvUmyjrzUyD
c8S1bCpdB5+EAyIO1y4hRKXS5mSRT3yBFnl5pzcmgkRJJw5+bZnQI6w1vrWqZT3dwIjMBQpcNPht
vN0jvcmEIf+hJ+023eFzVhJP78Ry+3wAdKQYWyRMXfBdmBRmLbfg+0x9DJvEMgGexUFFRJdm6AA4
YR8qt3WsZCPOeqSrD/Qcv4Jts0OFwAYiQOHLPWuvcfSbPzUPxkJRZZGnjZEQ7VA6XLS+NrD65RFv
hVFB4QzRFfuOlL+hP1F71UH9IkD7tpbcvp+2aGt7k8lNAmUbKUZmndqvXzYTWxWRWfom3Ta+og1k
L9KW1aquWISEr0S0gxjPSgXeZmWGZE1CMjbM2lVXF31Te52Ddw8Yugxp7nL1jBLotMUvEy+cvRhw
81DASME+vYk9LDN/Qrz4vyzl+bmtMQqAFIZT7FoOzCNoeBMIAG8QqjNAy7bwS/IpyGys8rQpl+z6
I+rqtM9xZCKxFvlwyTwyvn3wL19Tl05UbpJNLKUNJT14AOmT5GuFPIkRetlAoaw0qKd0esA+lpJa
vaeIfz2Iw/7zlH5GfbDIpjt4R1IcyHrHD0NB0BNRW4+ilxm+RnOsxa9KbsczeFmQ3QFn9m8HYnWv
YiAi7x94jJfc35IxdH4uhxERdPKqKk8kDaKNxq+neLEPnT1A7G+FbqhCoaCY+MWGroDAu64P7pen
cJLVvlIKVSDXpjI9tfvEDWMGbjplaXHC6wfxkKG2NG3Ign4cDO5jU9qhsWQMAw5WVuzMHKkHa8WF
LzCjgXbPH6oV16nv/HtheR0jKNdf+Y26cV/Nx80txVcRGeLt6Kd/tUtt37KjGJts1eJICJjdhLRA
Sp01TBBxtfUPcgE7klLGBZF9TGTjkFFn4ZCX8OW5ZeuQgGR8fJ/auTYd8sO4kQpGrfLhp5uGvPts
oAzzj8Cq8PIz/co6qFxzgRJZKADidBPNIR2iD4S1Fs004H8gwDXAzCMro+JugSDSPw2l2ZGu9BmD
HgPn0QG//sxA0tHrdcF81uXyXOVtZtjmKQg9NVJpXJQi50OFrhF+o9Nx457dx4iL30SmsCuqpXcp
WG9Zy2LUPPn0qTsk8N6DNEZ8/IiogKZe+g6tohXlvrSI+uVKl2A2Xvk11za/wacHwS28BURNBtZX
kWvdZPLYfQ6C/kt0pI+vhTslUmsNRK7gtBc2dQ328zjXpgx8WqaDHgnteaYgUbubJpz4b6VI7s1N
yIHPnuIWpHEsZANLM1Hfg3voMZOsEmkfw9GVv0uWdDMRJLpjER/34oL50uHgGcvylYXx79gOnxuP
R5fG1oFibJJ45kd3qiKf8y+9jUZT75Jwcq1Alp8ZzNkLgzJuHydOzuXjdm7S2NU4sSxKojGJfPYz
Ub7KNCZxh25LsAggZyU07z1u3j91A8u0JaQl1tqlLodcT5I2ZPWzr+T7PxcErqIFp2D1M6qEc20/
1rEABgVMw7Nyuoc7sCRNStT0Xmchjav4YRGhdrL2jI5QOeqOOlI8GMe78JPz+wQmXL2H2/PCylmY
3XwWWX+iT0okJJWPCoMV+NF4jQJa4FyNjj8DpQk1QoOy44Jj5v3r2iX5S6cQbiH2wOzmt6r6UO1x
iKCrVGPd97t82CXmvP1ZCUk2Nh9MDC3ew3D9Y1qpmss+HViACx95mlLuJD5HViWodS+d3eA/KKu5
biyCfpcFFSwcdMeh3azwY+HnccDvYWvMuTiZl9XkXOIuC6Ygs+N6XMbS77mzyZSZK7WaBCfT7Lqe
+qLOVndR/Ts6XvDfrvJ7iI7pME8Zxam9S1mnc44XHxp0vO/z4PN2DDnhQd5mFm8PqUFAkl0rUcFp
PLYrIj49cKQr/WXNtaOJbcXKLuRiFGvtVGrG7Puyfwwbo0RO5akb5nNzuuHY11aEpDCi5Y9OIuL6
jPntXKabVYj5TG8g1AM75RsL0DoW+8+HNsnh2cgQ9DMBfeVi2YvKy7DyitqZx2MOehQmpPYdAgE2
CaNFqqT9iLkcBBW77L6O2f5PECgi0JXXhVLCSL1pIaDTCBX8BUFSQuARt5oAhoj2zUteE4FLmmYv
qcZBD9ptCsS2QqmJTsIGMxiL8iKCzH0GTxIVQSpBC40Aro7m6ehdp13QCM8NtieBHfNKkALF4k1K
+Q01bt74hC9QV/uQjzUqfOvy8zKYBXxfcm42cFvcNRjzcfUbDTanNrNVjINnQNTRekGdMtw9uHvd
9MLA7E0rwo4AfDcjjOHi1liDyevKEn4UlmrdlGxpzjAnVLoFPqzUuG26QnN2EVHPy5wij9HA/yjH
j/qfDW+ApSMde+2hcOD5HZ6580d9u+ZtLgVbD/lgg0MjoYxk6o7QkKwOql/xtWRJCGrc4zKJUneq
UpmV1DsugYa1kQ9IZNVgeJQFtCFvjLxcxxrCPgIOMJ4fqKAAXcyGnU5EmTl3hDLqxKj8vzl2/BRI
+rAT6+qq6hJpepCdVgMi/ovDyuPwS/T0Z0q71T7quA0AWO/W4JFkJeqIJod+t3CMWa2v7DOFkyjI
L3STnP5tBsLhU3hMolwA8cnqG0bCByAMm7lTyZ3do+sIIw9mZdulThNoi3SYF59ZYM/zIVBPLri7
jL118kkDq5A3cDICW9G0UdaB+dev5UaWIhBtYhidBCB2ZX/hmM8F6umEQ8RKbu5mbFzPAgm+mKcN
vIvGMDGbmexkH4CsYKJdKONfU7XOxCZsVbJa6OUrYquHgumLtzAIzU+SleEJD/0STb/LAq5nDow4
6qm8RfCDIMKuV3IHn4fuAHOiSXf+ZRItBKUao64CjjtqxkOTHLYALsNVoIUXB6MSw19SB8kOi9Sj
f1LJE4JccYoIiOBo+7Uhd//PT6kkVIyxqc6HcedeXDByFaQvzvoY2PkGd0A5KFWOfxMwAtAu3CdV
zVpEn2PCyEcpo3tlALZ8YEPX/JvKHtxZqGcXlHcpvXHPx7FFmu1W/EfSSTnCGRrgXl9pZeYcFQao
I8ZlNdNg97LL7RZXMMNQsJnvukUiYVZdUn28iDrO6vKHptCXa+5rM1niGlg6z7kXmz8m/Hsp0E08
cpwe9UyhBY7OofrLwne0trqBzk2q+d3yZIaIfG2JFZZ1TDeK37ZnvaviAImm1G5bBVsn/9kOPlbS
vG8f+x+YTvaqXtPp2moEOcFT4EBAcgIbPJZozKOnT52xOlKz6EE9pX3mKWBITUC2VjeGWIPRePUK
x2iiMbjMkmoJcQJwSPoPIY9U+DC9RiiuEWqGkwes3zMm45DK+WdvVe+jnIu5wtPJ8c/urbHocIOZ
ij2s2t/V8sVB+A5Ll2mx1DHZga57Y8kwKZqrGUEfcIja80R0A5bXboCwN4uVvQzRwYVMkobFP4w6
sHVY+nhjm/u/LsF2APAZ+o47stld3fw22AFD+c5pALww+N3q7F9UkY3lK9/hvkWQM/U42Q1LAife
CfoU5KylSYXVtRQ7I7k9Fpx0rsH6GwEMDhFLFi3hZqsXzxiJzl5VlwG4NUMyJhXMf38Ws3/3ovLY
91kTKPKEdMAcbBbKwAbLcMvGoCKJdqHnHM7nq0Tj2synnsba29PyhfiW5UwN5/aFWYjluWaHEqL7
ve8PcQWrKBRonpFIvulI+EnyNvWH0DHFEtYGwuwc8y8I2nlqc2qUEyEFVd/dRBrpxh9a48g2ChTJ
DI5L9J78U6tR3tciSMdINzuRm/LbRQrRg5vg4nPkLMeg6Qv+hTtTpeTKoqzYcbS4dfSp+Mu9BM/Z
15CN0Z5vU5tUR8n1f2ijXVhhuV0E/QdnFhGBuWQQzC4CqLo4u3N2clSkiu3SknvtWEcVcgV+/zGL
pAnJlUjO7cB0LXTSq1EGMWDo6+Mt+Z808pDkGGu2FmzVCH15OIeFge5I1a2QWTQZ8jf9L6oGxXbE
VqKuo78a5yhtsaxKpvQP1YWSMPaQbb5GEBHOMnFGP/oc5/1BLiviYJphZhrMSoPH+rZlXXZZ7cPq
8kFxVH3bsYPlXdRcBRiEX186Pe7SWA4UnoJo9xUdq+rvqdGCmbWfF2qgfDaH3N0Pj4X41Yh6fzTj
zDginXV9ambTGetUVkA25Vsnudi8lsm53kG3nHQqnnM33b7mSuiFEsY/3eD2xRJ/KofJnu0m14Zc
AqrMwosiFN2ybk+SIPBFfYFgtHg0vdIHI0gpSuk4pzFPcsWeIL5G4j3+EYManrnQrkHSNauAAgeK
jYVpp4v3KVZLu7dPqMT0HlkjsyXz304q+xiAh/EsRSM8F0215o2fxgWqcQgHFBCJSUrEH/yjnuRp
HszYCJSb/LCYC204fZkpaV8101SI1jjlGPGj7bFGBXAbMpbRUTsdrrbC+QPJbmtPHuB7ClhZtlKq
5MXsS45hUcWLm/yWQt6eb+NpCW1rfr2TfrhYV7VZZzMxZJQrxx2ccvCWUMtsiEEkdNin71HqzVRs
mayFanwDpE3jRegEDX44DEWuL7j82DEhphOEyqGyEi6cxS0WmzAcIZlRjW7CTfDwnUm0jSSRynVE
nijzfD64LzbWvyfD+uQpLjoWwty5lgCdHo8PImOpy4/7jL8vnmPcL4HbN0QvKPEPnG7638mOUO6G
Ip6CTyTS0c0KbHbapasLeLD3kcNCXQiQQ6mfoylnqKogktDwlejDTioV3hSA2fPRq+TGArY5oisA
FFmKikTUbqVfPbSzdmE9Qxgwf4SGhB1qusLE+juGDrSuSprZhnNKSk7Fku7phXkKdnp4M+iVBW09
z5ptyE+XJknUYn1aygwaOuROJqXNu3BN9Y6TPjC0SbObEMf1pBBmw2lhNKEdGrRF8PiTVcNjUAnq
w05IomZHJzEaUS8vc8tPcgOrTkZYf3+SMJd9N0wSdEeJxzx3Wa/MVwUzfDZHgjNDq4IIlw+W/b4n
ZFzeNmNF9t04nz4CE/aAgPpYHzTZCHUZiGEO+G6bzJ62IEGxLFiKznaw+KMhgR/lwI0LxvAVBDUV
TsQ6QHRsLXhXVoJBjNRfHSTG5gy1KZLLDe0LGFVnkgr7iorQe0ZdIvDlkvrQ5rRa4u7e2yv8ZIYp
Vze6Q/TFNktswO9dWpQIxEVO12TUGgX6wC7f2fMnz9WrSV7rH3CS2WF6544Cv5fxKE2ASG4OG8zK
kKhp+b6Rs5lk0f3Txsnw6WmVt1sXeWv5QADkQhXZPGLrNNu1dFA5K0SHH0XlXoEYbYEE/bdOFjru
mzRKYVuju0sutJFAeaLiMG4M//vkX9WFZyuNQZiZ0ndUjHEnL/SxwXWBKddXsBR94Cc0adihjyal
KPIjeU9EkwgLuaWuxct9Imx2K0TFfRCGwecjG+poxHBwR9by8QzPOIjjt2yMkjBbDDy7VTyItUMb
ab8o1E7hdBr+7FAl2GuLBts5yk5UX/qYCYbChorDRXyZfFDRRPF9DKbz3vEEHU79/ulsbpUu1uUs
avBPv9p5fV5onHdE2sr/V4c7g06VFzUTlWmJQZrQ6trh+8H3yyahWnhtItf3OUUNLTVKZWoksqic
Uhp/ZoxsI0esVuCVwT6RprPeL/13ltrfPy2qYx6pBwdhBu9zBv15C80jfxxlJcYpyu2xUBuW/KHz
NufLul3x7jD4YVJJHAKEGkzbrh8qhgLMJ+oIdQ3V5peaDzBhKPR4Xa8xGt0zM0q987iyzAmuaucQ
Nf9XKCzHSrHMX0UKgNYudiB4+6wI47oeq3mVchOYu6t7VClKbusaxq82sVvVteUPL2XLjBRcZ+SC
yBTN+P5U/tRwOV+Rx2gxRCBk8UkFfLns4j8TrlnFcNAV/4v+KV5DM6XHHqZZzKJNG+HnP2dDyjXM
LmWjqJ+kckYwyTneClehWyc+uUAPNJObzulh+RxmVgxP+wnBQq0QsSlnMKQ+DRKwifiWR8wqTWcV
u9xh4j7spFyY5jawoIoeUik672fngzcmyPQlI+8oaF9e8MoWTVcq97dcXC2WHdCXx1XpBg7b1/AC
17IDRTE2uM7QancgCOn/xhFBA3MScQTsI1G31mY2HhuIVMYrU1cYrF84pIxGJq0IwupLKsiWujtg
gHvxoDzI6wR1gsSCu/e3miUDAkmvrWxgObQZAJ6EYkYwaCx0GHkqxq7oOZOaTUpGX4qRUctQAf86
vi4vekn5gjuUXTWCHBLx8U5c/UaMEsTq0RowRuy0K19GIShH/jWuB2ijS7vY2OySo8KEY6vtHo65
CUdPJ0AE+ujTOi2KjmhzplKyCOkZsQy1/HQNKW3E6BwlVhVEirj9iQFpDzMW4UVeLmDN/sG2RGRl
dF84RKWlf6zUzmW2WlMTT51p8X75UTUXLS43D8r8wFpvtlilAvOAa0RfVKdKAJQIYA0Rv4adaM6A
D59yNLQYkNFzUluBMNNMk0BIBMKtEgDirBXJttNcBVakwMPQjtRGQ2gLFpr1VtYMSB3tJK85CxnK
csaF5P1lUhobOLqfoEcYhhp/qUesKQmczW2y1EnONY2yFHvK5kx1HEh/2u4ew2ou9HviRtzf6Rbe
zxCZYoHGkCHJ+ilb1QtHz/9iV1PxdqP1ti5ZhVzAhXZP1vFZr/qiheJBBmugSB++QO3zEPbGoPEa
8PasOmiO6qV6Mc7/JS4aADx04JYhHOiSH/Ulr0aY+jKX+sSq/WaFgLBrUUVtBW7LM+yOban51HJA
6/G/np7EguTrlujAqzR21K/KBciPB9Hyp2YrFwOVZt1o/6Plq7PXbV2wpUcg2JPc4MS1NKenXMP2
t4B9HC4hUkKWc8Iq9kc27XXnKGGdSih3AIDbjPOsAr42Hf3R7todumXGdzWQtRdnRBjKIvBYgiEp
LFRqJJw+Fe1fJIlAYlO2i/pqVSdv/br5dvlMuEdZ6YzG/5ojlCTc2C2xe+T9lV/QK1rRRyzEGWHU
SKLBCEz3w+jlMfsl3UtTS+9BVrgwb4zzf8HC3VWrBKHLUYkt2rwA2PIJHEPLBKnEgjIvQ9YAlZ0C
WlMqgs+yvTHNxQjSzoan+uWseFBG9TPBzaZUSZQZZXxFyZAKYZK4IdXXtQHXvzNLXjt1vXnz22nO
fe0T4Z/LyEBemH6MuaES4j79B5EMZCeZe3FrmjbwAgcCs1KJcrensNE2Mr9E35R9650jCm7V1Wc4
jNxuZKY3xiJEMG1Id31GCtcuJij1bZRkx5pprZBin3h+RV2zrLFJBrN156kH3m+Aj1WtUAdIXbXZ
YFrGN+kpKvtnREGBAXPIw7anwCUotDbTF4oaNf9/Zvv45I5PldREKPGa2AQFpBp8lcQQqU4aU1ff
NETg9AKr8G6UdhRdoTEswGYW8z1uZxBg/JHQOG4lAmS4d3uHtmWkGOfSqEWwdQp6zxCdM8CN7WSI
dvE2mhc56utrAc05pmtM6o6DCy3J7gqKVfPfToZ0rhidZ1UPWxvucbLo7ga3ne7D1/SFTNI+VbIf
J8F8WRdkX/VSCNMp2UzeTvIaMd1C4vkT/66cLT9b83UJLCoPH0kyvWU6/AVWlgHiM+d5rM8wpJCb
4K2c7DWGXUfTGs/nvDCaf4kOlbL8XJIk3UxYXYkRfWtZva7sMlwC8qDcQ612c4RHcnza7zAFjUOO
ZNRe0OrVfCTAsKI1PpFoz9sDHfoIFGzaydi3et6u7l7QHMZLG2F5wUDLrd+aT+NL5qFdxkkiMTiJ
w1OUcb+kAIWYbC2ZIEjnG8HsibSa1J9v3KRsl50eDpoTvZpHYNg+2NVNaHzTvITzPym98OzW+wl0
L93SE3ETXFLpaXdLd8Ej40Mlj60UXf9i2RNXFHLeeqcjsOarW+QwoZeNg5rfeL7S2wiopFdVD2P/
APFP8rYLIK2WNUsCLReOGQve5LaoucdS3xeZM+Vyp5tT9n5LIDBYxT1DE5lVy93HD5BxSkVW8ujd
rcOc3rKI0tYaULhI1kvSmpCk/8s5m+8z0Vkh6s/9OrLnyEt489wE2MdDdYz6kBkXtOwXs96iZS2J
GTI9xlv2/D6ZEn6D+CO4t6FHr4Ay46pa6MFBwTgyncINYLUjImcManp7t8Rd3TtYzZJam6l9DHcY
wtPQ1UIwtJXrOidH9XmqIKZxUwEGb36q3aMBQHBg3prUjnaYXqRT/NMWPz4GrfieM6kguOqhW+YJ
MtIi/3kHv/AfKKAoxC2j3t0/DxdaJ89oYXn05oVJ7Qlwiwfb9vkUAM4Eg1mZZ9867QcQ+M/J3gzC
y8iEfKl0tawFKUB+61kjTzZwLyQudMNy7VgBtDxOsyzk/1tzCHwo8c/fmrZw8IOUGSqaxiwaCpWT
5DMh0VvF6XFkCN2uI3nSI6A5dHRlf4t33Dsg8KV8g2tEJzIUZdAXgLbjjraQ/K1uu+VwIJJN5vs2
/B+mX0UjjwixZ3/wrQJ91plcHKpTG/S1IOw07gl8DVNlBqzSBsUXbxJK10nyqhfVcurx2x8CGOL9
SGAT4RxTeLxGfmcnSN7Hme6IkFCRc9kx/CxulrXqH1B1fZO7A0WSdHtmiLzoy5mT17dHBYqZryBS
s/AjsUHKOQJspeM/CHScVj/R33e8xVPRebgkANYxgDsCokCrgldoCEqeGmN8b+YaDt9sPZf+tkRv
6u2taed09sK+nBK0i1gFAWJU9ErMlRguAE9HGyo4Ao1+RsXTLmIC+B3zof3PAh+ZNxjo8bK3yyD0
XuDvdoo7nOoGmt9i/4OqH17wjaUOW4PrssT4Ty+c8OP7wKAUuK56WGT9a1uwavfT/usmQg392XQ9
UFU5crb63381NSDNbfYbNPlQln+FKFwSk6I9NMxY9MvOIQkPpWiD0ZGW+El9Jmy2aJC+FVuJfVVU
q+Nn9/Xfd9SSXuowfubNEt/ycrbTwl9Lol+NGNdqsuMrxpsMbSKtE6xSeMG5oklkWHXNW+MBq7eN
Xaig4x2UnzcjEAvTj6wUghDWC5r87RyW40qDXTg6OFev1i5vxQxCTZHctWT4u6XZvlwan4TDdSqG
+CmeUYUOVr6eJBJMrvq8aLYtkLgMeGt3mhob5jJNf+iRAsR8mZwLizv/YWXN1klMk2D0Mcjj6aqC
gpcZTgxsDkQ1LPSAaOD+0EU7fYY90RPe3gW4i883GbWDtIcxA6BMRTa2O5yhqZpw+COgQBapxxxv
SG/zI1404Yv7hJu0AxUTWZLoYDWHUt5PRDbhasd3kSynfk9V5RXCl1QsX6fciC7a3UHQLQMiy6mw
i2JY/j3/zdfOSEYQlUMsvUVO9sCcS6SL2jhbE3zSwiVHodzPhcGC0RjdedLyfmnwviCQSon4L+gk
LItKbGq9TUNPutwSPpJHB6gbGOz6aoLkv/HXihS7jG715igDRsm9sXVVhNOGd/3I7yV9wSzNeXIv
IOMFQA7OwpTg7eYf02An4piSs8DdhPHMhZpKofpy9RHshhbSD2uDi54xBpq/+7WtuKd8otgC4iNH
pOFLPkwBHPXLMX7aN9HZqoXcOh2HMohbrgQOBXVr/nBCpPDfpMMnpwMKSNRSsUYlSwbJs39Dnuk1
h2CgKjh07tapH0kRvnM2RBaz9vJo1dIJk0FHXedqdRn8q1oiGgYFSG/Xa8IoeRfcnNDfh2Wj9i6L
j0qhV9Ifts5sAbb0UDVEvHmPSoWiaqWSPzSd/h54STLvE1TeTKYKmqdphNat6yhkNrZ/gxvlhVaY
jW0iR4kbzdRNANQXFTrBjzOzVJF+YJ2/1hiltIrMhHeCtu0QRhonuINaJY0DAfIhwp6+li8s11OQ
JahsFFhc/JgYC3GlpcpMhECvLkcyHPAb9XXOHg5G7vZXHKV3bLBTqdCxmfkvDOQUqwOxv+bZ9Xpg
evKAjiR5dqCTDc+AZVfJLgh8F5fXjYbEsjYJSVShv9EuYuFZBqa/fVtsRDTahd1W0KUsbrbxFGjX
WOXRJ67QAVbO3LQ8V5x/f7rVw8gQU8VoEoiA4dN9x3Ziaek+IBnTatJUvdLHGfanoyA8detEjYBH
LWDEzVrt8pqoXgOIyOE4+9g58Z+XEhfqruXB6/G1tI0B7zcilSC2b5sBcFlVWNKDsTjl+LpivCVT
3T30D6EZQoJ8+AmZJkDWxNiH5yPz+2r5SOhAClr6v8n4UQTRL6yDKcnjFue0V4THCWcYs5vSO5wW
9nVlvptJHtpx99DYPI+9Vg+ShVYEjU5wufheB36330Vdn8IhHCvUi2pmz7S5gXLpOieKVtEj1wmQ
GW124aeqgYv1L9lRgGhGg5LgRcYgKT3L4QC7W6fS2QgSGMWmsO5hweyXlr/s5fbdFxXPYDkhL6C+
lP4vGo3PsjJWZfXGP/64fj9hyWjTStpffY2HrHcMaqleDXHRKXwSf4upcgnqCbPSuD/XQxBpjIhF
A7Xwm3+ccY+cWbBj4rcfL+OzUNOUbBFOLTfgcb9jnRCWHfacPE++bh36+THUNNBs/CVimU0kTM1g
xjZc7E0lhOXnEICtmaji8uL6Lk25i1zQBm/ovreieqfHGsVFMtfgFJ8V3nd7N6luRZaDUX2n7Q36
/1n80qEGDAOgDbXHCuHrz7iKGYCwS1vPaKhccehDK/DtZlt+NA+/xJ+PTDlw5L3GUtDkK7n6podq
g/JaXaaSIzjpXBy07ZcR9UY42LQK/2Mv9qrpcjULPWjxim8ZNA4gi2cN3cNkfpNh0r+BdtD2E6I8
CYegDeRsE/EvgQI+j2dxCA0M84hACdvb2y6aEVQ1KfzI9J5LUBpEnvHliGjHrSeniW8tPoBYZZ2e
6RyD+vN4Eht03JW9ZuHlu7T1IiL7Ay7JeMhh+RX3DgfuPsckkXcs8mOUzlxxVcqRqXPY0zS+mV1Y
arKyOHiVcipIjhF1wB1mpFTuJa10DnDSCpk8IHTnMJM8KHO4473KT3MQYq+ujdrDvT2YrhJ//90b
ENO2/jmCJJtcSv+CxFzuMa6uSIHcZ8MgtQY1ANETahtpA/KYlAZvRtEoILRM1vLLLaeJKselsecj
rzLZ6dtNTFvAoj29yliBup5Zi/sbmQBXBs5xce0+xxlZvK7wD3lGjScXzEU5qxE7DQLIOqse6YPQ
S/nz5iYBWhPF/A+Kc/c7MROkXFkrStSj/MJRhztflt71kcAaT2ntpY9XNphJQ045XWRHorYk4ZxL
ulwr9RK9SkdLZWAtbfTcxRaHmps6JjGjGbz/y+oTw7p1rw+LlqL2GP+pAIsjwieydHaEs2rsVDHh
/uPFATuDjO6t7UwR41Xhf8j9lW+HDULklUigaGSbuxFUU0QBPZyy4A4JsFWw5M10c/cYA6qb6G1a
WXU+2Gy7zXx7oQ3Dphr+XafO6KV/tmlJNVjRTIth1hFVKD71B9ZPbmbv4sj10r6kl0oaOFL8DPGu
YNXUAFk1VAVxwDzzZM9+GdmdTl6eBzEGMWLd/apfLAVpv5/VXg7YPSLIhqIDtT0r4QBWSRA3vozI
ZxfxdW/NqOlHNgxFl23qDX67nQWNzKOzCwNKJDq96NRthOapNqDLM8R8uZLWtwh/g1mojFPXkulf
oKrqAA9eYCSz1QHUHdV8BsgIsrGLlubWqTz/29PBfY/NxffEZaMKmSyOWylAtGxRqKROYOQK7N2C
BTMrg3U5U92zKfhmHAxmQFXFLhQFkg1sfyMaoqU5iLXCYq/BlmspKLyf5Zi+rx9xwbFKgB0g6ss+
GVfl+dTibtf4irzhLiI5nuZ9SLCq3n4IqjPKLDjghyHbflhhuTaXUqSlm8ML04j9K9Ix6fbiW9ez
CJwiucAywFFr1y4iVw/7YMKx15QpFS83+DY4NVAnVzAJbeiZZV/uj2AFeHnrms9EG/6GNj4ag6Re
W/M7itNwe36A7T4OmoZ0qMtLz7H0m/MIlnFqEFXMmsMQst3LMYq8ERA75Z2w/oi1vwHu6PEL+Q0U
bT6O8hRkiOZvcnurotJMtMJ0bcYnzy3dawcZzKtVoj13RnCTxuVzeu6heVxp7vS2W4VhQ6mIhhbK
vedQKnkPIDjn8HqatCxhKFzGDtT/LytVBkAmFtr7xN2glhsDwfaH6HNT1fN85DTh5C1jFd0I5wxi
/1OtVpRP8QHQ9BgsyjaDCSu4zaiClXoaWvew5owg9PnPCpYMz5nMDTMoRQ7YlOEcOwpwnu17Yj1B
VcZRdIZaDVS0pMnXOawqnr/X/Ro4nPB5/ns69s/0aJbdjCIBbwFmPEeTjJZC3nGlc1r7MVP/Dydm
6gYoHFoFYo3b+CD0bm0VyDECoqSiYrny6VYg9SJRB+ADlCm3YJBgfaLRZ9D14k9/M/LejmM7OI78
+x4MLmcLRdyz4QxLu6gjgdDsd+ed+/dYtiomfUAh7EQ+WvOjdXQbBf7T81ucFrqWlJJB0S7aYk78
e3GoR+aWxi+lhsKFilyOZ1q4QFjOn5AuPgvQGKy8eGukFUNYtojbrhNuogrlfT3BXuhcVf56+FeQ
Ltt9YyDF/BN67BHqGekjt7s6ubb0f+80Rj+0CEr7M7sPMDoGiYmzLQTDLWQF0XmimNtE/I4aPwg7
VaZYqGxIfsiUXKyE2hCTnNr6aXqrE7n8Z62wrPwVFOusE8HcRWwEq0pPplKKm+b2xkBk4kL6jjCO
zTVAnrt9vZaJWhUldxxPPTP7wKUr7hOcf/NfzDhHdh/MMDWt4i0hItO7eDRx6XOjAzDnh10iAcbg
6aXTc0XmlSyU5Yhn34EgFbInQ9q4IF+u4a9Rt8dPocWSwBhPKVgUhM3bGnV3XGOXLC0nd6C8vije
Vz3aI/wUbaAHAHSD5AksGeec7d8A81DapxsOQc1E04jhEbBCUcfOd0RqNTxVlXLWP0A0u0ip4Tcx
891qt8F2pQJm6aLiy/Y4vY84vpxmD3eHs1LTGEAIODpGWg5UdRctOu+t1BlU4huRFl951I0eFXyr
yoTf8zsBgAkphIvG9Dko6B6E0sT7BW91ySAXflFLVEDDFBq5Q6iyQa4vDL8lpqdZnJga+muTUhh2
PGkRGdWKUAtnfbcISCV3jy6qRk2HPFkVSIJPK0Penr1Ffe31PKHEigIvSHintI0/8PTmoO7YzNT+
MGDqKltXj7zqcZJKSRVL3ojYSvPKkAWPC1Z68J/QX/+vLIo2agqZa+z6qGELpDj95ZRptxiRuKy1
81MPIC8P4M6+rUUOftR8MIkO4OV0A//QkzeGPtITy0qhO+/+1B7OxOw4bvRXsAGyb+koyFo9yULT
wkXMK9TA5VTGSkDxGNk9Tiz4dc+jCVatPEsK72pXD6318+GXCzR9L5gzujyk/m3Sl45uIcQHADBY
+FIpaic6sxW+ZzirWKGfyBXBf57zgjB9Y2w/wvyFP52kDHCQ/SJ9f3Qs7jh/aObbII6mB3roUwjq
1mPmgOdbzFx1nr4gMZA7K86owex28U9L5U7QTYfr2kWdVshAVnVlE6UObNNw8/dlIczGkwNsfsmd
Em04eXFHQ3aFrmjxEl+auGHqgAcyYbsddPoCzmFhPIHnQ4WzbmsMpc9CK/W0dkm2tcoPHJzjYJ2d
Z2MoZS7oWZ6I+vYhDu1eZrzDuXuKLDHePlXLfYFzhKEZ83UE6AOjdkeXNto38vV8H4k28lygaNOp
3ZfZIRW43ZeFidVlemwOG9se1p1PVQNrJ4ZKwZhKAzPMmRbZI7GDtEebdZqjerf0PDgcH5lSdqdt
v3M/duESVwnBpDzIpKE2D/Ql4UuwzUE+0DESpkHiLz+jYfABNJUNHJGrJ3MUz8OEFIUvtKdVXqp4
vaPcElGyjVvqV8LNqZQWXZqFrc+kHAvnkHz0wbmqVz91zcifdgTMn7/wyTC4UTUJf6VoXUhGzAxN
eVZEBbnQWEFjMMo7E4kiLG4DWsDv2AoeypQwDVJL8ZjK3T0/oRX+gnNYl89y58L425E1AipDlBLF
QU9wE6JzsEKLjznu7s2Kgo8k92fHku230RfYSJ33xLWg10zIEwwcA20/6iOqQVt4/kdI5agyhMOv
NVKG69T2mBbXedSDi3J6VcnAa/gA3Qyux7ZdhMfUFOFRYFIH0k/VipZ7lM6Ems1z+j7uzG9f3477
k3BDm9CuPx8GlmZd1HZ/eBKIphIlknUh+Wab4mtX79V9uuEcwr8lm05CcYS3w2jSoqAJ695e9KU7
3O5wVvvquH9zP/3UyBIo8k9CX24RqUrsweGWsRX7zosJtcOxdRIN/daA6jxkhk8w+CpaZKYInGSS
2LMZgLVevDOFNbwjY7m8K5KxiT1sSsrgswxFoqOEon7yc0Ldgo6XC6G+uyAhLNYCj4AY3Xk6Cjh7
HcOJHFaF/7q5vZmUKW8wazspg+dCjNH1NuLr6mhC/2wyer9X4IKgDpFY1jHunF2MGEWSuRQ/7gWh
IjC44lRGzC2J1zS6Gq7upSxf5PdMBL2DhGiJyejFiPHKlKBAAiB0TitOIpF9voi/YkMGjNGNI4nO
Jn78AYwmNFYQoE2M/GtHkZ6SNuCnEkNW6sCVpVzyzLfbyPT477DYtcvP189L5TyVSGPxaaLtbMt6
D6YOyi8Xl94xEK3Xpv1Do2jQCLbaTRozQ0SSS2jhY3gGS34S07uzdJYyCq3ZfILZUMzyoNbB1flT
5XOmDMNtAFzK+pEt4aG4uPKOXDLwwFxZ15k9Flcv0ywPiGfftn+nuWbiHKHdQeIk68w8zycA23kE
iNRXj+H3NmamFHDbW3dT16S4Eb9DAwHvE1RDewJaLtUo37NcJc0QpNyHi9hEmnB70oAwz6L7M1ZA
jFlofF3s3K5U8KQkZG0EkxBoTzCsFL+wrgQCY7F+LiZ2Sq1VrFHRIi3qJ21iDHMYjfmTnxO3FvSw
IJ7lFrO7wrGWTXjw1TQ091sRwt/kk/S7kKfwIFNZovGz4zRD9zOfpS/fEUsulQ92JeDUoZ9fZLnA
EIFCPt/qJbVSu4oSKUR0789VHNaMo0sj1jFe17q+OdvhL6gJdtMt3XCPDha/PIEx9hyLwwYQ5gG5
mhmZRmtgAWpmpPhEy0Cn0Tx/nGBvgaizgLeFK8uxlTuwJhm1DMKTZA7Cv5nHo268qMS1gT9lQb4d
2Hbea7kKywR4YisF/bm7d4MHul43plTVifxM2Pq3dg0Cit+F69YTpOmnXyzgM0GFehpoL4a0gWfw
nxv0xzRLNVZBt83Si2+H+KTlfSOf0JFuiqQhM51/Br3uGfI/dQ7hxzMZ8aCXWHyiL0r6cL9h1hw5
zvwt9bVzgb0VRhsMF/XpAvFHTW0NklOh/3gzcKezjLiFD4fbPuhQ939wMW5bZW7nG824t3jBENcJ
5akYr1pzNrHibMBRQTvLhOdfGPO79u5LNf7Zzotu4qJhv6L92ipYH71F2lbsygLwtPU1yQxgU4wP
sAhRfVmUupWm12GX55CyX+BTff+RFAdn6KHQ2IlP72+/5W1Gyq59/bkI29MMzueWVBIjAHyQYkfY
QDfL7Fn8blv1aMiNhvK2KUMWSDBYcGtlVklistMU6a9B6aLTN7tNm9FaQ+yDaT1x1T/wNggawVjq
KbA5+R+Xd3PoyM5DiZ+9KF9UakLNCEwVAwrWsFUpu3U8shKBt37255v0W/H2RPW4rLgtl9UQMCXt
MN67RXb/YgC1ZEQot6Zln1SnFS0dOMBaODuzRZzmguHUtchkYeV4pcxvFX2PL+BPsWMNBlZNc0A8
U6BLze4UBOnIEZyXIDhjrP+Fxc3CfM0IJ9Eghqk5R8yRJIn8L2o17488wNaAZm6N8tH3y9p7JqO+
yFn0HGGr9QREV5xLDAbfPy1U0td+3keK2TAlmvwxqTvrNBbF9YzSvcby+7GxZx9Sr7J1/DGrM6ln
y26gGy44U1nbvI/VZepHVbmhAGGvlaevJMysxDMLb6fwEhfInB362ZimSZ+Y10vBspbsggGIEKm9
C88ArgFmWrWCkX5fuy6Ry0+Qo5+NlciZidOtNPth3ZjmX1HmP4g8rUooyCepq8jV4slTB1GixsmH
gs4KyN3w48Q9aPEySBK3Pga5UMvLtDuIAYoR42pPtpDvW3KJCI7vGPOFNeve24YQ3eMxJuPlxir6
2vdgg3HWmOu3cO/KOl/W5ojhOWRnaYSfiIpdvPOE9GtIYYnNRbWm3H62KqdZ2cg31JhPlBOsKcbv
Pb7yiNLAM8q5vDX52i1GPDMS2zpOyowidxTTCKyVrycRsPWbHHxt0jWIaG1nminpE0/PCkNcZdBw
+V1pQ1poAEI3JKhdl2/UoZQxmNJUnGIFnMSEoR+z6Hs+c6B2ElcPV/A+yBPBn/VLKMOYdqA1iCWl
tKq2MaLw3SJLuMgAFllbKMiPGbmFvv2x9qCYLUu+PEqUCaQ8S7h6LVoI26bQ3TUKA0gWrdAoygJe
zWs1ZPISuD0oNNmU9JlxVYDlbAA0/3KdTvzqRyqW/V18X6zB0iKSUlrI7tDBdgOg9FZQKdKHdnO+
FvNnKZlgfY02A+c71/tc0jWpoilHTke0RCS+ugdYldfed8Z6XPrYZZTgG78Zo9tNc/L+xpv8HeWq
Wz4t8GdPVPV7fYsdzYkmr+QhtueR08ckf0PcYJV3VevarCkTr6G3s9l0MpoCmjY6gwz7l5wSp/tE
zUuqHrzfsN6vpEZfsFOyWN1AxDnxfeeyinZvcacDC5is4yzHS2LwAB+zlaNOIr8zJj1F47FD+O96
Am5B94M3xm9Gc6/BiPcgIyWET07wghNTZr7Ifn5ocitOW71cztXM9bxmnrtbpel2kw7qat2C730T
NlBl3NNmoP58PvSCtdP+BiFqnJcuWYmiWIpxE1PZrpwB9uvgmRI5sSau7PdQdgJVzYWL5x5Blo6U
7tUiFty869WjdeF00khkeWaM3rGJBimz9ZaKzYiSnxsRz31NUlU7JyDjbgzDAI36mzn+yHSC1NSF
WK0ReMXnU5NdzERS0klZbqxVbaUHpdQCzgAegWJk3dC/I51FlstnPxe79/Mke1ipHCGIqPWzuFhL
o0yFhAtr4teCrM6VAIM8CQoRSkm0MwG+nioMhrHirGDHlApOv58zyW9xFdVZRuhqby60QukwUXbT
nYkd0RLsrlmfr0k4PbS/+xfM8zzF6qpLn8Sd5/6MJPLu1yiWzzmEZdrNWNqzzNoySvX0Tz6I0/pG
1nwscXi+3TfUo2Ddoc0M9fk5EeEVCyhgYA/j51PhvQbh8q3kJqC4MbchwUhImDt3dBvjrHkSIRYf
e+vhgi1X/jRdF4rNVR7aLa6C6klfAPBK19UhMce0m25r97/mg6dSKqY/36YGU5vrFqlIgRg3RveD
tCvg/B3ll/GkwuHjyY99BtzYVFlYICB06p+vPyh4xuLZ2ZoZvyqXMfYlTMe5qPD4aaYX20U5XrFu
kcKMWh1PPRPG29MlN24A/truSKzv66/CvMbyiZ8x+kvwEsxN4ddyrZaE3OP2VSVkTFdCy9VKvhr1
FhVrzKXjVvuj63EHHHwIz7O1EowNJNgmjhpC3+NAsSBTqhG3cJ39KyN0kg1FLYcU3w8QnXK5RdZQ
gOesULjSsFnwhV2g1MxrVFXKgobzGE9g9NNRGBkOatGFke8Vjd1+M93s1J0BCOxBv13K/k1IG/DP
xLRXIJ+L5a3FlDQD7BYWNtUUG8OyXTXrzpEZl4bz8lqTF1XxeLl2iAwPUwdBzUp8icZddyd46FB9
KvfJ+xHbWnb0nnD48OwY45lM8Jpv7dk10c4akApCbLaKTuTPvhJ5iwNkgAw+6pKv46oLps1Mdf6d
1+MhvIEeljUU2Ksweq8P2JHVwofVTCsDA9KGx6biKKYHQ0XglmgLLZpSRMrddiwEkT7BleLNWWbi
iA8ZUELe7tFsswdFc1eTkDAhz3fTrA0CTGivfybw/7wBJJuncTgwkQLfctKY1lPCH40CdpIu695U
GdLG5lmCj40wZBzdRQJuYjEik52hXs/BvVvHcuR1RMHtjk6+pG3lDuG9uHOfFClxmvocxsxt4GfQ
WL7u9EEODBpyCiPkPuC6Eiq9UWZdbnPwXPbEnDjMrKwgI8bEdcCwkCc8yYysYcj/loyfFCcSLG9m
0lBOKAT+VTne2YAWdOuMU/3KOWck8ETe4v/NmxcRgvgcl2r5LmefCwFfd+bbv4TTcW4oA9IIXj+m
sIoazeMiHAPuOPWS1v45luHUXXVoVEoHdrSzhhyEpGQzfqkfV00wn+UNn4G/IhkHyCYU5Bu8zPgV
qv5+ANuQnsUshGP55+fgIn3sdZHBUdO4UVEYRsCZqKvylYuIROqb8yVfQdSPj3mRz5q05yusZEvg
LlPJKABnVktmDOYQCUptQg5RU4tzc9NkhW4oDgTEb/9KJh5Ecs+SmD5g/jZxsOeB38Xkey6Yf9n5
prMUF+pnM58x/mQNSnsBsg73N3PdxY0paiZDjtM+LB/tF+0Pg6w+Z+rpNa14sWtyOG092oi6Tb6U
g3VRVSillynQ50Xuz7sklIY+4AHk9vwvdkQlw5K7DKEshth7ArGNbuqJAp02nLOQwveLJelNakA+
XoX+cAUfd2Vw+4D4P+DoJwbQsXWPRdKePybi+BZ8zaJ1cDc2fejugsV/gODoF2b6yRCtNkSc7h5v
39GVQNTskrUNPH1St8oG8F184L+CYw+fonn8ujAu5MN+ZCOot5YvxuduxFx5mM3Qgy5kWjYQzSvJ
ojHMYhnkLWuIo1F4M7FiaJI7mHD00tGjIgxlRothun98sWzbewGR6RCilu3YedRc9dAX7Oi4uwr1
xzIGJXVx4mh/wsrnYGBMVG2fdgZni7DwyhHvqZe6aBRZXK4uDNY5JgrWMZb6aLWlO+9kxNl7P9Q+
oH9k1avwYqdabHyIGoh6ZuLWYZEcNcMhMmeWKJo28Ew4yiSZ8qNmTQC8kmYx8OSXTnXLxCDc1IRH
YMWq8HsmRiFk1RimY3+6mLrN2fVJm0whlBPBzGw7zV0AJ8Y6+SjsjcPDWMExP2E5kLA834xBfZss
qMKtI/ESUqjl4NxKlynaGZKWw66TYL/Yt5DYeihDzlPLSRubpwI9jGLot60Zu817pmig1J8ZrFac
nyguJ/OPtJ7sgyLVOHZzZNr0aYPdT7Bgdnf8ZBJT+muLC/0Cyn4rYql/nuXTXshdjV9NCZjMfJts
HHjoBXsmZoiajMulSt7d42D16yrmIkR3ct1BGiuFlwZA3yXuzOuoe7sTUXus+a1vv9OOFKbXFHy4
eZzmMOx6XQeDFwEdOgft/wPkP3yflGAcN01xq48Wf/D7x7Z3Dq57kUplCc2sKiGjUDzI1V9GFGVi
sG70m1HPTbDWnNcyKcMo3CKdB4tcl+Yjvi9CtWkmqOsh2vPCbJ2GD8Ppy2oJ/bOrVkGOQhyp+PHp
l+4Ud3rahfFRmpUskNHAMu+QQupxG3pPOmyVijzRe+bzsjvWOGAAtuzE51l8gjWVO/LH9YjJ3ezB
k9F+BEti1+4Qx3f4U3I3Ym5ydpc3HjtIoyEYhzHNLlaaM/N01qQiNTNk4rAYT05VXhWUBiRqrJmV
6Qf5wnAx1RNlAuM3jNrZXjSNh2S7VzExN4tSM6QVsTPWnztU4qjb+WUpK2EgXsmu8gXyAnPMNAW0
AecV/3G0s7jeLAEbc/BBeWWOgF9Si8whbhy6nNAZTYuSUPQP7vIXAMxd22Iqzws0lkgVbuQfSnhU
rcnbBRTxDVTM41DFl4kbqqO+Z9rRDUHTzP9aHiP92erGDjn6S7qJIispQXM5bBL1GEz93rn6jHXu
ls5oQMDIzGtIP6b/ASUbSnG9cU7l/W1jO7G/yRWvAh3lqqpjf4/YNev+TOG5sQ9o55KCrVfg1p4/
IXurgT85rI+ZaXcy3xbflOpAZL5GxZjym0rFKaGoCYq9OCXUXE6u6WgjPHI/XiuKZfpt0BkpX+u0
3VxhMx+S2hHV7pAmYFErySqar2Bz8NyM9v4h2g09JOqyulFMrBrUU1Iz3y39uSBW6exzJJztKsSc
G1M1S09OS1sRrHLeNfj7ZT+9tLIjVWG80rNzNrQkPFkqs6hPw2vcQloTLQ8T/TQ2fL6OLR6iDZJa
kdfklYupBOYi1HAzxt3HiraWw0+ATYgcUikvN4VK6B8yNC0u6qaFbBotySgDbVSKkNEDMUL25P4S
AbDsLwnN6fMbc7gEtSO9SeZaFxFOqqCc/X7eVkxKRrm5pQm7qkH/CTHcY1MNE+uw1v8WxsACqdyN
uujEfVVSjfnrVW6sQz26A2UtNPFp7pozvywByJ/pjO4ae+WcQZSddvHCXwsEu8uR1JOpDjm9xPG9
Chm4pAQt/nY+CQ/Ehiuuj8zJFp66VKRkW/QNVFpDr93gaJn8btXnBxbnJKXNdM0MsA0jksyEHz/H
KOIzdqtAaZ3ncsoHGq7GZgKNVy3Y78rRsHI7X5XOkNZLrjJ5vNFDVfimuP/4tqLYLUxlhMCLcM5H
EWnEZjmPzMZNecJ+OS30INAINHz5/tpvopEzCTOegx2BM1M2sq8mBzyVmPtrfRve8JyBGEhbZO5p
jRTZS6rDdD/cz9D8Ex/KCrUTSrLPbHY3xq8QDi9Q/mxMp53XTKOVBFfqA1P05Dw5p5uEXRKkgJyd
jf+eYkHPMPI/vxq7uW9obVlGRvA0qdhaBqgAlc5YIuUL5ls8uWJjJRUozt51AbJ4BF3m+C3evj2B
W7mgYNwY/jdpY66JwM82KfIMgWRsxLtHwd5sMFGCW15TnbI4oX1WX8uLQ6cif8o6lVWyA0CmfNm3
kWGdtuY0ThkotFseWpdx187vRKW2z/BQ1vnb/WAPqAYq71KcKzLKhedQ7V3JIbrfN0iW5T4/ePj+
aCcjcmCKzBCxWAcquTsWIFhqfrQA8Two3sEdmheZRKXC/sGwz/gErY4x4+cshxTDaaQf2d82Ev7J
taupQpoQP8dq4D9pyMVGNokaeh8EfnJI+Q4lfASYtOIVJZFYMUKZ3ImeFqFyt6esUkzH6M5+Oa7Q
eLB9o+wccFhZMYfh86kG9hwd/NCTZDt4FoYedBqnHqFn30qTHuEvE/1ijI0ElecZoAr1Mn4UvZ9M
SWpGU7C5q3r8k4GESItVJhM3SdA065sV7g99xBZTMRVAIAC7BmM9eDbKfagDZ2ZM9YXXLNSKtZIl
VsCmHglHbQL2gWXE+tCp1S27q2R5YRMwsudpxxQzWd9lkOor0S1KqBclpEAv3+GypIHaog2Pa7Wf
26NLM6iMDRGFrLxNxysJIJSkjhFIDv7s1g87o/xz38+qn5z6jNE56s+G79ANqr7UkpXOqjM55ArF
qVH80619qz1TZ/nGcSZbpC0xBRc4DrYEDSzlVAToAROjPlTY4otdrCs7s2GA7E0OnG/J35vO7C2d
scePD+ibF5Fm0JormDv0cWE202Pasx2laSK1mngRV1d+HjSg9a+p0Cc2r9S+CyH55xwECJ+ku6F9
ePQ3fNMcW11sz3bqLHiRlCEyOLTlRSU8zeh8l8KCs+n7snl+YkSErZnz4n0Vn+jBB7eEeXYwUKHu
q9E/lNI+FCDXFxHkQAgeO8lveaqjPPGe8JDFsqppiXur0D8NzKZc2GU6DanWy45yvFDDrnRmoZSs
TPds9e2YTgFQqcfMXhjQVkcnSbElI4t4kWtnLdHBGJWRI+et1G0OZnK7LNqVprODuTKqDLmV9awo
3PRkuI1zzHosvmRrp4OgAG5V6hySGCnMkLZLHx3RrIpIlvMjhgvTIHf7hW76aKn4BydapcUiQfD+
zyynlHzLhCs6YHIcJBEm/R1YE0TxBuUVxRB6yi0LFsJP8jraw8Tiewhye8JpC8+fPhRJVIQbqFXg
FFdcAzlvBVm9MzO3LpWAmShxnpa2bKGmYCmSnJKkRXzV5ROTxAXVeZMBPoj+tRp35mzhpLoNQvN9
bmi/mqL8hIRKUk9INJDOivB6OH6m01CxQNyrILsITL1ki+FoOiqbYMS4RvMEUgGBNFDRnDiT1oDv
XUuC0nekl5WhuODwjOIUKJXq3RJqOWBTyVmlYlcgbSQM1btvvtXKprWOnlHqJkedGaIwuGkXVLQb
dtzXgGGjIA42Tb6kulrFVPjFLzpr1mYTs+tJZONiQLfUIHcg/AK4sIziliXoT3CYz7UXl8bnBVYA
KgjTVOzDBNf0TAMIZr7IIu5P+AxkXKIYsxS7TjPrk0WQqtcLFcpNrGK8yxTwlsueOdTilMWfmoPg
nFBbH42DYaQ29bSw7rYPlBl5n/SSFOjOrgRiv6h4Lt5pVRfRbeGNz4+tAuckfF3t+MRGd/AXZ6Bk
xyu5YtX0oejiazsFJN4H0qdxc174NAGVEongx9aOSbNt7SC/IgVuff103/PGVStXwhpkdxwB3/bM
RHjJv4kjLa+K65iBAs66owGo0l6G4TtPxO3aC6MusfDVb8itbd7PigHKq5JEoXLt0stbIHBkNLjl
xng0J6B3XEMf8uWvCRzA7SU6GrtdcSxE5GGn6BZjdYVuAaDtxVYYIbxopMHKV+sZKkjcRZY6Q4sn
OCWKRvnVl7Rfw/r2oQs7tuGkQqtb7Jya08BbZuHMm1xauS/FTH6kuW8PxtokozM17o5TJ+EuYe9x
grcKKZmE4uMZ6c/s2SFE+/b7OlJALllQcGOLy6ZPTCsJDQW08j/hI945WD3ZDp+MbQHhpn8tGSOc
Veo7YJI2kKQmkI4t6HNk/aNOfd3DJfw7Tw3flx4XRVW8MEGaSLd5pT6L0Z/IOS+1QQWbTt5Ac/d/
yKi2AdvAy3Q9TuAgPaADniGaXfD0Mw+B5xkAZjne+WPnIw1DPhLLPmPCiV1ORCuptCuONoWb50Zi
cPh7vXEqBhvky1ODhzmMpJp6fPMsSJ2C7awIRTFZ7ktgZ66EHzVhtcAw4ECXnOOOMb7ZNJAoYY2U
iwMBqhNJDlc5zKILpIvLSiQUmhV8RCqJL+pX3au41xQTy6Ps0T20uQ/46fv1tFd+ngkzyjIbCNba
CYa0hbp3SboLVQnD0hYjov49+d2fyIUJW4SSI60Aqai0S6sUvw3V1WBO1piaESdLnHCOnMnV+NSd
hfyfdcOwa/Cc9qHc6h3o22IhoLP13RLl0jmgbmYExCrWSFzonZknwWKIL6v7C9E34Dxfz0JEVKCr
fVPrK3AJzUr2NuC2ninCpzcUyZWgk73wjbAS95jYbXXkUo+D5nOaazB+9SxG83X9Kw1MSUILUzgK
1WAyZIRZIAcoGA+kfsMEyUevjwlHYM+qCIAoAJJ/7pYTxzPsLTWQzmhsp3bXChArmoW6ZWjQ64Gt
dIs45PLc5gbfQrG3M72SOSHfKtXvrDAmia1OnPFXvQAKq7o0gQLNFAVloW+GTUVPJRLIwBmp93af
NpgP+zBGVzvd2Hi5cv64qRvrJetRSkdEki52jnoqcKdUdHz4I2UvZubb69aQdUUrsZnZjqsys9AP
qujasCgb0hHcLjjXH0lqxo8eZAfiEKIp7fo91acIilbP10SEmYz9Q+quJri00ln0Kxs8xulR6uZb
19AYaVcnxfjaRWby3HSgigALaazMNhpxs4B5aR+ruhq7OgNPz1z4bPW+PD1rWV+xJMUoHyZb1aEA
su5lCpEZw8I7vkY3ilpHQIigzNueXKRs/0WH9UlA31eeDgpivPjvKWkC3v1lzJJ2dBeBrxzLl1KS
XXLzO7xS47PBMUzntPmUL3QONk9Q/ZeEkpwfjxpOAMEt4WvhuUuhJ5wFKSi4zZJeBoqdAGKrLMcg
GrqaZVhe6fq2Q6nK3JQYu1t/Q0XtroFMwoFqVrTu3NdUKz59C6xYOHbTtiKS5IK0Q71m6SDxtT4e
L17/h6IIMGR22jw6DVcg9Vf4WoVE9aWQb2tFUoDSAmoCQ8/aX6zChBKwwAIFxdWV+srjufTJLaf/
PJgvoweloArTnBlKtYQicI4mmsr4rI5tVWsakIoMoaB45yCPuIDtkmAODv2C8iTykOMzHKdKCfZi
djY00oEk8nR+2EZrp4gDsFFxaVctpCEqRgot42CZp3N3eZ+sb4GdsBIFWqy7XtD1v9WmS9UOIQkm
Jb3y0OQy88Oq+Gxa8LAnwsCQgbqQcRvifG/bpEQtmJxjNOej7dAjbBE4rBA+K/jh+Gx8ee/Wzm0C
WRh2u/hJqTq893W5r/juVFS33Axp/KjnSN26HBb+3fW9pMFOYCzCnTkeRCF5YGNv4NeUcCknr12F
NEkxlLNEYdgvWNqNUsPXnZPe3wTBE2XozYrFDbKuXCw0wgVwpP0FLPxwc8NjNiU816C2V7NmqxV8
QFewfUT46eyPMPhjkg4uxh15dZLVNKhpshLH5diNBTjNVhCCSJqYp62I+pNyDs9t3/tXjeTAX5o6
K2O3YEyTquqirTgbTu8LOWoaexyNmS9blqh+p9WxfuKaxohHYDDn8DdaJjYzEmLJjkMgQ3boFpAo
hzHZEmo6uqVQM7MEJcnEAuok/ohq/oMTdyo/9ky26dOikSjBi3bG1eLBbazUNT6E+icYX7vYT9ZJ
i81JOPvJKGVNq7lhQJERF5WARkmxk5djcPzq9lYH+W5D0jfi+T6pMhIZ1OtaRNf1elxe9emqKPp+
CZQYUHnlipVVv3R/Tc2NVGjSWP4C4AyQDGOT3SUJjg/VEXvvwrmWwU4HeMN40/QO51ozATvNcsoD
Ra4EoSLOZfYFY9m3QDJjRITXkS1IzSB5bb0GsUyoiP9dxydMx19WCr3k3om8tORozdRwMpvUTxN0
wz85IAwZ4YE+QyOjRvo1arF0EP/+xas7xReH0VPUXyXAP74Kbv6eX/qBp6/6ltcLSk18WCA3ED3k
qM1nws6+xZVPZigWUGTgJZD9Trk3OmIblZKO5am7fqE685mKUYHs30OpUzLu2nFXt/LBL8f/Lcp8
6hluo2OqbRzcqzJyocZVnyGTvybWMQ3q4GWPnao1enwqS08nM89zz2HV0AS05jnkCTe4m/ORnnNb
Qz3aQbf6EcPYh5o+yIeMb5NGxh7eKwejPpkdpzNuWstS96kFtk/U5lh98j6cMtoCaXLVpgXza9We
+3/mxwCfOOL5WctQ/OVWE5UWttIVUOYmODQ38+brQiTZzrgpF6+teLk7rYwnvtO/tMJ6H2NRNPSS
da/ENo4XeiNwEhO/Ey+/1EewZmkUrmrxMQMpP2CjA814Ewo22r9wkU00zUyI4pL1MGtwe/nBxIx4
zjE1wK4dzuR9d23vnRvaKiESCSWR+6IS6ysVycDWH4/XeyB0p8H0FZx2w01hlx6TchdYgmCoyboK
/AOyygADn2GwgptxxBRw7ZRHIJ85cxnZunylx5dtBW2uSfWEChdjdky7lUMvenpBCG9e4dwRBPM5
n1izMrtAD9lhcIgL0yu37b0aBKAZGNJlEGGUivi1P6yDHwHqj7rZAIkhzMq+AfbX3tEfQiIZcrmO
JcUWlErJFkTfp4VzT/2SuzEdsZKM0sWsMTZuJGALE83HcIu1QsYdTsbLch6iZjpet50W7msNwUTp
g0vjI9l5ZkrgbPOj+LeWF52GnDnPqQA/C0AJlncRhjNGV4mQSEMPh9h1wcUyccr4WUk/boWy5d4d
qFZ+14syNDqZyeTT+TtzE8U4fxhdO8p6o4Ew7HVX3EZAm4dVBmlS4fBrwHYoOoS/+UHOJSTHQS5S
s7iBCNI0IT9IBTg4kQLgyZWeTgG6G385F1l6eU9yqWYsKl3s9syth1q69F/hjrA+IMcPNzAvvKxH
XKepxW/89c9tvR9OWb8gltQcsuh0QBPbLnmo9crdsYD3mGfFwRbH39genR4hw4Be77od4sqxFyH7
DFvZcrPbcskOuZUx1LKx/QCrusvWbz2upgLoJg7kVun8pIPmOt5tSB7WSDBUweaq6hIHXNyagIGC
R2SVBxkxwHmaj/yLfvA0aFwq1qq1kGxEnfzhNNZwOY39ceUlAz8qkiuuBkyLNvFI4em3MTkyD7oF
/IQGImaRhdhziqymYRuXbCBrFgWrAlIw/bsZ52nQx7M/jxoBT64UT6SSyPo2rUhyEDXLyE2sbxzE
Y10xJ/WUxcO1FBjLK6uyha4AZMlf+afLdvqoBOKOhu8maDzGa+4txXnprik4O2AURwdqrqpXbAQ1
EjvKllMlVU8UpqR6r1j57ToRgxm+q1cWPrYgq1avwSGQfm66ljKIhjYnXaI5Y00t1VmZhyaLPb/Z
IO2ek5+1r1w9a4i3jsw7dIPgb15OH6RCp+RTw5ABu3AG68m15AFf8EJJdQ+54C1pohAu6Bf45TyG
dLi/mxHNPd9sfPEer5VhWUEi60AT8eCx0/aI8g6rEJmkQXFgtthIHD51O4qT3SLwzrgryqi7ywi2
Invz+N1TX6Q3Bm5jZ38dpLxupFZZPdyd8zaKzsuIBo/TgW4uSu7ZYMyaI7rDnR5q08RtKcqVGmYW
l7hYKNU7wGF8n7fEj2dtxwUuI5m9EQql+DCBzU8LCimITyVG4CPHwX/ZiiQyKpRxk5PN2Y6EOITp
2dJHFsKovfVFsi7r7aEdMxClFdTRYojaPgMzxB2uE3Lw1XjL+h4AQ3udjoVm47kmBZzWqUDfrYdT
uvD65CH8ovvy3ADKFOm8A2xvpOVqlxcYoaB65XC5SEq5g+Oio/lcjKKbagNsfRqUVxUiCEK64D6g
C5KDrZHiw4o7hyYw1VFtdD86zqa8Te9IkaDJtjoXxQFRbteXY9+rN/yTEKSe9q9hwSuBYw97ER3l
FiNWHH7Ni+khKlb3VHpNy6ZDhAZuNE5m/rvwMchn8HrwKi78jlDQrY4gXNwKOq+pbfRc4vXGns04
U04RC+gAdUSWbGB6IC+QiI6dCcBs3CEG/Wvm9n6P617V4VEVSAoa319/nMUyL2W1wli+bgylCllR
VIk4ZyQDie9nAqp1tTDQI4pQXABFmiJsfUKB/isma6ozAUdETuWlc5mTAeiiHIxA65F/GqWoJGFv
YTkxLBFkZ21AzQ5RqBwsW6+31UXcncH8UR30BgF2E0/yy60DZnT0rWkuWMhFY1I5q4R/GBUieSet
uRNjUxL6m7QPW1rKUl7J7iq/bLe0m+sjwKiu6uxDQWNNtusm8ZwxB6oIJ8g8CtNKEAqNrZ/b3QXR
ZBFewA5xve7iav5lIdD/HwMenuTaIl6tSqRlgZZK8qzQQnejduql37B4yCvb51O17XZUW2yI7n3i
i8hQE97Reug5lDrD7v4Ny1AJku1h3oS44HhwfJBH9hJiTHvcO1zKg73IYAvzk/OejU//tk8JPSf2
vgb/KvDmlP5fYV2RkCvf976dQv4j+KSeBTu1dc6vFT769puhUXBo6V0K1wASJSapJd7/xHalDIvg
gJVR1PFE7TMfkbRMVmnEB3Gn9OKLUwa4U1JtxerhG+W+Y3OyjAYri7Bni+7HWFRB3r4gK/D9UyH9
bNOYaPSrwoGH+2ZJq35pIa8zWx/2YD0qRsJqL6V52KRLXpduFk/AoWfbJYHBN5k8RVApYIoYEZBZ
zQULZfbs5VyANL2tYP+9/O1OXQSCt8z01RSzs8xMx2ocCyEJROH3RIJV6ZEEfQCTbOgA8lixB01h
Kj2YdI/CL68SdZVIyQjewuQkNbXlTyRE7UT/iZFeSmoEAcL0+BgA0BVyy6IQm7EI7ghOKwKBP3q+
K4qUE9bp+mFjB5ZGd8XpXCT2M6+psEuENVuiqlGE/8kkq8DSxuP6Bsu+CoG/72tRILeIsqiZgjK6
Okk08bWzPc3XFgdSX/bNyAAjcblHHGBDQcki1yR3MeAzX95UTXdMnMav1EMg7VY7WZr1BcLDvajf
qiPyPm4K0krQwIbKYa4GkaBR6sd2q/cFsDRYxi6s3WGSRbgc8dxcWV+Hh0Tjs7JrUDmleW7qO8Vl
4S5EX8vHUTIJGJozQsqrmCwb86v0CjGG4M9KWXY6/OziHjGSmbULL6nHRPDsYq2Yyh1RwCNS6QK0
U0l7wrsjm3hjuaPrUFMgutfQMYwVSWNvzM0/+oZ3vRa41P+XpiMAtmxnzLfXcPyjj9S72Wmnb/Z1
iHoWFKOJzKinF+QUlXGpGu7wTsZGTgPmIRtCggX6HOZ/71Zm1YI7updFU0PbN/lR3Uk2NdOuQrW5
C+3tDvOyIWkYcMm6KNNpbiBtdI0Pk3fJY36tOv7ctwTz2YZJ0mN2I9w0HIPwoltK1KeBjjPuZkD2
8vGZLGWNOrfmpvyne85t9I+B50SRLvg22ujw5jegu6GrDMv3TP3siWFh5jstuJ9hx8ceiRTBxjVf
CgP3DRwilhHBwsgS6qMn1cDr2nx80mPXM87c+iXFRGumoUmcGS1rAQ1MeTJrbF3yj6lv30cfbNZw
BibUZDWwqeC0+JV7XLkGKRc8gyrikckdST13pn1xIBfq/not3HyXrh6k6dODr05ogAlHmZmXSTaw
DU0IRtBfp3Q4kNvXKrdSHG6YqY6RT+LPivPKm4DIWqmxdd+gdcfI14s70sK7C3E+0njyAS8GEBZD
4OYdxMIyB5Qpf2zOQuZgniwKJd5H0t/FU9Y6myAAt16JV+UyOx6xYch19LyQQIS3yoW+ycG7E8kX
rbImWtNL9o707iSnZT3QipGPra5XWuokI72wd4u+xv3XOhN3SlyOC+kamouaKO8MuwGrZrZErabZ
7ucN8SwsNAWJ7gsAXslSGbHBLMlYhlAHtvZMW65YSFW90f+5MxF5PEGGa2Xwzs9oeNp9JwELF5JO
UPgiugZVKn40AvB0qM/VCk1EKLKhgBQTtopOEopWMmpyGnzHX37Dy+xHpHzPytlz4G1KOMaWUsak
oUt5JgEgyuJAmS7CY4UiyOl4bc3W8mMImvhC1FzGFt5oCqwHQYZ42IlnrDhJY+Lvkj5B545fxQ9J
j6t55GB1SNq7L7KfmOdToCBhPvtgyX+89h3rvOOD3mjO2jXQOTv+Bq3h02Blsgzyjw9oIbGSCDq2
rwd5lCr/ACmDX6Vojyj0Sgx63Y3S6Dd97KjSynaqCr/TvXdPcgy1z0QDTXTLGQajI3eBdfPf6LnO
aJzONFVlzKlEr/fdQlwil0qQW4MTIdC5b6AkT7DRtHzYFzWV7Ywj2wV1iTrr1rDdUfaX62dAgj7l
dQ/19StS9QLeEUruJMvlDrF0hNz3pOdACOxTIXVUpY43cBMm2qbBirZibLwK7zdoijTwIGZccr2F
OKY1ZvMKiIySdqIeVj4StqVMHOJqZJYvjvluGqgVtprpWQ9niTYp59MAiq1JgkiOtEymbXJGLlIy
BC3MIEFA1/hfHCSheIOZ/i3qI5SYMlqpqYOYx05GaFnhLrAh5lYsknQCi3bucRsrSdN4FEdwL5yk
TpUlW0HIE44DSv+537aBbLFA8LI3l+zTtWCv43yKFzBkixYAYKZ7naoDFY+Vw35q0t5W/L0h3yjr
h11WcOo8VT6DUxqBKjfXlXDpCpjy89XXKr8cW/DSd9aKl16MV9oGFeM7XX5iR+KF1wKYwrtAVpnL
W8jhuVZls/9zL4HCAZeCBdXAwNIrW7BoYYe1iJfquCAFtVrsZJ3WI4si8x4mPrXirYL/yo/XrqTK
G9lTKivurSn1M53T0WqS75QGnFj7yoEXZ2g1w582Qv/DOk+sKDpCFoizkjWYzrv38v2COmabLdVw
UDn1a+CIHrSWXjijJOyhu56xckoq17IL39qikOx+qB3lUu8ztOkNBuZegObXtQkbdHAO36UiMHnr
jOVfKKC/H668440zWUm04Yt8hS4J+JGgtWGgFC7mKtxNk0PRFgbkX3R1bl867lY/3KTx4pHGQ25p
Oy35SVezE+eTvloUK7nNLG5XPz/xwgxjobGUARnxATRKmue0F2mHRd+i0h72ECDCFOoPr8m+GcTn
8b2NPtXQpqroZpHctopeRVRfyOamn89ciW0Vh3IsJmRpdBb62uW9F9Ynoxm3Eaei2r4qF/qBi81c
VyjtNeTgmpMVNA+kMipRH84JkUGNHqmgbLKLzfxIAuFTITW4HwFlds50srf+Fb6cdQ+1AUZMMwLK
fFSuKryXi6nRa3zPy8FUmkfm/4e1TQ43ILlujzubEHquXIqwf47cTfwDNqMvVrsVQDGSqp3oLPaX
fOe4q0naoMAyAxqwuDW++LmTkwKIZPAUiX7hmvr1d9Q/Qw/O4vc54hUxyZ592SGZ+LR4nmGV0nN/
IlgXas/6C4hl+yFV99po4croEbUNpxKIM5OEZ+prR6Vd0wUjW3XPrNfSvu7plyq5y2rLSvFEl7lb
LsRMtVj96paRs0cSIViUb6hJ+P+rttoXq8v7e7z2cocWYuaow7JmgDnZ/PWFOwXoLFczIbXH+RNT
TNKUExuEtshl99KYccY8wyWtpHXkfAl0uwzBkwPvZaJEpVBShmn9MKQQ4kwhmZIDxg8xFNraY1f5
Go3q3LswGGPENr3O80ev/xZpavw8y+95piOJC7sfR+iaj3RxQKakLiN4s8kVzQoWujfE2dSkY528
MM5ROyx35mPbzdn3YD33uZoBuHUJSVeyW8LNXi9cCtzXSwoJBE70qzKHnYVu1RXQPkb8qXWZf/fj
cL39Da4CMZvpuALX8CBNu34XLZAKPBfhKgcrW7tBXv3z3ZP4VN/0Rbk7mEu+mzVHHDZ0/KU2rULq
vQAsqRRfgtULZHf2aKe+7abp8lMNeabWp2wOEmr6z5N5lq1RZyOnI/zNczUSmD4dXQY8P2+BaTKh
xduX/z/XdWYCwqdoICGHV/qHculkQD1HD3hLoaO4u0q8AuSC3T0pS9dReLa2Q9NBEY1Mxxdfv/rN
XS6L904Y9Fs47cNyDIjvrAyGhJbVfBgVmGSUq1S15pA12PO4gYApsh50GNpmt98VwfS/no1nQHWf
fs1AW/TCutRHDpEA94kozgJbSxVe06sM/PsMkY++bIG21xBnnWhaz1GBcfdKITssVdj5gsF+/6ib
GyfVO1h3FTBzDHgcrWml9hKpQXzFB4MQvL1tTPHp6wZYWg+MSm38QzDSJ55vfkq0zpc8jv8sKl8f
iW1TgxkOnnrHTF180ATtZ/3P10WL2t3iMfrQzexJl9zB/PrZcfLl4SogHDTNP6ANwzA59l9DSFS7
0yIeE0HPDgJm2KktcbK0aSyfKLYXodTWwIjLRIus5MpkS2rr/jr5ggo0021ZCJbR3xnsHcjlezZ4
ng08AuYMf2iiRDwh2AuDvdbj7aviqMB8JDuKnU5W51bD6WCpCyuE+E3/FZwSsdvehn+szoq3Ysfz
JQg0Wy4eaRnR8uYnDtrq+ecXHkqRNAb2napWv4JFlMvE+MeDK8ZnpRwz7L3L87nLKigIhEFvj8Ly
x8S54EDU3Dq2qz2ug5TZ2Q2NS9nV5Q1TElk98lbGq9fWpOm/C3ONpaAj2k0vgdqZ9iGomsIU5aua
wf2BoiktPX2kCVKn0XgQHFWFli61AZr6B86BNv1Pu8ewXksGRd+PKCSNzmffgA8qZe6YwJ09RFwh
YQEPjvKVjtqlMz1BQYfKcO20ZSuc4FpyQdyTtNMtF3dp3sCFjFMeyubJQk3LKQbZzRrLEnI2hZLL
FqZ/uju3kureLxtv35zDqM/tCTlCBOmavsnXDwTWCxh8UdjX48U201YeZUIIPEMZWvNhku7jlo+f
fDczGma2RA7Ss+NzghCyNI5X/5HvFIDSsRIrhMGy1m4qTljexoZ3vFAmC3sinJNdck84CT5n8Zfx
IdrderoebML4643W4sR3qOJNy+ulI2AklxFvYo4kupWD2ldokF7nMRcurimWDuIc+Y1xPSUMdWAn
qxUA5R7oTIogRJ9rt/1EC4G+rcyzBrc4a5n2azyAXufg+3yqZNFCPfGahleZDtsBWt+k+PEn4ZMp
6tkeJdbeKQshWTDYrdHynySTRrQih2hjRjU4WC8be2vqUh3A0XmVT3hChJo6Qq7kAmf5hl16TJAd
hkihKbzR7tcu8YDdCbryk0XxWJBqllses2JzgtF0A+zCpxLLFPRAgqgW/fGQ2ovLoKf5sqEExwGs
KS5FLNFCPYaKCU7/W79ao7Zk3Zd3mCSq0N3gk4GxpnST1/kyyLKa6A5DFwdDxzj1hEGZoEEU8pjF
AWGFPk+68zYAryTZUu4x87Tf7zGd6eNhaUCwQbfNpIqbZCAcAlocm8leRABZjFeEuUcubCsxiGi2
bcsn7rb+9EOKxcNhxvxm75AKn3QGzCVawn0fQ9YRFGwF0Y5iyu/uqoWJQyXxm1pDEB7L7jdLYJgF
dtHPUc/0vUvESE6OmQqyg+tovi0TLZ1dMs0VAdc3DottGc3sYokVUasQU6TX2QRl8rWNPZsEHAR4
iaMfvGyyXTPP4gQiM+pPjLithQOXg/uL7qI47DsCa4+Oo2gO69scs36ujIkXSb0Ru2AEFH4vggue
Ja8cZ2Hnhid6cF1yIEE8dG9QODNk7easZvscOUfGbF7QNzeRF1/Sdz2eb6CByiXCxZbkao9TvgrL
x5jv6btWOa4V1BIyZI1iLKhmMrAdbBD5QLqaQ8/IqbVlAYFNRIDqYq6lbaGcF7d+joh2vIyVrFXK
pWFe0BYgHUNxbFTwi+rcPlLn9DPfCGqeyGY3DhMgFt5rjRRQ4NXFpPb/Ar9kiaOI6dXEz/FvBGxU
FHpB9p+FfKMgLZanjkAmloAWCVvV3JwfxwdFuDwLCNRVaFKdC68yUvMo1IbEYgEd6NGjDz1T7BTP
2YpR7nrjD6cwWdCstFQeO+1X2yr/r3Ds/F4s1TtMe4WLdOo7xpB3pVbewel+uofjvXXnQztqTwm3
Vxf51MPpRrqbaDhgN/K+MhUqkeJZRT55tDml52u8pXw1xdNO0X7ipGFd0PLBW5ERC6qNgz++kM5d
Ra4Yw3FF0lu7MwYMIfMlC4xgJ2Z4fRmRirRV+3q0DTGWHRw3o/nGjJUu3XqEDcytV+XQpW9f8GM2
ToVD6X8wB363SQtCH0emgwQChUmEN9YEF0Ji8nbM7l8xrNjuzkK6mNOUJOlwQcbGv54H81rNevTt
f4iVKkPjL6Zm6sgq7Fkd7QBr3bUUHHRFUHU5L2eCp2fliRViHkh/5uQRQbzx0oR21W+z3XUWocwm
WqjZ7/nHrFK00GULBTcUzvOJZC5jYBvO3NTQQPyUrArDydq/Uce6bzt9lHmFSEQPyU5qSFJAoT9r
VKRdtMZe7SI/PFC64WMmGfWy2fThj/5KoJmarKer49ahbG3OVGiNuCirq6qOvRcpJw8yGru8XO9x
JrWWXUaLBB+XORNR5D7H7XrnOL3Lkc14jwg7YHsKCF5jvef3vpIsalyd9WkXI//sOMfkD5T9CFVe
s2N3lV6RjTTn5zQC0JzqZWALvlWUnjASUabtQW63X6FNP7S8uJL9dJ+eg7ladv7F1l8TdEjKn79Y
xVsjCBLfJ3TNZgDWUOLIm+tZDi6SiqTJ1xJrgDeckHTPi2bFN+cvupwUZy+XMKROcZANhy5Msc4W
btsRm2pRETr/W9Zll7+D9X20T0sIkSTY6PGRJf6Zumu2vFcmtUSdpfOjH+zcjrZlMhwl7kLa3LQo
8tGk73oxBuxMPLftvtpv3R4s1qyCid4au0G48ed+9tDZdnZBIaA8mlbyhO0xjs3f6U/rgGiWulCz
oS5qp9+b4dc8wety3aZ9cC72HWegyRjN87JUQ3XtWglSaEzw7q88HmgvHDrOzBeVcUOYqWOhv/Qf
xHvsy3H/rI2sWld/2R3BZ5tr4F5JdYQdM8DaeKC1IjvHUQEgbzhiqX7vh0zoJD2YTe7Rs3w8IvbX
Vyb319XH/mhhWTktSuoWH65jD2SL+es0oKwA03fyw43Gff1PYitoYjIZQt9bJPqsAFSdZ6pmIqo8
OuprOe7EVSTrijv9mTMTsa6z0BoU8/JuFQtc//rmGqgZn/my+iagm58RdAE8yPVDhk9xSqoVFlIf
eacrxEe4LYH7OWnkrRnqAMTIOoNa2WMtFbbRjvkAdtp1T94B/bHuUuWwejIyOUzhODt4eSgDkwBi
Jdvhks1+yIZYksoKsm54jp7L48p4MEDHjCXaSUNwPhKj7mt3iM7IEoFoCUiCxUjoFU+W7L3O36yi
15+DniNO7uUNR85U49Bnn4nH55QZ+g1M7P854BQEZlYMy/qtid4MIWgS2FT4iiBnO+qZm60VpWkM
uGZQwM3zyuLmRs1891chy7ThZBtZ0WNCBeAkBytnzdhFcLT39y3L1Uf/i1606HSAm08Qv66dJJQl
v1l7ulC/wjA2LcZnFD61WdX89PoZ0T3ry/zSLFCXyJ5NQNXNlF8Sl625OkKpD7kqL1VjhM7uUEcq
1AlnTHTIJKMJIhLQjWYH4erM49ibE3rZ9ONKJDE1baMVY9o1i8tnJ1EBk1l5hTOSrSYUz4UNtX/c
Xg7ar1LxyBmS9t37Spi46bMhAfVwD2eFjme/wg/im0JyMo/F03hRBQ8cdgS/L4b2h3U7iPe/diBy
lXS7l5uAQfuq0bPLzsQKDhXTsIgZJm/Jx1DwvAj1D+gDQLrmEVGY5P9Ob1Jix//u7Z3Po6lIYgeq
oGuBBq3GaSCNaKt6yB5Rp3FeepkUtLGr3p+6Q3dIOpmOCkqBsXnqSWUdhRF7qCapBGsV3EJNtq4j
1qwjB3xuA7oLe97SNwyB5ntkifTQF15Waw/ghAAXMhVHSymJF7gcLTjghjrKurI4gs9uuetncGhI
ToIC3Rv6YgR9LF/6j5iduwGcdIa78+KEL5p4QiVKsLQg5RgRRx1huAZKY2S8agirSBOw66MBXxLi
L1TytmP8BWEarEnvMIodmwDmVYS5HS1popURkqxfxn+wcZQ5hriwZmlOP3Up+d9QBs7lNUZqqMRx
O4Hc4HF4OwBvB8b2Gyr8o3WIDmTgTaT/a1ZqlhBasJAteWKa+UM3rWdOVvxK6kVrpwVd3sgiGpsJ
2pHHWynOTiGCbF8C8fzFDDaB2VYXTEi3qdyYrlFmtIpA8iARFb/K3QQFz0aBKihxW/TFqGCE3Oq5
1Wx0SZ+v3A9NIlcAbS/uqCZISQmT6BM2UOOYHMjMDBPNXv9P+lNKsg8qKsrB+T9FNZyFtmlj6VR7
mGR6xhVvmfk2oDRNSiUBaT7n3Rmvf/Xapn6c0RZBu88sPPLsfQIAzCRRIDhFqMzlmGE/QIHRpNvX
b/ttqSzrIbthRt9k0aVBHfdx6p1DKIfORm3DlxSuJBvp7MayvNc5TyalbDQPnNW8npdMtF5sEl8t
6tkfwub86ManKT3UUGpve1/C6SP7P4jpLmQhIxo4HfjMIizMxbCUXSTE5x+1l96XPKUdzj+pXOjp
wjMU/Hpt3mcBflzg+2SFfulbrgaiHYV2yrd2N143aSA7X0Jt3jCio3HpJOy/oiWGl+EOdvKO8wmm
D/BdnEW1ZDvK0EHa7kGvFU9bujK9nRRp+vdIUwg0aiVWi/1l3tibkTAq/l4GHMU7RGqTBz18FAji
z7KguSvAzFYgBTsLV1iBK8d9jwnOWX7lL9aE2An3gxGqky5LjAmomfG/W33xQtoZpU9lcHV0ek+s
WD/cQJytbVz0xg4YyyRLT0yAUw3RKYizsTYfjGoaJQfJEiamz5sjpk/cY/FW3kEEMiafnuQ+Hd2J
U6qxKRfwFRGuuRBGx5upJYc4IjRwzXyKiUXE6XVafJ2f3RAQWD0a9ipwcIJHUSK/J9rA/ei//5v5
J8rD0DlJQYpM7U1wBR9ey1uF4/GozqNwBGAmznB6FwB34BK9LJ0bgLHIfc3dHEW56YEfiL9LlksQ
cW67J7Ls8PfWGKRUgBp/hHeLu8pJBEXmXstK0jFNIQPzysWQf0FC4i9ZRln0Te2DQ48z1CBrk3YV
aYLHSgOsOWle/A1dOd1DRLaQCfeiCKidspbgP0VTvcxqF+S2giP0VMDMpMhIUTQRf6AQAZSj0xCC
cN3kecZVpO0Y+UW9ZQRCCvvGABEbsPsbRhbq4J3TXYtnJ7lhcK4gMhkMsY0xdvuDqHnO/7k9AmJ0
KO3tcgFDx18MuOTE8+OaNdEhREc0XXLGJomHgEfqcYv7HX7jS0QQ3ZQcXY63arjpyLibDxtMZJQB
+9Rau80UYzqJLUKbaDuxPQZylNClKXuf/pB5oDgQwwZVP4WK7o8/cHqyOGttb6yI6MwR44amrRKq
reLQtewoZYPNlOw0ABHGR5DrrNsiOyIG1QTUWtLMTvkIl2QDzU2ExaaRdTreiMvSIGmpu/ICKcIT
A3lFOS0mXac9KQ1sEWa3hbyGz4OPvRwPV4BnUuJ7VGTD9Zu0v5O3YbscafYq9agAV2KExJl7LcIu
es7kDQtD6GAwdsuUcT944htY8/DCbaXuadwU+stGGEMAWsY79djpoprHSzQGTlQkMbN9TAB1J8T5
oK8D8PbUmGn/XkyXlpBDH4+P/+HJyrYkQF+heKqptFo8uMpsB+lq04R42y6hqQmqZMepyJsLy5Vj
/o0BvUdsffHUC65ZtsZnVV5elJsPYt685Dn/9KT1hy4H7QEK/Vn69ObKFlpXyb6wxMz8/CGWheJp
gNgRUsgpO1wUaz4ijaeLRlCe0/v8pNM/3Rv31lfov72lZjqOTo1RwHmNF5+b7xcNxVH/VoVcxZpJ
D3VjREzwHSaDPYs98s/ME9I5HMYD6pqfjCJ/4lL/TdTDm2617izCZPN+84KkYUnfTOZZ/idEXp9R
0gQhadLRfGEFxM1xZCnakGZaxtwo41KebfsHWXRxv9wwP1EPUPLSAiFc6d+1gTUgCc0NCIU99gwD
Va4HqMz/bVwikTr0L3IPkJMOCJVESkbbTDopE1NOUPzywIIFUuj48N4Jrdw2AGJSYwCiC891M7xj
EqwfF5ZiUvg+riRRFjgICEcyOSW2UAIfRb3CAGCEfNp2UOeWtjw0HnA2dN0yMgaQTzOAN5Y1mnDw
aFvsLoryrA4uTzIzYtoCn5WfSfv6QixeAjiNTZ6lzc43SJDRdQxuaAjPEVtFZGu14gzib9LyLYkb
ZsILH+5kxjSKPPvwZnV1dlOR7pBeifQ7Ur2BqWwBP4tzc5+zb1gwOveDGAODiU4t1mdPD6yg1oP+
HQaljALs5JouFdRDwa8oW4EVDHCoNPXwj6MuQ1GzUYAcx9rStgjT3wHI6pf+8s8edj+umOJimTX3
fzsoMDGP04QKaPCiMpvvvyAbVC6Ns8RT1gjIKPSYGo06yvwc6bXqZHIbpaVKrmypdJ3KSf6mO9ZP
dtKSnj2NNrrpYWVp/HD6UVU0l72bvqXRI85zQv9pxxgutypGyBBNnpzoCWEb3MRRKhIYB486b3Gm
Ptp9uAy38A5KV6Y3LmqSqkDZ55S8ju3b3fc3qYIZVNWZ50bBE5w5znurV5mxpxUhSkfvPH3ridgd
Fkexh5gg8VkcFoZuhc9GQatKFm3tP9tczGGA4ZhxGwrTZAzSdW1z+WOCe5/4fRY/Etyt6FBdy0Ug
Nmoq+p1fQPcyxhuuGw7UpwWOC3MJdkinoYMdlkk2Q90j8UZ9+LG/IhtWq5qvZn0B1+AWEFvWPeH7
20xx6ZbzbQMzCDG79DiUCGks2IylnCvLQirlFzNkO6HCFI4Kq4aIj1JIh9xrmPe7Jq7J93IJDAWu
d/ZWWUo2N6GEe6qmQcB59ELKmEArzHQOwCNiqywod+P8HGi3jOLkNY9bbQQH/zMyN3e3tXmdKXgx
+cQTIhCLbhkpt2yCE4jIVK6JFoADOyESk6QGcOuCtQwq2wtAF8LXeD5VWEHkwNswSy23kVVIqoS5
L63fUx3+SjmX33pFkVlLv+3R0v6QiXO2qz4yxZpIibsxyMDUsfZqwxgPz0R3WN+XtpMvErjlnLKM
TECVROrIVWP8WFiKisw1kb4ajUzcQ4cksfdGJMk1vZY0CG9cXpoUe59r7v3TEIHXV0JT4LkaZuPM
2t8JzR3Go2aHxawz1d7rFa67QfBxSHGHoUxIBBRflXfm9dvd/OFi3AImcm2ld8sMfWJTbTDBqi33
esgaFl9lpURtY7jjPk7oiuzULNy0BlRfxPiwrGpR8buWq9ItCHgaxz/t95Ldek5npLDa7khRYMx3
idMBuiT7paYwko7wlSGHp/iedKGo85oAsjjB8TJF1SyH4uHD/5AkEPPhkqWMYItYFVIXpjxmVr5Y
1NkULDMhxd2V2X/clTbKt/mvxrqdOOJFfy1mpWvx/ozwy1AqpxnE37QYsxq294fhG6Udgm997KwS
7ogAKV/FDNyWUygTW/olU/+PD9P3oLiH5E83Po3eVW7fXcizZGh2SnB74t7xZM/8Q91i4wAsVeTj
DWStRcMMHI2d3M5A0kknSDCENt2SB3chFRdPov+16vF688M6CIOApPUTNALT6UIW6BoPX7r48kw0
YavyfiOC0BLzj9mNBH9IeErC1SFTpdGW0IMj9YDGsnpDlsnU8E+7tEM3kfzkEKAyDP/xjFRY3xnF
iwUE+QmlS5DM54ueUusNmwfOYeBfDYG2KrYLVguUDar4rjChU+ICWsipeyuiR2LhLYVBBRRRb0IK
Frav8YpisYJ99loS0tQwNIxNOBQsP/bT2mEP4pbMtHpu/fqcAucrHfdfr0Myz/fLvYByN/wYXeZg
XWOLBd4mmsd+tgDLzxuP5AwezWiuaEJ2fzk2fF7lHmThjRsFZu2fg8pHGFkSS2lwfRUc1mcbh8zP
++RpbvhE3945OjxdNY7pwGcIPoB80nYjkd+njJmsjhzZSpMAVSVbvaGPicMfJhphm63HfIO63+nW
UcBw/D+tD8gaYogZ53tx/DDdJ0LtS80vF+Yw1uAnreBPpDRsOj73qpLiq8MTZLImCidR2ShXEuTL
lL/prWWsJOLie4bTApAz45p5M3lcFOnZPIHZOvooZyTnxEAsTIDjG6wrqUfdzEnM03tyu8UgSwfD
2T9Y+VIjZfgsRbvwEfH28snlRJbfgJ18I3PpYQ07WI7jUiA2M2eZo1aiNXb0dE4lEWtUyEnjydTn
f7BNvLB2ePpDy8grZ0ihGvGycQ9qPu6sbisPh4G2tzc0qfGM8ZciuljfnSDSSrOiGhUSs12dhrp6
B1cnfPupNzHjdb07eDlD5haYPR4pczz1A0TjdzmDoq/1lyVqr8mPPUdJ3PvrT18oK5OUbIqbR7YE
qi0W8FWaYqfcLwDcelRThaMPYr9WHmetE/1X6H4JWBP6FVG1fe7cI/CjOkp1IOq55l+Wi0+ULhMk
d5zuZtirzMtYwMlos84vrV9TCUCn9J5vv6Zhh7pQbMZM2WhQTx77VK5jVeHm1f7j5IfvUEcOk/9m
4ipmwcmrrlIOyKPRUHSHe9G1aX3kCaOLKLuocjWQW/H5coPXjG0xFGBxmMMwUWB7MxMt8Uqz887G
MDs6NlDlIwb2FZPF7HhcHliYRfrWRk0gJd7/JwpcA2iB12UyDN4Tx1hu3Ji60krG0gv+08DMhdZu
JsDT+5dx9BH83tSoYrRNxmrsCCJstoX3jBxxasibFZRuR2mKGclDHevdSz17BkXcDkfMjO2kBk+R
GblLM1JnoWxwruvaKAHvs/CTqow4AROM5BT0BU66ga+guH/Pe6dBGTDnKmTreEPbySdG8C5+LRVF
t66haUEMnRH95t3K8/5aUv4dtPVtQ8vJQnJ6mvnTnixIDd02ERvERTmeJs5l5yXu+fl6Mz/0Lm3r
qm66ccWhudSaYIj/gtirrdrPnoNMMlMlSXbH+2WfP5R3P9txhgj3RXhMaxkGATksd7s64rvUj+e1
9LE8m2IuR6s8qfiQbzWyrYksOdLlphdq3i+Fc4RwpbuKN20BVLfrE99XCCVY+smYUZB0x1AtIQyT
BoveXZUaCdrC6s9OwEGzZtnGpuDJ3w9rllGYmzGfKZhnQSHCdi431rVpImlmP0N4KuyWMH8InQjj
6PLaJKf34zBqw1fToYbjIDdMSN18uJvxW2Da0vh0wJtNvdFeKMShe4nFWE0U7GkfS0xfdNxiCndJ
vpfB1wEbsNPeWB0js339EeXpp/F8KK0NRPlKrlFD5AASXUTbWKx20N2Pco6+ljVkQK/59k/W9PW+
bUK5481VkLDUFqSHOS/+D26Jz74uyd0CHnv51VG078D1svBJebTHLEN3pt6dLZrirO2ZiCio+fjn
vxXbuDZJ7bUnceH4iXhfS2v1UvtQgDMuVf1mlXXBBaX/HB2B2b4+sSUx8uXCrXK+Q0U4SxXcPDb7
H4TS6W4FQ0dGWvXcCdofScCImhtddI28YFO6fdJm+/L/g3YaBMTcYbf/hseqaxwP9ido4nqD6Bfo
+Qs9aVCDURvMDy2gqpid3tLajGzj87G5OBZ6jjhtHeX8sT/2HfgqaWL4BGQJz99S1N1GcQhC+zVT
PyeEvydvD8vIg67/LxZ1EgOP9TLa4tIjPkkNOzbJJY/OF8Mwgt0zbrLp28Pk0ng0yXYaOjLyNFTp
OlvWoM8DcEwNEmGsTfx6C1PZMuxXM2cRm43TR+LON9YDUXMGojnkZEAM34GQ3MI3BJSyQM20FjZw
4KH2tz8M9R94m6Jnpj30EQhDSreV5YnEUdgrpYnvd+qBACkyh36qyc8MagR5KCnzJVfdH6eVA+VL
oQQ8yuKoy8Cf1xYdFDOei+sqEEDFvABD9GQoaxgWdlmUa1T3Xj0nSq+mmKafsfSIGk3Hww7FN4j4
0kg9U8AVTjDz61M+AzUWiV9hPfn7dNQNXM6OxXMCwzy4wIrg4tNdQJPYLyVMObIJrC+8O/qaiWuj
To0rimEtr0EiEsr0qy389bVArLw7/QB+YGj1NNaL7WxZWUD74kye/nAPBXIQ21Bb+Q7Uaz5Z29mA
aXy5Z+YL+IbhKPd54qGlVkL6/E+aackebsGFLcI6Cpx2f6k+gJ+gNHF6pypKPdJBODjxpHjgrX2O
7kbG/1oP58FWYmWUvNR4yxYvuk5tNE4FfpUxPLsd6TPoJJq+waxLaEu/G1qp8+Ml9Jjc37wFgheN
RtlRNFSYcM3pAFjRbx/uFhUFIrDJGyDneOJw+scWvzOdpxdecXspukASzPvaTOPaqemXlCc3l5jU
8agMBhpGV4PA/Qt9Ft7kDTEPe+nEYIVYA+KDSvZBpFVoo9alY6AxiNmDUTHuMeXw9WPIlu//7eKX
bLvihOhNJ279ZtvU2GM9YPPG3LdfeM3McTtixUZLCgb5awl9b0VdOh4mhm7SRf1eKVsjROcbNLqD
yYI8KcFPgM42cDixp5kTpOc3USVMZc5Fp2pQ6QXximIxn1pXdldTfQ8W1+mm+RNrmJt205LCTwlf
wdByXshY4Q9WZT2sAvHQh1R9PSXXoUyJepMsRa9xB3fCwH1TCW+E9TsEwye16kHl7oDQ3sSN2GD7
+WxnGTSQmd9LlZCmTCkiXvuZCKYjbdq0h2tP6W1yYFWkTyTHPMcqzi0281Qb7q24drfR9g/mX3Fi
pUz7H/HN/CLwi/zvinyx72uUsQPuhm7K24bioK0VVEbh6YmNVo64O5hTdSPoRl236UTWJcQVqIU5
yD0TUO+nq+eApy60sZBW88A0IcvyeQGNhSaJ5hpbQDQYaSRH7E0EdveQwS1XVtZZgY96Fa6mo4iy
8towthWl9slpHEQwLb5+NOJ07N2CefCIXytK2jfNR/Z4sdhSRbmiMcyaQHU5mXtfk3QscSmFHOAG
KD/FiZy08JhmFMNnDCOeCZ7rTwlTPNsIDh06cVMaDNjHiVl6KKjZuYIcE0wyfAoxfdtDC4JZRf/n
kXgaTkxV5bO+q3026v074hTh0hKxMANhUpba6D83Hybw0jt6tDuYjipiqkvMV4ptjWKRBx8gaB9L
EiqrM0h94PHnVXxWNApnbQCRw1OpztyxMWU5Ygvff7stwaSEQ8cBaoN2VqoQrX24FIGt7ur0oTDJ
U4POEfxBRKggZbGOSZIOYBF9UDQcy+aMplp2YSk8T3NtKkUtZ4ACIkc+lJ3JlKSTMfocMIcxwLa7
qSSS/S5W7FUmkg/28axJOuCqalTCY88Bd4ApHUGXjR6yY6hVFt7YKxsEsrwp+648zKZ0T/WOeLXr
nivly3lb4YgH2Z/fJjbv0qloToURPPK8UyRgN0g+GvuznQxJ2qFU9vfb9lZghp/arrbItd1WSUq2
6BrUb/WnxRZAH1s/QPG7up6nkAUKQkrc6aEycE4j5wL+dspnGPrTP1c5MoSdes4ZbYR3798SJpRj
8t0xskmG8COZhQ9SDUVgRxXJRSMjT/BPHws1O9YZ/oJj0FGwP1JAAa7WhXy0HpIicJCdlzah/tpm
rB8EDDqPA95nqyoMfDaqF1iOJgO6kJmbcRkNAeQ/dgk0j1foCr80ZK0+dZvK/qsaBUyJ68tf2uJ8
rM8aDolwGRhzrZ126F9rXalYZ65NlI57k2KZ2lZKRypEEYszDSsX86yTXhmBf4CvNTwiBUG9TF7j
RoC5rNa4nFcK8CnMmfy7nYrJLJ4Q4IKrPtpFeorwxoT21Re0aAnQjwRI6P4FTwG0EegXTs/Wj2pq
JWy1QvV6JUChA3X0V5uQGuQRicT+z9K1YLJe4+g6YOJjjtt+d3wRXO1MvHc/Jtpys5WGG8H3Z6x8
RfWyd93jOQfmnerW+BdTtE1KXd/VRstI9U1cfTYIFmW6nUuslPnLdqOVyPCeUUfzcPk5DQtLRrZ/
Jim+57wWj11IVK68QFUBvx1Qg+vdPMbTLaBZdT1XXAmt685KUJxSR43YGIyYB3ODb+CdBIepfbba
B5CTubp+Qmfl+pg+06hFeT6luYWEU/XSlABbAKwhX0Qf72EyPN5KtZdPZiAAAt/AFoxipPCeRTn0
Krj/Ui2Kb00CsrCkzicvtFAD/Z5J7fXrSOmLc2lPOWT7hqdeRMB0KHJz2IGLLe1qP6xfQCYlBFRK
DnmTnWTv5OIgkm1dOQ/FJTgao7hTpexQaZvyP3iqgOn3RKZk2zXr2QhNZYp3UbWFQi5FGVrTlIRx
XeX/ebn/Oo5hp7HBrbG6zjSDF1vvLEbAE8aXT/bie//5drm/3OC5TGty+1W4mHLTDRb+rhc8TpwL
lh2H6N7zaIjvNpc+TKBtCxWGXWuNJGvHbkVmzW2S+0TqW51iADSwRgUf66PATzo5D57ocwcnZ018
hCUr71PP1aOVjYVDuw8OVIEX6/Jgfkf0Rt/3+QqPjXtEpfuab77aKL5ywsjYSPv425s+9zcDeDhd
2/rfXsQl6v0gmzPGlI2/2emxHkRTFWkCUyYSxWCfYYzC13Qxqe1pwZEJ20NOeN6IxWo4ByLl1nTt
Eir2j5XAH+9ZZ0Mawb9SDquiF3kG0jMzkDRgKExutxsWt+fjPqnAhppW8bsuGJEnZXMiuw154/mg
X+4VRUMKAnqmMIU8o8B+GKTiyl34iJTv0ABHmY0QJ5kCM3eq4MXfhuocwi/2KJHbhmZz7o4qx+Dx
ST9mV69Ge5InIgXFOhZVxNtnWXxL9AoBF/wPfPI6L602nairEi4M1iP+ohB4EVAEbXCqvp8VzOM+
kunnSx0DU/xReADqd7O1b9lE1crFbyUFU7xf5mcUIF9bMTs7Qz6ir3HP5ryKF0HmiN1N1WWtRLeW
W5BPUvHOpalrYAB29Ez/k8dgOxzumnUfUfRffq7oMJbEMIJ0OaZDaK3LC8+Cpr3doHn/B+i/RbMa
9ca/3ayuCB03jZkEY4tZFOip8oaiz/YeLzLG6+izSvsVcBIP1uEIw432OdHDK7RjA0LiCqp0ouy2
1IV+x2wfZypKyMzk1p1Bl56cZ6sTwdSAsyQ0Zk5uls7fNbg2e5XY2IQ4oWaTH5BPqBROefW7ipMq
xNHIDo+klxHVUOjHbHdd7IrdJOsAI1MXISKvl1xn8V2yFOGpaIqCIJ41HuOySHquZg8mQrpjeYog
KxbN7pjsqqScyUWcbQGIib4sc+ICDKbIVKklxgy7PiUQUZjgnWwfGA40cxsE1dlaeRXZzJq7OAhC
FY9j28fxTu0xSuNhBFyymaiBX4OlvKgs4Sr8sbe1Lu18ZlK5XTp1dQVNS3kqbJdPqvOBUKsE1KGo
PcKaA+UI/Gb9Rkc/51d1Q2Uyet1s0CR8b8TT3cE4s2G/3rVtBWEazSjHhSVD6i9Y4Za+1ZEvD/VY
r8aGzIrCURIGSwf2/SHUM34rudNrlQbKfJcTUTKnVHxgeHy92YcnHv+f+2crKREDTi0qbV9OyKJz
CbWXQIn0/FtDC+SabDcuAcE4qFBYP7xxl/E/TzogvYlJu8zfLpSEQuUhyjVCm0hCU/oxFjXZQxoP
/6oHkwe9D+sPVaTWDe3UEOeWG2h/e2A3HrC9XtOfZgziwtWtqV/JzAIIwVnz4HW1wMz0r14CqLwb
G7vl+VAdp4z3nnxWwiQQshQzbSMHsB4/qTlEuq3rdpJ2LmTK8eUkyK+YmGwgTx1sV8MaTLtYGqzO
ZE/fiCI9UaVeFerOIlcna/sL96OlOimy4mJyjikg0ltAxCH1+7VsWooTUYeKmJi9xNwTSjKy3oXv
+YJOT2DvTZTGeFg8zIi8DnfyEPpfEUjOdARfozOb4FSoOfKh03xGYZjq1WGYxaHtQ7EQ9vhUjRyF
shTUVv8FkiBPFY3KZjzbTbHEZJeJgBaoNuLUV6VpY2BuhIHtP6hwPrn71vwjJLgfiuPJZlfSEOSG
IgxNpoaIUv9d33Ges0ibs92Ss/mhUIp1fJOHS+jixn+64T44t9r710vZXiHeQsXDSmzWCIjWJ3F1
/3cK8I4NaOr0Dq/QgRCUERe4ggCTQGACtpoieFRBNxQb/BbvWH4yT61hP/21vJSja+7Dyf/VDe7t
kV+fyUmBNM6/GLI02trpJos0ebJG3lDe3bEyhPgaSQz7VbjEY6ebMSglAty2Y+2R7Hsc7a5+zbh6
s83QE+R1UNfWfsHTkagLrQ/5GfoLB3Typ5PCcIO0R6BEcGrG+jVWdmcgyxHGpPTA5Yb232mwDLH4
N+4sjOYAm2+FDFldBRHHfdLUJ42L8iBCBte+GE3lD//h63bEU/tBiYhmZhB7uz81dFgiiHMrwp8M
S8hBec7d+qVyiMKvM0NYpETb6RfxIVmjYrCVFdKM+gRD0rbJwaQ54o8/g4hAH4x5SYoworGtbgGu
8kMy7SjNVzQLTjzSNkFYp5Rxzt5R+URwIkswMiOX7elzUkxYH0Dny0tHYn0BmEvFSuU9k/zEHhJN
qXMzR0i73mW3ufQKdcBnpuqwsyPXbXT5IQBJJ8Q3F+OluCJPwKRcpZpohTNcr7y3KfjerZwZheZw
dZA/GYEqcmt4sc1zdZCg5N1IXPmpLD64vdYMwYad7FMyTApHx7cNl33ekHAnVb4tWN+nSyhA1B+C
LPVqEpirGn+itae97iAdvO/Uv/JhKb09iu6Jeh72FfSlA7rDE66TwZNubFquFfX0GSzO8frV9FTF
ENid4D5ABNtB20LsN0uvtwnThKAQDMuLfsGvf65MSa2RivIlJh4u7ckmNAQStbDtawBxYMGjwAjg
dXy/q63mKYWWBggohWPXqn9uEHeg+4J5NITL4xX+FxAD+nM580XbiJCnT9abSUpiTqfmgZ1sMBbn
L6RRBL5Wg2vDJRJvAOMQTL4Es0kKFP2uBn+qUQm70cy69PwzKtDxMyt2g7NJnFWZCfmyeT00bIli
w/VKMAtVtBQX2PMPwCDOBi+nK8xLxqECmI/n2a2GjMaPGIsCJVDklXbh3GQodA0gRX7tPrBLeVaZ
f3Z+Z9S9vHNORM8k3DU7p18/Efek4jQP2oBq7Y6LH5b6EHWO2U5LCMF3zmMaM7dtw4opZLHZzDi9
orQqEcDliJcBwVpcvGn+154qBo4s4UH6QYgmzC5OO6eJdk22s0rccp6+evrFMnBQvxc/2h2lMj9I
ExC+ZJ9gHrZGfpaFfgW+LUo0VX2oSpgKdVu1HbdZR0qq3WuzGwt/VZFd7BVH9xsKZEdmnOZejvV9
k0oF/dRgUVBlK9S8d9gd3uh6a0TnCadVcVbEqQTS/NSWPzeM8TdtW0XrWW6dybtktpHWZ1X2FT3l
GL360a2AU5peCa+MmPkBsdC45dvdd2RFzvSb8NJ5cOd9Q5vWP7hWePctMwqyhGRrYXsYtBuE4Z9Z
g3y8/7GmfBcNmxZ114e5suAIDJRqQABT/CfJXX7okIZqro3ZkBCDbjvB+2Zj3OEEo6MSBMWuaFcD
WxrxPaqFmxwUlBmApjy4R6b2453WQ+AFSSo6vCyzWOIMStZ+3fjbKC/C+Xcze806PihQ6yxxwplE
ikLKw6gdVir0VtVqTcuw9gJiGRZvKlrHyXtKyLSYROxI4JfvDZMUnDVcH1+FJfN08+eXmMuS3rS7
YbYeLbJXZN+I2AgupB3E55TcKnrL26oqbPbDGjZg6t/XkjRFpEZh20S1qcCGM+b/M6S6oXq2Tfmj
99n1AVMuyyn3YmHL/iqkdw5lpxVtHuom/QFObU2ORx3MYFv4+wyY15qW4qCD61FUjmUfN7wnjSEX
T/VOqHZIsT9EPgrxNc9koDDbS4DbFCcApVEaSHzaQ9lZDSMhLIcwoGSfnp60xalG9p8cMzk/6o80
XoiO61wFbwGdQ8e5TmvrRnalUDUUav1hNj023eKPgfdfrasPbIEcujSYMWu3vOokkjDSCL+Y3FJ1
kugNf6+ZNeCA6yDlRrog8tbSlOQ7Fy2xkXt18UsGsNIoglttlnjcUCukG0pZ6Kv8BTspRfHxsYCS
W35xiCoL8lpp1vtVND3upQCTxEpum0pfSuE114SFvpFl/SX0RGLO/1HnxoNY/pU2po+Smz8qthh6
nNlNSHgKtRXewSaNbeSCkyBgpZU918BTgMDBjzai0xXhVTGT8V9zS4LUrLM+fCyAJAv1iV5SOfQr
IHKC7zgj52ikPKoTk1vhgoHVuhiSxWgU0BrYNQXGlFB0cLn1N0HfQ58yJD3aEejbna0KXXWJL1AU
SjDgtFGek5BOVSw2qfl5l5aWTiZERdcvV+uSy2eGNA0TIQzqkRkjfWHZz1pOUCZFk5c+bk9UAQkZ
FrjAi1FMwxvWnKS841wa0xr1suxSAWUqSXy9A/j8DX6vRRln4l3ao1LQgFtvBluwXcn8AbCsmkYI
b9WMBUinEeDIUOlRv4JKiTu6SKJtiEPt2oRI0NIjxTpY0xVKy506WnBhNWRLHi+pOb/ETs6jdMJ3
0grzuZD5uWzbCfOYx4A/VawdYwFGcSqD+xVh7bN9ml2hCIWUtwSLitbhEyz81hl0hKdniSfNcTLf
AfEwgH5FjKb3azjBnXJkblkSsdeKlR9HlH5vgHNT11oSlqaGnHmC8UgKrm38+HC7+K1qASYXEalB
/KnSR7ug8J+9kda5w00wnsZXtCpJfgWMUerOGryl41UB5VrOxaHwTJ7arye81xfMSAZ3yn4ljjcd
L9E9t3UYI+kcXUIhJc/OUVJ8O5nHbXlUVGPD50dc1iSBmBlMnudO/MBFOM0hJPy3UIPC6eKvxOcI
MFe5/CzjX/q0qwTmOrSGkMBKHuUipNbT1JEimcefxtcF5ud/85zb8CHm6xP7w+5BGDkuy/tnUwvE
Q5l8hDluHzv1OfqxMyI4epWRHTTbWoWLtqmdrtWI10xMNANQ0GO9jE3dINWHDInbR70AeQzUBQ+6
3jp0Ikk2VtharKTzUNuBAa6fYmc8RmT/HHHMlgT0cq7ZYy2L4ytGK+xJDQZ9LNo9KBrXHugQ6liq
HvOcKK2ofLX+2yhQj4wC2WikxnDpPeIsNIUFxQwTNsuOzI2CmTKVMJ7Zqw3UuGKtLd0UPkvRWUOz
R1W/aPW8X2aZ8QID9GH0soBOcV2+dGLM/P/dmkXWgUZ8mMbDCL0kCSA5NyCZFTvsEbtxhHGp09a2
gYESp7/Iie0EI2UFMcgDi+8JBmwWbqHUYoggrgz0s9vm33gxQu6N2+N0cCy9tPkglSvpzk/ABTdn
+rhbPJAoUCd0tZ0rDx92wDw2r9soqi62RpGqiNoZ5TitiMEAl93h3S2JmMeiYyLzkqsOsHV0ILH5
ORYPlrCbV8KGhzawqM/zswuuJzt+OqoQrjg/BJhZPRcoanpltH79UUVuIWuWBqqDscHgtRxQAFiO
nGZtilJakfkwyE/Yuc4oNwpaf3fF47qgkqA7iBq84JKH/owYx11y9PNKHSP83i+3edl9/9nRAnIf
pPjXLHA6TdqgHlp6rrfjBwkR9O4ta/bpDyk73YYfgYzIaEdaiStKd6oIcXjcOnHkxas9GSgEUW8v
8x/dnKPDUYXqiUOhNw06ZZ6IeiCtodek4+dPvnYT3yo+N2PcZh6aK5p38riHCtfp13me9hzCrq5D
0ON65h5cmkkpq1tyBaTy5mdipOzPAFL2tBazKrmfNp4hAfmVlk0JA1LlgU4+/i0xE2eH/+s+YV20
aLigmnOydNpYjjggnnx39/clj+yXx7KEAJu3HrN7c+H+p2RPM2nc5b+dZtE42x1Kan65GFcXh6Yd
AGvtdMa8edYElXPDshg+7D1yQt67zaqTdfhzDd/T2JLlcexm7sRsmoaUB8vXLmqZoOLLzUlTbr5u
JCU5aFyeOQUSoMEqtQSzyj45EOEQ+anPWPNqTx7AlodPR/sZbxdeuyrQc+OGk1xalBin2Z6TpHzM
GZlZzyefQ0/qSvasfmM7ecaOC20+5PQae6GcFTmLZ0zUM03cQ0QSx32s0VKbpO8JIL6KWteNBA/7
R9HW1FgDQXQKBJ+o4EJdttwhXQ1C0aPeR9BxKrqNlXuLM2Qmq7AKWnLPOULUoCX5JNLJW95GuEm3
sHwUjab7PtU8ilvJVffbz3Homl/YUG7Hrr3evbnwkslaVY1sf/U/iC7+Qd7ZeIs+9rXMsjugEVVF
qgeyRj5+wK64xesDH6b2VghRD+wu4NSLqwL5Xln8aMpDDkkEvdZxCWkCPIW4hzyuzi05T97oMrH4
wCWAt0f09EhtWH3d+EsBQoLYm4ib/WhOzMaRC3gV1lBN0X1Q12/FjrxcfwfpYRXTn5u4DSuz3gOB
AyNRzp8fWKrvdFslq2odQxZqbOmiqE9+ax3ARAC90nZ671akYF6qfeFuKv/swsdrcO2t6VXSLEpJ
SZQb4ATZbsQ2XaP0IyWCjF2d2JymAipUksuGGrYkDgflbuINv1agontKAgq+bTMsovhQzAAkBBh6
ciAI6ULT923Z1vaGI5whJlFON4IOg9aJjaS3Mw9vkkMsAlrrZMa6iu6IKj0X9jIl1aEO9/bN32Lm
6UzJ/PiiNUSp40mU26iFSI5SIBPD4U2vxiKU/tVPJyQigSAKqnNi1DDZABSw10Jnc2DooL9/RtMk
7cXNk1bzenhb5IKZnw7hXhrpDXIHv0LvS1gfDPqQ92Cs+9zW0iRFKkuvf2VCfmNVFP/Ud0z029hb
PJMGraWyLuoqt5MiAg89n3ne9LYAP93tnSHdzwimlv8ML6xpYgnGW0vXD8pKu0bGhU5pI4XbRx4w
P/b7W2sS8PHdUiN0szmIg1ANHzYClGMeklUq0iAq4NODUpoQUMa3TiYCH83kJcgkx2MomVUJCRKp
MoJeyip8F18tEfWVZMb7x1D1JDReXgk9Tno8jh9Tq0tX24PK75SO3nK6aBnIXzx94c2GowqmkEN3
9OaYPwE18fkL12CYxhi8oDQl7ARx/Yocro2j2JfjqDowS0+w91h9Ok1a8XfYlZcXmLdesdxWbAYk
m9U4CGrAnhyZ2LWJOlJDXTAJMuWb44xisgr5PX4VKUKea3xZILKIgXVSu8G/AVBEDXpolXICFiIc
LBaZkfkkxpJT87ST72TUtDAEaCuWjJtrRlgr8VR1w2zp20pIWnGvlmC3DH9PYQwfFljoeDIH1WiG
OLFBLOtDIHNsyKvq6srsM5pNyvLYkGTpQUEYJsi7aErXQoyF59IxVqS5/Wy+UfiAhXZfEDOlnRc4
2pmDQk3o00gSjkKi60X2IXuvyjrCG7WaNONtsAqFBQBcaumrshB7ZYkdKWlHapQ2TBVm+cb8NRw0
f30+qgjdCv1QJPWaTrgPoB/6Z57TiyoAHbUhw9M3BSxUnPT/jtv4JPGgvdWmlpjnGYB+DgTdSG8V
yX7IJQpt/s0rghUtGDWHlQ6LN9Ik48T+kNsbmNtlWXL7UL1o1bvM7jP9HjSMnIrcaW3YLI09NXVv
rp7Nzy3dYY/Z5cgAP0yNeafRfHCcQljNKRkd8spRcke/bUORoAvkIBz5Wxmn+YsLEimxtq/komgB
STCMgboCciO1evELCkeD/RlgZny5S8nXVeV+If1KixFlzsPrrR5LvonYwPKsUpFmBkNXlcKKxCm+
ZzSoCWRN/rtQAdVGCAocxXENs06u/rsvaWtX7zy7iXfm/L+KYNB/9C0XNWelmofD4oHORBE6axma
t4X5f5wUBsxxSB9ERe8PHYlwpAo0zWMOwD/BwIOUftiq/et7uP22CrvARKkfeZZpS1gA+dlydsg7
92uPNdrmdJNLFo0plFgA2O2s8dof42whQzN3wjVCmsiN4rI83p3aSeL7ZMy2cFXaWQeTuWLB3Oe8
QK9iZ9OV95u+ihsw6ondsrhjVgJ/GLnRE4+mBVVVkC6VOfkiKJnRovYFp87fM6cTKVhC6DFdYM1Q
Rmb1Ty9IinJxJtZ565SMrVFuRdq7S6ageLdOIV1XLzX2YNxj1a12NKNvNjXkR/6FxfYQ63qqOFjn
aHMVom53LNmOAtp6xTKElfXt+kBBV8sevDvt2Mfv8488NHyvkOOr1+EHbd8BPc9voNjzRgB6tqnS
XQ+tqPKPI3m0EB/YYnNU+vrChOunm43Z29qMxyftgl8rC1qpd5Xp52XjM4RiCnzjR9aTcLRcyulR
qWAkcURXO4ID/zzmVI62Kz+OGDMBcuDIVi0v1GKKlStBwiG5rUfFo51xeEBrnCsZTF3JHcTZNcoR
zZlHBKdhyk7r1i2/Rlj+62tjLVD4HUNwuHSKsdBiZf31UsZ88dE5XF+kLd8UOqXikvNIpIR5g3I2
k2l2SMyMF7bBLGhQoFS6pDLLlNWR/OiYhCMIznV3xDP6JeXN0tvHpqdxhC5rqS3lllrwipOXWJgn
7xmNf5ydTvblIO4D2eE64Jtb8pXa/Q7pAlr0+sBmY/p2hifuIcQvuDoavxkxh2V1C53hYEuFCEfZ
f97LG0ICJUMxSdWptc9/6xSDllY3ogp6GUWSkiL2rASYGpgRoL4+6RSIke9aNf3kYcO1vTjfX6m8
e1YB+Pk/loQAM4PI3hU/CWxiV9cWHmREtibAWMNyUJrXR70/AmIbaFWlswBZzmrr/4eQp0F6vf5X
T0bFu97K3nqCt4Lkt7p2udk5OxgVoFsgPe9TOz1CNKAebhSnqTjvA5b+q8ZHWC+PT0uHOdut3BsY
bWgxT1gSQV7f+4TNeARkpxKAUwwMtOdwunQEH386WWIg0V/WHzU4IkHv8pSiRsnCGU07RvHDSETi
cRf2cuIFDWC1ukLHK9pjfr4uahPV/40UKhm6tgpcRVOXILJxFzb3c/WAWS3pKu7C8XqwVfTjR5Dn
JjPjJZnpxZnCAF6sY7j+cx9qSQ43pu1fmyFczgewgpIaqBWI9eWM/lWxKL4LAmlF8d1jpzv98s9k
QQnBOa24XEYm0tl4a4nqM+D5vtG8MW0mnlyjdboSQ4Fzi/qOZ4/VsiNaClgrijkXmDWiGQwsyA+u
CjZZOJKnMKBZlzIi/sOy+KxzLCe1HzKRm7nt/hPkkbqp3NyyFs7vEZdNqBpiLxwHJoHlSZ3ljtLM
DuRxjNSDq2JgWaZR4Bfd0JLy2vDsEES5UxLekL0e2Z1od0EDJEIRc0fPICKA3dljNtXJwI1nkp8J
rkyUnNQtg9MKVHnzC3xQZsaNnMljMJrWYaQRBibB7wbi8xg3t8FEob4fQcxd7l+vy4WURh1gHTL7
KTUS/nI9t3Ul/N6guX9E6rY97ou0Mz0UsliyuAUzfLsp/Ujyu59ni0rc3WmruIZpvx2nNfcEqbIr
qK7iMMQelUd5I3qwGk/w2O3bFnk60zMGpjDL2EoFS4cReBKanElwNDO3tXxnt3b5Dh5AKWod4/Rt
yqHrjcQjLByhq9igoDoPonk46/JXcPayQG7EsHHwMqpMruyZqJxyHH2oK0ZT+kJGaPJUHbPt0/1q
zTSI5E5dqIGw0ZELM+AwgguZMdCR8KfTx1euonv9lrQbhqK5ki0X7w4IkJ2PCMZHqI7CbPty7+Jz
vDifiBie2XPDOwNJfkyBr24Ti/VIkXwzHUhIO0DVEIPomRiEUpo4PUK50K78M8PP6sxTDU/tV/XA
QiU84gpGNhUZPezrShYYkmVCDq6BYCb4FYPs991WhAPeZ6+i27tg02hLLGBsQ86AFsBRAXvk5JIJ
v5er5eShgMQTbwwTpq5Y1nxMaVXpPVnd/aIkWHuZYKwz/0AgdOWgbROy8tcmcLAQFf6QQigxZp0h
1TqIl6C/iwkh5kT/spJmuK/z40u+1bDOXvN/OSlmCpAGKameCwhC8323VY7Vb0TWv68XZcLzaZXJ
Z1Kcg/jQQuIkWqhHsnpR+mt/SzOv+Nk1M/00Ls1slTgL37kA/qvTc7umqC1x15eGdRGhMsrmRdcj
YsVgA/J2nemp7Emkpqj0Vp+TGK8yivPvW3gZHzIp79SgUg1TsqyAodz6TpuFPziPfLKi0RK8klv3
oNiPpsVVzylbiK78zgUSCzZPKTXf+nOYd29bDHbzbi8C0zg1BTQRRBFM+n3a07BMHNn+fV0RlqWS
vTVDqHbV5Gn1FuVPVHp3UZHXB0UhJUvtB131EOJlrXXNsygwYgoqa2zX2kuvw52tko8o2Yv1tQB8
XYpkn1/tFK6twDYpTVPoO2OWLzSXhb+f3cMHWntdQsm2ieTXjJaIHtNZC9qR82N0v3+KNMhm9u4w
MfTGCpECi8H8odV4AQ+Yb3jzpFHkdMlivw9NUT3rd7E3KaAgaWcsj+vfrcULzDtDDUw/0NYQE6xd
wyFRUPdnFDPH2QKew3CRJcTK/GThtf79ArMLfolBDv7ENorHLB57XRnI/+PualkXQ7xk08VW1cr8
x0gZScCtWTG7RfOR679ElmfwLT7XmJ6LQ6dOKs9LiQjlDe32CaPpM5l8kqQGYm5PbA7bxatbkSxF
DBTs02owfHJVhPGR+47ExI49jeqCvUli066Sd6O4MLG1AEyLHMzQLkzhxuvNSBhLMlv2uwpyecHH
SkpYFG7V5641YVJRJsrg7bi83LljEkPsKl1TGJtnZH4+6Qy4CasfVCtiKshu3FV6VPZuMXfK1QMv
zMSqEsaQgCRVGKC77pdvtcyQ89fEXkrnGPKJ3mkbM8uWg6oMywBoW8yHAfyZzTiJS/BYPOJnjReR
LyRNTdpkD8SkHL6AYGDWurS0JPhD5ftqhJu2m6x7q++YOOJkaWPxbnNg7fnC313uDghh+MTcaX7t
eqggLQr2+mExqnJEr2YlEtzI4srp+xd5VnEw956Y/EuQSZaKF4SbhlLxMs5EC0+p96a3hNPGqnVJ
t3V85ncMDshuxF2ud8ajPg315s/7eAippCvaAPeyw9yOo7sGZC64JAFjf1dJl1tHRSp34EbS9tBa
feTh8iGBeY+aOvq2uuaHPmEyOK2rOg+g04nF5dmambhrVTsZyL9f7mwHzmWW2GsmoUKCg1yAelfw
ZKyycewRffvL8GPJ4iTJbohRM5Lw47WIOFBlyacM+yC7ppMTvMrr/4/aiyak0DQVEj9e2i9oaP48
12tPc3LBQzfuBgWQLtPR6aC/x7R6iaSzm2gSop/sqeAzTEZuqkLfCE+OXiftjMeYe0bQ4qC2bAMB
cF/Q49D2Lp86aTF+6AY226s1yA+5gPagqGsZDUp0Gq9Qgt4A8w95WcGYA5GJUs4adW2s956Lp89P
SXs1knMgutXN1+nM7zq+SZ4E6MdsMQGBk47715N9o+XXFWvFGWMY2UlXcRtDO7IL00Xyvi2VxiOz
GwXrMFIDk0WnkwBuIq1hYzLwRqNgBXB+x/1q+Z4eHl/MfP25JiXWHiyzFI1Jtz5njvk8rcYuryr9
SP7qsnr18+Da54gMPepnhtx+kq68sOJ5lJi0JZLQfx0fyWY58R+yLLAp6ksknTykiFoiMrSz2SiE
HCjZk0tSemVd9j4kold4dHo30x8r0KFwpjHDaAUQ4W/YOCbeegaGYDCsXsWyXgVAoQ6fD76Jh5jY
6fD3ri/6B0EwVUW3I7WE6ckK6GjnuiUkyR+8Jt0BQURKYWKvRFgjYwHhB8HwKhndcgxqeJQJIrul
fjzZfcxLagMwOv5WzuA5DAJW85m2OJW1+cF4WIL9EfzuxtXFTf1YqUwSimPYKR0vj+xLUbBv6/UH
iOYRTReZFM8ccLJJ4CCbKt9NafX1/irBl0tQB3kILOx0ukXU3cbV7Ru0cB0g8yeOOa3Ub0UKnFX6
qp5BoCAcb4sXQPuCMqMI+W21ZwMIWjeQssfVoxIL6ktFkDqGeOewEjJoJGqREqh8mJ4WaC8p/zOn
q1NjZIQQYkIE6g54zHhTVep4ppLJGWEDG+zd48aZU9+L+sjTx7q9rr4DKL6RYFGX4SUnaUm2iRZh
Y0p4m8teU4cswobYJxdBysrA+IoMYvhCtkJTDOuGqSnvLa5Xv498b8spd2dMpp7qy9TSHsPzlp3g
Eh90bEqz+7+6Vq0cczBAVGbSE7b5EvXmhWLKnR4E2Av7sv10xHPONp250YnseSb2swAheToxbSM7
JGFRysNHrAN5BvyeW+zruP0GZYq6NCwK6MB9lCgQime6dYmh2JuezbmcFtz7az1JvOQM+M36Gc20
olAi2ZZCcTzTMZqRdkOTkDA0jG9ME+3gRBQBNTQ8Tqc7ewqcMemp9eJGNfrsNcMbWetY5+oHj4FC
3vzR2Uqj/B0XdDj2w32dzZkzIzjld68zUfL+jBes7y9qy1TTSkKlNHDQ47d3UKxul1iRr82QNS8v
296okklsOl6bgENnmKJ/X3/u0Ji5MWntMvnzJeB+wk1+mko6+AJHNLAZdR01HOPZ2LUqeuc1kV6J
cuz0hpXPjuGKn/13OVIBXgerJn2Xa2yiLDbK5wIqXx4vKHjpK0HElStNQzyLNIhD1HQHD8BbJlZI
MW8D76o+UJ+qCNzZ+tXptsEUzLBEV/oUlqacCErFQU9jSdjWe6MUv4EMgc8DdAYyJMqZCAclPrQL
Jilo839pzxMAPjkSNQ4Ybwg6pfXRygIjO9CWIvc1McE+k6tZb6wZ730r15w0lvywueC4qx2CY0VR
NKye7UW/SwDKUfOJY1qJXTkD9H26vcirpezy2w0Em8G4xKm6n+mO+S/8xKnYwToFESSO8arP62Re
CT8F01iOC0M+78TxfzHS/MCYGmpeIh/FLv5Ak36dD6GGwf7459bqTHG48nasSimCb6QBgTrI9P+n
qyidv6p7F1cbtVg6tFDU0oM43+VG516EQpNEHtfF7adLbNlRLcBylkChLH0DIRvrD4/Ll2BnEalt
JM3/HMW4/ywbBFaZNfpihjAVBb0bsg/T82Q0RWdwlfaVaYuTKyrizI0J3ENTI3ClWruoyEGuSA4h
cehPQ3ilbqtuo6QJ9xEci9O69kRqLqRAcQ8wV45NEXU+KHtLXP9n61qZN0oU1GZV8Ddn1r9MnFeT
Dg2sR/Zxc5NOuNnUowB6ZbeAFy2TLruI91DyNktmY2LJcXNQZ2YkStXgYdriMAfmgBxtDocl0b2u
r2h064TanPQ8NaHP5AyHe+pcx2GeHhnob8ikH4dL/f/vZs3DaKZB6Q2j1W6Q01773aKpj9qttb+6
V2c7vHsW98LtnTpq2b42WEodlCn5VKK97mYy1OWk3o7JLBjBendjjER3Cr+1HKs8FbV1JvGaaC3g
4EW7X5txQxntBGiEoeVKFIR1qH3uwupKbjsnc/CE+ViOsYS/EoRY18HTtdEwO2EfFCjnFjlp6n0d
Q0EcWWoUunj9Z7Zil7Zwhuca+yqyxCn8Oz/U+yLsXdGrP7iFdNWiOO676//guoN/NlyWglawzAWT
FFD6agMmZu0wDJxG/HdMeAVutsVR50UOQ+r0zNcFmN/17qz5k0mfWpCjrRfoNqjSet6aT29Na1bB
1/Qvkg7G9k0+iD/K4RNe1qMr9LiACWzK4zkzFPvj6jF8M4iKx8MrAO4tWNby9lvVKSX01C/wX1/Q
j+1N20y5bb81S3UhNGErxxh879E9qdTomde5D4HcpJl1nwjLKBPbSiCmU5d5/7GgTQk9N8ZUvX++
h7z+iWWbwVRPGeEGlfGOckOfeoK2deOK+gDqD7qs+MrsWyuESyhBNPP0NKEkRC+/4ZiQrCM44qPh
v2lzuQohojVtpyyvwTe0N6i8jel37p9qoYs9RIR8SUGxF47qvsb9Tv/nh252uDIBDABNhUdOmrfM
/eWCmU8mMq3jTK9aahENaHAw7ixrV12xf4EDKWmfNfN9MakIWTssfZXk+qioKA47AjAI9hWCvYLS
xW1FXB6rzz3ZtQi1rL9QC6KIOpmQblgAL5zoESlNPNlAcRdh0QXOKPdhxr7u/1nPLYlO/Ss1E8m+
6qxWIDEmPH2WbznaZo2oAXHgTNIuckBuDcJI+dZNL7OVRh0UXVn75dDOUtXNVs5ON9TbpB/9g/Js
YgVufzaDsEhqjVATqHlxHDatT/guAmtWHCaHwIQbgE9LDZJgv0uJcj9fn4VsE564ZSy2V0eprtZG
mQ7rca/xxi5x9deHkcRdY13TFFyckyZyW3sbeL1tnrD0JCFXP5OlTxjrzjld0OeotrKOWy1Q4xr4
EYShRDoFv8Pn9EwQTkz4GF7WMjCtLhGZSvw98qyuIbvzHxUJkk4Ov/jvoikR1TUaFNNcyNTuu6F/
BbTIK3BZGgyodZ6akp4YjghnVEp/UceqV6A4+o4znHXs0Q9X6TbTWFyH4lgkCZGtT4lbSo/KGpSd
kPDretVD+5oFY4gx5Vc9wLXSekrne+aMaBR78yoeiMcQiFlH0WwNecLFWzj9agapfhlfdxYAMRbN
R5+ZZJPSNIvq406LwvYGNTozzSa/khItHpEyNM17OUvVe5hLygCtWLGc1h8OmY/Lsl8fHhYqUsHU
eOtmaGXGvpzi7+i1XxifhwoUopVgf/LM1/Ive8BtVSKeFyW36HkK+bnaaCO575lDTAq45nHopiMJ
Vn+oZT13M7aioqp6qXy5Sv2yqY5aGAA6qkZOGIkMyAUQrOzDGoUIk1Ih6D4nzJnMBpHhZohvpJc8
pTsF17cXoinvGkxjz3jJtvSQVLvkNrlE/62z/uD0fc41jU0ffFSFO6qL2Brvbfv8Kf2weiifNAFx
nN+nrpr+NNl881+LzWkyxJ1VmOTeh5v/nRg4y+q6W9Z3zpy92Qfe+kHKs8IA9BvrUXpJCRa60wfl
GMpJUygTexCkIfxqScf5lRl/bxHdVmV6k/e9SJB13IVLAvsYRXSktM7WINktsH/lfY0b39fa2vlE
WxsP0OTvdv5ef6des6+qz8KTlCCdVS4DF821i2rVsdaqGgQLRK2F9oXlScYzTrodz1weEoipnUYq
dVHs1NgkqaDMrgsko0c7u0j4vrLJF410wX8PcvltS7Ap5ElpZCncLU7wlnSxvaoqT668KYpz8n8y
tLKuM+XKVct8Ch9wkqqmHHrQaDgfRXGwT7fH8d1BsJ9XyVUE7//DFtnfN9ZDvtr5qOEmrS2+gt9e
7KMxTg96DaKdmnikb5hanM4QxCdh8ov/xAvotKPd2IzejuKxz92Hf9Dl/Ln2pP8zus8WSRFJ0fzc
ovmV4lJXNjSYyM9/D+i3LgjZTKA8S3gLR+K7Norz3UDlh7rdzTq89M5Kh7j8f4gRKCfNXCxj36+v
G6CZWD+VC+UOFXJc/WM/YB1R8JOtiY2kbdHH/K5SnebSVnAF58/kc3RcGgAQIchdqjDiKFjdH2mm
dIJccse6Q7zziT/tLjiORJe3q+8wjG37JvHpurJtWycKsZtIaJs8/IdxZmZZQKkaaVTY/FzqMYoZ
aFUTD8bY21NZn/GuWveuhL6S4k8VvsWpXLJeGNsIq/hZnF44qzRmAAM6iP35A61Zme4jBOODLUP1
WKW01VNfK9s7ua4fJ4yDXPovLV+nz3OJbr+FP8TKz6OXIQDYMRBe/Xz3KmLt0ErK0DuMKLH4Z7rm
OvI+IYXIka105QES7iYndJg4GIESy1oDYDe/wRvI8lEBgin7prAKHlDgNqO8v8DkczTksn/P8EZ/
/H/FlMUO0Qtxx0ieo5sxOQ5NiEt4xJrNPJmImaRUF7yhJcCKyWHHtpqXy+3RyWD3lUnoyVJw7Ffv
0mpOhh4aLluJfe0NwMqQ1N9W4GdoYdf4NavAISl0Xz7eSehVtS37i3TAnReidAXsqj4aYYDrADV7
nGIaqgQQv3e6ceaxugM3uTy9qFCTRBc8WC2lvF9tsDwF3qOy2VKZ8/QWG/47aBF0Ua1xnuHsFYfT
4Tn4ovd7Hgk/Z3bUjxdMyPvH1rxe4pSGFhdHQ6q/jd29iyDF+wnOOLp5obVIscsPtjzCdTxbviP1
BDBSAmN4+lL3SCwa8Q1KnP49i9V6ZbsciTrhr9Q4jPnbEV9IpQmBwzcJ/pdZNhrunTGj8meAneIU
dQ0WSg0D7QIb+H6vbyXoXnAgGsI0c2xn3ns5KzvrPZUDm0KkFgOpmQNfb9+SLxXBJVkCIsNm14q3
KMpKSW0YkwiG1X6wVLkanC4RP3empJND+a4ET0zzN3nDt4XFpSsHeLq7xPTeV7k+cg7JqijsS1G8
yTudaJan5Q0mTDzfCxhSGNjuucPLzSJGJr1c9DQUFnhrutMbec+ADgU4do3Bwdt5ZkBe0pf2Puo0
7YBhdHhu/iqraiZmje/4VMIsJqZybknWh38ltFdJoQbSwWZJczuFXZNKyyiCIdPDmKJrVWlwSrhW
WItIMuuahhKB8qqJYs2+EOF56ldd1lsspqM5FabbBh7kZi1fg9Uczjyf/sKQqxxmtLVL1Qyp6CNQ
DMQPEPBSbwSmX1gM9wFuRng7kfY9Q3PaU5d5k1W46+0kYYwY3N6tiN3LOrhExmVF6p90f/n0PQIo
Nu+Rrobg3LWau646SrxDmR3F9pXX7o1OF2w77JB34KhUMVLanGzboDvfOaGwg9hXQ4/pBgD32w4i
x+qlFEE9Rtrgan/OCQG0hHlNC4eu+kEZDW/EGCUZOWjxyATI0d5tIPpYuy3m2eYqLczYtGSz0y5S
TTLKfUt7nhaBH3eZr/XirnK5f072Nvi2E0dkCHH0XpWiLmy91QdrenHWpMfzLxfyfPaHqkTRrx0A
mZ7l3Fo9m/egwue/mfDynVTKNCFKwXTjhatqbqe3XveezPKxWNtiPpPjJrxnpnP7+7MI5Wm+Ymcl
nPoY9QB2RWFUVO0G9ZSQySSvHga/0ATKQ9X5b+ukyg46jh9XxE2gFVahc23Lx2thqwULnWdMcSDl
fmLmCdR5x/KHleP7KL7Rou+m1FMaM1l/Rp/uNs3+T4ezHwGyLppa9RhhKWopY+ZL8PEZklDeyq5L
pGpB5AYzZvUNhpsOpfwJsZ2o+26mn9f4cjlCBF32BHwKKrVf9ap5TnqyEX4K3wVI37gSYPyKfsa3
Wxp772HUKqH6FeyA+qqBL0rPTZc3pCx38bwdSo17i2I0JddN92Dz7YtR7PtArcSg0Z5TTk3zAGls
7CFCH3gsvDnfjN9xyIBSmi3ZHMfiO1qyP2s24Bddb1FfSk5LUDcE6in/KQahuMmJrTGZRnBba6th
iTdiEiHjqHUjcUH6W/8H+tk+kJqlD2L4FxUhl/+cJQFz2U1ZNG1GyrmM1/ODQfhuKoAPxuFHT2tn
mFnuNMAVDsVsXeqOUif0C8JLNPiwIIboXE/IaS5XhTHHHzajx4OUzfs7l83QowHFSLqftLam3mbq
25ErAw65x4fA+Zio7qd0lvwxoU8qv0Qjt96r65ohkJVlKf2x0KC9d1qt+D1tWgx8ttuDFwr9+dC8
i5p2nruag1xaLT6OjFI+R/8HNExROFELDc58MiKjvvJ7QcoIdCaUBdg8MY00CghnLRMDMgfeLAXu
uZSnlDAjm5hLFMdvQ1OfbcCiaamPoq0Dmcug1f6cfw8bvKi+ltHIm/Rfcq8gNmhwRQziL+2lSrjZ
52IC2nBW4DFfjnwcLLMC2M9RE3hT4B9C/55TvH031u45vozq1GjUc+l/Uw5pldHQlfO8SyWj7qN/
zAtF8N78BD6qiVAr2Va4YgYe2DhmI04TWb8NQeLfxzHCzEUKkh9YaNxhuVccbHnV0+/UdJVm6q9T
ktvcli8bza2hKKXnewVCWu6oS7uM40srt17NQ/Rh8D4X90EXkPNMJmuzZuResolKlWRc8tW6+/S9
c6vgpnkt90R6tD37TUbhj6E3MK0aoMPFs4ZycUWNCcxpCBxb6zpEDmLpd0QQ9c8N7Y0lEm/ZoAut
Ub//TYdyfF3TH9x5Cgj1BvN11SyD9ZgbhnJ+pESunSRDX7kBDDza6+VXRDNEhCgZFUVfxUuk54wr
KjUFThAyhEcnqIT1kLpj2C8oM/e2B4iuKqJUKXOL7LciDPyq+g/D7vOeIZZxSV1/V6NkwLJOQceM
wFkCh3r5PWZ6YlpeFNa2UmaeEgAI51CQs0ii2auQK57EJqb8DfTkzdrBjLRGmG/hKhNYi6Lc0Btl
JV9WBFU0qpjAJZ51A950SMqIkgdJhj/eczMZL0xv7G/qhcaPaGF1UbdvtkgwrgjmIIDKF+Pi9OqK
D02sFXdeUJneczucKIejjtgA2p7l21v02H4s+NfqxiDw4z3QhTlKiNpv7i8lfIlL02JLf+SxK8ib
B+F/994g3K4ee9vG3YuWdNztdPBeWfmVu2We6Gs3GlsLhkPi5T7J1U03jmiTFYyQka7npRKi1PwF
3oHM4UQ+zeBJFV3rWzW/5ivaQeL4mALSuyFVq6qzrCPzMNNRHX6Cd2XN1J7AxusPIAJcfT971hmV
7u7f0p9nBBE8xD/Ntxt09sYgn4WZRqtCHpnI2DKpFcQMTyUKAigrIWsqzkBQC1vYbkk2EoO8SDiS
v4tAo924bqvmbXLngBwc0phieXz4FoPIzDCaMAeLSNYWxrf3jOXbamamJPEq6ToGap2/G6wBIFAt
IcudDddAzTZkroKCmpxDOU8tTKe3XZWkF5OFqwtzsFzCGhdcUnd+QBJh5AIxCrJFDaAPjtOtKd3P
zbtHce/BXACPhA1GcQlAj6EAeHDGRkRWT+7AVERo5wiuPb7nH2YnvOCwZwz+HM3U07GjUr87WY7i
GWMYojXyDXwM3VUUOwPjupTT51O8rKx8+k2W71WslM3Htv+ZtYwnfGL++f6088OKDCzRYevXwSOb
mgmdt7pX+cYvDhhryWkHhaPtV8Tj5ebnw0Isc5hQCs25gckfSbsP/tQy501oKmv2GQyJSj/u1OqJ
LDN164symVgD15gdFY7SvoL7Gw/xsAxQC/1ib4tG0W1LoSRShPhN6y5GRZH8W5a6Z9VhKcOi4s7z
XJjDfeu+5sSYH5cKaSvftIT9m3m6It5HTZXhmiYeetYtIxbsMZnO3HTry0tTOq8gmTqsZpnYk91V
J67XBRe5yhHbga6xShXKI2jDoDePfeY6nYq9pf8pX3KAGEApMUqa09oPz8MtOHSgtnVhirAuv5Br
lpOG737iBrfB2mijhE9+/zLFzUBAKXYcSaNuZm0EqNCFhwjbTBDZXF4CF7+CoE+OhLDtGW/iNxp8
7lmIRqUx8Nh5w14H6EhDXmSuTQJS1xnx3hKGm9ddP4Fbtt/5/NvBkOJmlVxCG+Ul/Rtg+Ae0qMNd
yKOBR12su+oq5vcwaeHgn5389goIXtX9XB51acrzFMutbtSRfzyY+x8gKcFEJkZNLAo4j3zkKsNG
/2lhZWqiNTdYehcp6sVnvcp4KQqALEUMlvf4cqXObTob8xZQUp2PGIsJtiC2eCbGYJKKYBZwaybj
NYkZvH8qiVxQJST/6YoZQTAmg4LOS3qp3jcAB4wXcEeXoTepETXYHBHwWcQAKtEABhyVaWlesuux
yvDRdkHcNVmxqs38AMBDOKAmlAsvi/34xZ8I1Y4iWh1W9wkWaSad3K5ZLiI7gvfpV4BF03daXiEe
20qI5tezYP4wPUV02c7Nku2MEXXxS3XSO+fvsH4J5Y5bZWsgfdxOdfXblTziremi70B8XodQH7bJ
+Yc9vVbR+ziiVSUx70natEIjhsGRvFiF88b4n1HpQGDaBeUPTlXf6Y8mvwB/Wnie7bOtoqOxlLzi
Fj4owjXnD6Ruw4+fY26aMIyfKbohCT+bsMyrOfOJzTrS+YUkddOQH3V0GRdZuxEio8xLZo760gAw
D5ZPYWTF3NaENBQ0p0yfZlP1M8CNEyEe7ac5TS4/lUClse7GmwJXCAYfdHRWkC+IMfLVPWcQA+Dt
dMMRZgh/6PPj8TMqARnOd9II7GnQNoWyqtUWH8/fFpNWrjV6GzZDbVYHlrkCmgN2hpSuDDp1DEJx
xzz3JOyDStLjSdY3ait/OgJ2YYeDoQxtHqUeHKhYHJ/3hVRNo1+javGzpNzyOeTRdcx69spZzvMr
z/Zp5NqWPEMnKLABywnBcrTZTybGBGQiF3AcsQ6vE8Njjv0YIXjAbdxMNTzn2AJmKiowJ1+VBb6z
yt2VWfUMZ/Hlj1lMkJyOAIl2GZJRWFJU/jK7AB6KyXGIiapl2ckWWqg8MQndidHKwkcK1me3+a51
9neqwCzFhEsUyVtk6sX+KFTP7nmZN99Yjc8L1OgflWcYZAa8qaK6kVu8vjeC1EMQag05F/RWMcvs
J/nI8nSzNeSy2QuyQioAFh5oFanlWKnSHZXF7COrUbD3P74P24s/OjGcV8LlCQ8FTd6ANibnKRD6
1MYYM1UtJThUmz7FnuyJcpDXfxyT4mnPZqAs7RUfuR0mQKisNm0DWCjhB8GFkbW9ln0bQeAtJ7+8
legv2UZFHjRs5u7tZWVeUUk7TM0Hs3t+Gg45F1RXSOUTkFV1faWzttQgcmZD2I2p46rEbG9oQIg/
adUU73MqS97qoscOh5j+GJzwB5VSBuLSEAHh7w3rKXHT5tGGEJNFkI6hXIEWTpuaZbyuyODBp0PM
ov9E6lFx8bA5UKvfE8bYhQ6f+s9yR1RAX05BvgMSEygOQhc1wbEptPkXtK1XnGwwwHVQ0EGo1wvB
SsTPSJwcxTouwLrX16OcX/FR9jxOoSHLursIbt0NsV57EHetfKtlJ4PIMAsqKOaAFeSJIHqKT93g
a+pIiC7C4AATUe/zaHFfhav86tYztShuau2KaBxrSDchsltqd20BQ+1j2itW9EvAS3Udf9lYz+CI
T8LTq9cHgm7fjhvDxb1AwIzgto2exMyVwAeQAZEjNXas7r2At4Iayx66DiouYVWMp1Lk3Rj46i7D
DmWOjqhIIQw1dO2xIbrDgLXHvJQM1/QvmUyWGR0z/skFIRa7sQoQJ1ttBOHzA6TXPIDqIJI6ZS6r
EWhC1VsHOmretwZPsdTp0LKodXNG5LC9Vg0oERwbpdCB+2b6VkCeeBV3+Fjo/TMyQhnuIINlidEo
uxKedTYxt+dc9bFHTRn0QXr9jTbOYgtavgxcIX71l8r7q1gLcREU0BwE6uChjTZbdcs6bkQ9Va+Q
IJZ/qn8iy6Upl0qMsu6CMa+S0cAx41TuWhTZE1NAe3nf+0/GHclV7PStJVOKwSsm9umdTMl3GLgk
cg94Q8kXs8J86GbmH+Stzxbvx2lD/b3lMdWpuYXHnyRMWjJEBLL6X49dbpvx3s6Tm0QVmQHu/Dcp
RIOmRhm5FQkdmNzElM+mm4g0vntVBdYv/IeXGGjIEft7cgL6qWRSGGriFnCSTDSgcJSF0BB6D9ib
aCQwS5oswRI8qvXfWbG2ditcY9ga5z48x7cHqDpdYTkuAPezWZ1CoVnTTh2xImgPrMx7FegGtqvu
g6XcSqVq6VzQthcsNucwVPGNVI5uDhbcITj/5Nfr/mDPvVNnU+uV5D7sZYQMEaBWh8fToaMJYJtW
E9tX6czk++zZHERz/1torxh0u6fO9bOds3rjU4wvDa+tcaqicGbRYu+ZwTR49ics9qAYuEkD35XB
AFWjKJzRtORypY22xGA8VrPHQmdw7ITrxppWUCXm/O6KqzW/PDEWWeegePH7fxGGTmD2Yutfwb1z
7tFfsqxIWs0qF2xmlJHSJUUzT9JMedRvp7vf/Yh0Joer7lN8QWv6yvNL/eJ0sVjicEJJazdDkntI
dk4AisCStHQNaFQ89ArhQM2ROXCWo5z4997a2JB9OmI96/768WuZ5gQxLAhhcpRFPrXgOlw0s3Xy
XNu6ss4Kq54FyzKiQv6+HDz1yX1hPqkonbgeaPyT5eM3zJFE04Lh2mP9PAgv0nxEam7d5Jc1RsGN
vqjPIpf1KXPr4DNtduJypCn+Ohzoh0eilfcxXByjzA+6gEtL3UcBU+rWB38JsZO30hMW5c4GaLvO
q3XYMr3ZuCZRDlei5cQPJHNA2h1r4LU6YVPiLI1YZBNyN3QVKc37gZ6NXbJCSlAzfl0elzZbAGoQ
8jGolRaglnKD4L26ytaYHaTTs4laMTbP338nHidJd8Y40g+SJlXPLhH6NhZLzk/jOlWNFMyzQ+NS
QXqUYDjE3WbBhqRLVYl2TzjkXwqNhysR+vZ7dApQeuWuA8rBTKY2YT44+A5l5hiiBfDTGXsBBONu
ep9APJS5oT30wj03cinBQeUVQY9CJnNvbvg46XFjWkVX1YC9tTNPxwPV6YzXIuTZz3hhbIS7MFHV
4NuMnahYqtU5WR7haEvZf0DOEurIVHaMySD5+EJd2ndQ4qPDj6S3p+njdsmoBbrQh/X1HIe65d9T
o3vyAoxpcZJ90F4pg6mOuino80BCLxxBKKDM8aGIgZbiO0pStp9n3HigV+7qx58q57iL3WvJE1Yc
jKWCdWsJCG+qXDy0RgbqFPpjgIBLkv4bETcjGKzeWZW5J8pDeIKJtaoX8o5Rya1rk6mZ/JDF5o8E
BZ9e58mvEvt3FAWU9WLMl0ROOTws5PZku8nfRyQBMXtxPaNSnCw5QtJTBfaXDRfUZBjQsbS963az
6+Mv7tSxc8yTnMFokCFdfAwHk9xpSjHYmUFneG7XzvAY/mDGPOSb4lRRibC0DiQQ9cwFOUMtH0NW
CscuGgn0g3240bPyU1IYK751cWZhRrhTKyKNy8eXzVU6dDTStHL78E3KNpvqgy1/Wfjd+v1/xJkO
MoknK3sCNneP1jMQfe3XHpJKNRZ9Tgp0tVB9fJtd+68mHGV/sIwVX7OZNi/hcGbfOv9tFrFPignh
D7Nd2FEqYfXjxPqVioV+o3+nyM/IPYN+lOZl/skQNaSleRi3ZaVevabZpXI54azHKKFgogJfQYXX
lsQBEAf3snL3wVz6LrOe9v2/a0y5Wmq+u1Qzt9m40qEVwOmd7LqPjJcz7JhehssW+TcNQYkTeBGK
xipMl6sjFjzjsTMfbn3A/l/yG4zaLj+PLxN/P72W7AntJ3siW9hm+w3VQvwvHzSgLrIwlpuAWauo
FOziMmJox7GEYB/S1UdH9zW6LkAmYd/UVZVWLnIAALI38hBiedhrqf5VAcMi7SqMjA3rtXynu6bo
AxUDwhZqfEINLXRuU/SXdeSwVgktdCrd23pmREBx5RRGT1epN+FZ7n5oicjfAkYMd0BU338SXl2E
33HlRnw/z5cCZ4EMwCSQMebr55kSMUkBbtxWPTCW1bxcFblKYQ5I+2zvAQrRSq4curwtpYDIAI1/
5UTfNBS+e2AAjD3HsOKgIGhF8G2Ryhaz2NEamQlRjPcSgfkA2YDzEirkJ9BciBOHUWaXG2fW5MXl
+amfagXQaS7SFBTLyBZdcV7H1Tljoezz8qeJsebIgJ4ZRmv0/ML2iGQ+pSl8VW40T7j5BA3nshMo
8I9GIToQzR0+90xYxaqJulxjv8EtcWE1D/Q55hH1KcVJR1gPP3fwL8UiNNWlaLjS6FFQDeWdskNU
Kv9/D0mtrVgiv5QIA7QmehhYbFo7E9iNjJH6XPjayLaFaNfL/2EJc+fSwEDZ1HwjETi46tRkcoWZ
GbHcR6pGwQ3HSvmUU31HN1lm6WyQZhqNYJUpidosOLL0McB7i6LHBvSOrq7nCNzyTCfcr+XEpXdW
mwi9mbEu60zVuINhYCf7QVcGD9Fja05Bo5ijasxQidwIYjUBbmV6a73NlngbtyWyzQ77UgOgpPwT
IGgBXis6dNs7c4a2pi3f/yKIaFdsbxyd920NEtmQD2GcosAvljg3DUoskhLWaEo0CqY2hYBs6qV7
cWHkz7OXWZEh7eOKFFYAlz0ntSM5kPjPwiPcDvr4+YGwoAPXsKG4PVxGDUzCs4WE3lJ32hk/ukP/
sD93EAboVCBQOG9zjqG37i7WLox5/94VQeCTcfGT+BvgYbTWxWvrbp2Df8r0Ctc5heL9D3JAkrAB
PZFg7HUhicPrCSAllsuX8eEWuB9bPi+//mwk5estSgzoc4xaMRCodMTLiJh/0i1ZSuxeWFl/xeo3
DTMgWc/RVNGEfcpKASZpj17Cig8+2XyRt6+JPC3Dt7dcpyNSfeauS1oW1TcjCl3UiWNM/FCpRfau
PsbQ8SKBTgSCFg1eUXlcdEzsP0bkCmTb52hhQhUWPYGn7MdWoJWgM9+v+4kUYO/dZOz0N+athqRs
S7JewfNNL8OklLOc9+xOi1qW5+w1Cu89o8zTZgKrn5SW/JP6SWANgTVywjlmQiMAP4rk9H2ZlD73
mE8W/Np3K0ahkdCF7Wsu6duST/eRit1axegBX3tTypswzcKIe9l/2r43U3yWJ44+/Oa4FqKS47hE
N+hVukSmzUQxcVzyAN2+GmkqiKxgQW/imARhSG4+l4CmLqy7xnNFpAaN/gcHmqcaVpu0pEuz1dzS
G1vE2wvYU2EpyzmcHKfEytqbgD4ALDEIlCTfivi+qH4Zm020jQ3kO/UcTJ3zlOGrSI3C8AvxLArL
PwcjTR1CrFOPjFdXXNLsmHAYWaf5TKigp/PRI3quqJOfcaxCal5zUySUzWiAA0N6pNX5i92IKSSK
zoktwO8xfdR2UiuqNHQU8fTlNwwBhJcMouL49d2eSueRLIz2EIMEZtO8wwJjhTuQpWbdiu4jF2/Q
WfoO8XSUQePvUTCM7n4dac2huxm5mTiioQdUoKefcFj+6F11RX888KNcGSKs5tgSPuX0cWN5qSjn
q+1QAzAnLO9E5WU9LkjshuIHaujGMHf0bOJ65hCo1LBSXiupBmRHRbr3GPDo5FkB9PEzXK2KOOYv
VDSfCVBDxBcM+XwN+pHk8jjvf4kXPr0fwGsq99MBGc4f9FWiOpJi3xpN9FCPzSPZJ2MKtZpf6v1G
9JsoXTgQaIKhExjZqx4KRgJ8szVFKS5OV/fW6vQzE/uBVvSeCo136Jm8T2o89v2rL6kZm59sStBZ
HNWGY5C6y2zlMVwgh0Vy/NDSo8vwTq/KDXfrnkVY5mzfouJDRtZiRsAdZSn7vXOxGslhU2/dxIPR
8kbqc+zxSFvi2TCIuWEvoEgHtdn0W8hV2K/3+n5SFEvnTfv8lL1dgwwhP/a4xor5KJo7rOffoT24
8ysXTZe8bpzj2TJhvTsfIXnwdgjTgz7Qv3JbICn8wZKHo0FnGlMZrmVvC5O4ch8AW0QkUPAzes2h
DaFdJfGV697v52t25RZ8eOTBngW9F9HzjcJrWgD4FLTcuzlkgqq3k7YzLj6CZ27W0sruiJjtgkTC
m/QR4oMD0UIyCjsduwTBQau0ObPE/fFtYivHsDGR0Uec/Hb5hDMTLgQUpywlUpslQqnob/pAg9bN
4FoIVPVC/Wmf3u8LdhKsWKCAyvRZJSGzMJDszN/M81AsFlvpbTnwNxXzJ9QKTUPVDRUuc+ywwfc3
f1vR6gQjzlF2WaoU0zB+k3Dcon0lJ+5dU6fnzQVaL846KAE0Q7t68DwvIJh6hXWLzVrMGiL/fdLH
Eg1l6qW0QsXoOeAbE8wKynpm2CQnQuMVq2eGalvc7Yaq9h9iwVtK4uzHa0dfUKPUvWjdLEZYYwbJ
doQEgzD4me4AYkR9MXBGhHgRjI9q4IJ27uvAfOq7PxH37b9vLb22Lm71hrhhaq/bB/HjcyObWawr
BpwkOCQncY409h6DdX7t1B2HnPFDUT5GOl23xhMPPjlzlqKjOeH2Lfxdx9PVs08hDVp/MbAlckpj
J7m1jrx9nktMAt/Vu5iJty5tG7/GsHeiZqWuPjUz69mqSCLfFcv9M6Iud1HFja0FgotS3JwXzrIR
OkE/W3dCuWibiS5clGcfLK2W8atSTXLGBuuC9ZtDX6JLujTa4EHTX72t1d5ILhd1ZVa0HIpmqitr
tA3vO6fNVGqzwT6LZBzemFTwtwjUlBKj4RBt+P3j90Aa0dPLXEcEW21/mn8u2WhB8e8RVbWDoxzC
dPFa0MTyAQmQnRNKgdrcdiHAJMk2Z9LXPcEFpxNA3vUiIj//gsIlhpA/4TkbTw3ALdF96CMknoxj
Vic2t1O2U0m6lodT0iDhz81z3tnGNASDl0sDFTbP9pmahIJhvpF/aV7g+Drjt64JglaehoxZ/K55
9ICMdhuaJxSCYWYoK+ua5zohcFJeX6GdGwULvySNXnTah/391R/EYbwHqjnUe+7KeQGX8DvUk8oS
RVGJ9Q7M7Qxqn3BVb6j/KF5UY2oVLCNz/lngUfuFOeL1JTpqrLK8OcKcr0pp9tRx29DdmpctD2hb
T+zJcb9OV8/nivO0uhbkMxY7okaLK99JV7WWwJeg3tnSZ94G12WSnrfYoHHgCzC1z1a5yDj2aWAZ
3+5IYKx2Nh4otBz7ojI/h6HJhb/ekY2L072iEGMErFtPZjfRThEoH7Y6DGSDPBLiyq3Q4hjnVnZ+
4jRuocfnCI6GUO7w1X+mXXdu8OfnWjoh2KDFFd8rcHRLlNQzyeA3bYBpAViRZKmjtvnJqB/7xv8r
tRnuDwgZ7pvfNLLSrIqw6P7SnoguUOg8lL1uK15uSfVtsPy+aOnNvm2nCxqz/cqXKUyaQ2ljWSOb
Yy+JpW5DsRvHhBVjlYBM4Oa5trHTlpqchWZA8GkSEXGzCk/Xncdvn5Kqw79AnkZlKreiZHnf9WFC
JeCvuiBmkv9tVc219dweGI+ItQC9vhtPZclTXcXijBFO2nbOxpSbRncQRckP1b6rmTMlnByY4ypH
uiIKQQW15mlLvl7yTEO9r1HVaALtmN0rk5KE8uupkLEXHle6NJAewgly6AHUd3XZfTdnneCGtIGS
tJHU7T6dyYZmaU29OkiOR3UWKdS+laXE+7RSB4fYW/JeSrVpA6PgXhF3ym19d85LZH34kpAF0OVC
QiTXOkMaMWbQXMQl+TEfL6azI+TGrDU85hWO1qWhpdjEXYvIxZ6wcMhXaesF6DnqktoET3G//kAe
e18w0jMboIB5ZUrA+geXd/tGhLP/3jIbDNP1WeP840uiP4ua1Dl7mWAJXeoK/AaL9Yu52qk3l8Kt
vTBobasDq/Wys/lOJzyatDjBXaq1JuicNX1Sh3l+YPJeJcmF/Y+sVxhzjwovB/pQoJiOt5M4O1mp
x/aKF5RVjuHX0Mkszx0aTUrAQ8BzGZAZtbqj6QNp4uRS9uKkrix1F4qBBqRvwTzSWig9aEddkC4J
y1U+3oWO95nxwDdZlDknJJeL2T7IiDwp+gNDCegc6jaDGU6MyQZAGm0sEs4Q2qczf+3kPajEKBNx
YpqsMfBgizNE9Uf2I636AKLt2MIX8xbAxjpq+hJQaZoRk/LH5qmAT1ME7UMpQTqPeZjdX1yaVVcz
A23e6lwuDNIjMUdvm5GLvq18LIYTpp3xfW8zX8HTon0X42L+7At49+6tjN1nMrInQPZqDwwM8+j2
0kXe+SuRfzcCWDZioACKM8gdiMT7I8q6iJ2l2hBxzt4b3bHwimbRjPcU7c6mkbhlEBPBzrFKrXHI
SrIPJtOf6z/IRgrvoAi0GxVrnmBXiwTiX7Ad1sUjkwPJtN1DEVRZryUegY14NPGueJ7bJ3zrbjon
+2hTCrt7eq/Rz5I3G3RjoxSFQiR7xD5M5PIC4s9LGacJzyWF1f9DX1NsPU5YKcctJZgy4QVU+Ww/
lgnTlJXCvLeagaeCB+9K/NItmNoYhZDdd8KmXadn/wZQ84rcoK7VEOoXCiovUmNf4UVayxdcAZpV
olytbDa+Z2qxnTytPZdFUdxjpRIWGk7Ui+2wEw1IeIz3Rrv6gM7xpICRRdNfk69Q6KnnBOBbU/d+
/hns0cXM+AP4YqexN78fYsCzTfAU7Uwci2TQxGBG3kpYKzxiEoG9FKKAEncb0JydYe7bmQ2Ctgix
hLrR3GJRmYZi+MtJGGjLrfp7Ez7HLabzukCq4E4tET4qE5F9WEdMZ+Uc3g1mchmzth2vdnwJFCKr
nH/kljCYXoqmoYDUHdVaFNyxBMoRlumh9sxTfJWamzz9tDd03/sRG8Rp8PmtbjgLybIfmNIJxHku
2MlLKW5J7gnWo4voY/Rtr9F0+xD++eQwHBBtrRnMqXA0/YJ1ByEEe5cJAO0I2LhRXMGLPIePw/cp
Zkw6DuWzb8ZcsPla4CL4zJtviFXHjRlV3/Onnx2m8xQU1Lw4I3kVogxz1ewMq3LZbqggYy1CA/pr
9KpNuAEDAm7/JC0wF3mgSKVDCDYFNk77ORuWnXMTm9pZG7kCTGp+rc9OuGVYGpSpvUCnvGyPYS9J
IBn0wTNkBirfAR3TcECGOKpcHbw0N/VTeTuhw/fhuWGY0LUDP/5m6vrAM+AqiAnoKhy5qrQGyoW+
HabyRRPp2MHHoSCn48h244NyBGSmPB83LX61ZMbaujW45R9qr3XRFWwVd0XHwDed1y9Dyb5SraBl
dHKUP9oyuyCVgu11JmLcAjNeg4z9R32tN74N3Lee3QAeE7I8Bj+/S6FHoSusu1PrR9kzhqdbv3K1
NpcUheX84MjbIFgu2SYZH+wHwIA0egUb8UoEQ2q0YYUvVe5pO8Dr60boTvhXETKTEhmA71jS4uu3
niNaKBXnzZjbRt3tRTN9VqsW2FUGYllIduIQPJFC6ED/ih11XWTjGs/oEBNxpabhMJUjHE1DPdxd
g2BMMK3Tm0kg6b2QsuD4svhHPh33NCQK5BYI6rCzOdDyC1C6WzvJZeHYtg5O10/ELD0FMzozaokK
TGMJsUyG06By3i6iKci+jFOi29Wf8/rD4mijrT0Lm3+T5m2ZM+qpMQWp3P5xZUZkvrcN6cmEpMID
baPOaW7EpRyVbqFHE7dHnJkStJ8NGjs8YQOaNHuXdyZGNJh66WCLGGtNvdnTCMRdIyyfZF/KXrpt
tUmK35xGiHjAeaXXVKGMfVYWLvqo1Ziz1ZPL9WXPJfd+4QH1dOrJ4p4qOjZ6XLlelFtaa59yodXG
2fSSGFOFwCIzPWEqX36DtQyd/crjJNLRqk+lBalnTppZbCSzfb4Fq1gWGCrGWn/UtBrtgJX/fJK4
yI7H7t93TFnpEEqIdEXba3vS939ykvGt4Sixz/po0BjpajZ9oxp6ehzgBLAOJnbQo9oylxHOiPFP
awoj7+ujOC4Eyq4YOChr8xCm49ohCHsJan28jqEnxrrMe9XkGEyW0RF0SxL46x8x42K+g/WYSoU3
kXQSdc23PihbV9e1pIZKRNo0Q0/NixgNLaBwIA3py+jmqWYETh5FDQRgpnZbyUdTTAvjez31FHxp
/19vGcaENy3zFvZKVL4AGPtNMlFoJeEa/O3IEcbSAkCLtOCT3klthWMGSN0BO6KlqO6KqNT8IFHT
mJ7/fKbkBRy31fUKoHcaZE8fXVAF+1CDI7yLO6mS/rWqngvlX1bLfYvnhSliZfDNyCWnqIJpR2Ad
IyhHgcff40z+/c944TwK1NnfkFBm9Bnkl8tSn/Ci3fsF914MEUCV3Jj0lAOkEsYtMMRGuegmOOd8
rUdFTXmzn2dBy9y1X76gaAZoUVsqkW5FNj4YCYiFmyzF7Ni4aLz7fpyOTIkaYeiI3TDMEAq9jRjM
TafGT8Ul3sERAVXmbnGfJ2PuvDZgaOFPcBsqj/4lSF8AF/Zp/mCJ15RuYTou011G0tGxyzu6uMBk
DqugQ6FEcbeDqBYHTWgveUgdAQoEgRZP2/NqvvrDmdmCGpG7OMaKAqIqjWdMrKqLEDd67Oe2AcYF
ppaYc+vyusbZm/9HbSFF8Q/UVwh0b47IryQMfsaV5D4e1nF3DJ0YEqGOvv4khvpCmKFwYfc6hqDP
qYgdTvT2KKlVx3I/ch793cj1xNvgfMtQdBhqbU2+I5HMYX2BEsX3vXqSOm40q4+dXRARzOjKfRNp
u1l0c6+EoJNx818Prziejd+53IK6Qk1c5DmXQiOaeO+cPLwo/lqyUpcaKMj+9RWz8P317an/iwWT
NKzdSkeogJvNGpL+Mf2Bk6Z6iVPkUIizdafuqzU3UWJgxLTT6m4d9n2c0JaiEVLr0K1S1EG9PKVO
VNkipM0tYbqFLHsDvuOsi26pn6zBbyrqMZqw6tSOXEb1Q/x8Xt3NZwyiiv9aBRsMLMAiaedfetV6
ZNnGS/nksuLa7BgZxfZscvRSIbUwVRIjfMggVQXPabrMWsozuFj3eSsouxDddHuR34M6SYWv1Crd
4i6Icx1MIfSV+PV/v/q6uVa6cyZpBgEMadKGIHfoUysi1BEKRPY+l2GYmweoLajbbiB84E/oCvRD
bw9PSo+htl65uFr4MVDjhejgFIjgVBG3JwA3nuWGISxYfJ3i083JkzDITZKPgr2paQPj1e5+ECc9
JsG0XJapFkrPcNB+0AI7YQy35+Z7E51PMHJg7MYoFgESHI4ezTE1MKroha+i7EuRhNE0dZkoa6pP
zIPC69BthDD2TV3eq8rfUA6tO/ZSMuDQ5NSfEIa1+zo0IE5FR9M0XFaIznLRBL4tyBaQ7bgXktOv
Y85dTes0haRFsZf5S5K2K12fFAP5OC8Pat+KU1zgcg7HqGPoQ3maq1rbwGSiZSiMPapmAwxa+R/x
SQ1czp3OglKsMPFVB+rT8qsyxUy6w3zX4SS4Wnt6cAGW5w1P87zgE+TE6swg1a6y6DFV64xWypcX
ovJnltqL4uLxgN78R994S5ZpN7iYFcgE8TpOOtZfoLsbIS7yRSMacelCxqbKNuy7v7nD5MQSLX52
R6GeNj7T0/koZ6pMUJBz9H3f4OOT50heaG7297zKtbuhdIH5itkXZtPTfF+qMYmzes9K4t0kWL+c
pQGHv961weJrV+19KmqebVoq+lnPjiXz4flDCo4/xTqRVOPvCgKyvDPr8CsJzgB1KPcNMgLGWLlT
rgLP+YelpavTqLtkyoMDByeAfbfwdshYVey2tF+F+d7H2UrCMe9QSWaRuacDtmeDlCgdYUvlKU2R
5m2ucRm510j9Mt9bPF0Ds7elkExoB9K2D0cTGZODS9BqX36q/YaHEtqOixrqErP2/B3TjRVJt+oP
oiU+qPkggXAKHycm0GrURtxstOmrVFEwpYiQebHFMqZ00qMDyNy9Xn2VmYnIFL14ZkLgxQLh4S96
Z0KAyruNBSe3qpHMVpMQf6JNpLr/2T5+jbxJ/YUzikmW1bLYKRjIELFFOHGMvsLHgnqxDD9mB8RS
v8BmUOQFsfWvTx2RTelyl6piqFuEyIOe9QCGZIx3MTnzVoy7SBGOna3tqf/wBWU7DdbynKZV4Kow
jfII1eQb3K1B17Rjc6aDx/yzbnXtgfPBSrhb2oejMLSYex3M71C22i1VsmxqGrVfmR3XtIFfD0cw
NbC4scKGJuC27rr+Ncr8iwq5Wi/w7IfVSm8h2ktau2xg8bH4eIESFqXK3cil67lJn3DGo/M7mGSW
dFC2oDctd29mRNAYQDxO1oY1t44mKMqFXHgZUvV95oUbXuuHR5NPOwEzWyPIEcDsKDindHbuxtXy
qeQXu8P2nnS+tZgd/XsRep2y5XBQH98kD85nL0Ze3lER+pfQbEx5Q9ZeKK7OGsi2qaf7WcUhgcyd
vNHM5eahmYMdhFGww+hGz21hFdO3tszmOQKzOSE0HC3aE6cvXGxUBYVGFs7g7cgHOPN5ICIg/xqj
zol9IQOdjM+BsyIKuOrN4VzQI22iG/Idd1guhqkQGTX0cGsLDW7IPCasJ+dHq7GQADHtloTrTLEi
ZQbUQEoW/lOE1a1l8bsoAU/A4a9nhVpQ3cyE41LouACjjjlLjR63nG37Y00g8/TV32f3g/nCD5ki
/V+oddgPds0i5bLdCylLdgroru/BFHSk6YH7plnbx28rxfD9R6fwt5Xql+vmPzAVa+G1zDoHLVtb
oXKqlSP603qv7Uk5LhaLtiWbDEbcCOh/AgqsR4vRku40vUfnlCy3hwCsIue7agUznErXR1JbXW4J
Rw/b2goGAPwoyI2KjaTjFfzZ49L5K3sEyVAXd+tFkqjZ6GZJPdS7RkM/sQTTGkNzV3VA8oGiuaic
l1WDeIZluOVU2lY3Mu9g1zctXb69oQSjIWKzzrEL/CBcD0urJEyZzRsn3QST8BHvjTk99+6UAMUz
z9Y3XQUrcQ2DungPv+lAzCYNnrrxra0JY6S0wLYAFHOpsvruj9GavsaNeAcc9m0Rucb/8XNkpmaU
9t9QsesNAYxHGbSQHDsW/hXV2g5ZKvUxuuVX0Jhpyq4VTI6GRyGu1EWGxalTmLG14J5drdnCSE0f
+PG63ffEbr64ZiuvKLWqBFVlQz73TaDPgjZmI98PgFpI73/BAb76ttNeqN2rOI6xLyU59Mhz9J+D
VR1A2WFrBvTcBojVU6JQsVhN1GeVuk11gawcudvVUa6Yu5NQ+1MqILuHgZeKsbZUf5xtrZZurXnb
RfKW1MiEPaSqCttbLvORxFVFdMKKp8i4jowziR7bV0SIVXM60JF1XFbOwmjrFkzDNybtz6UE1M+c
ZGs/guo0zcHtJxpBZZRDTlBjbL/Wfr9YBZF1ZAJ1hYStm7CQKn3qk0oHIlKwfQKEyoAuNKU4RY9w
ZBM5PwJe6052L5BB3y5vwkrik9OXfyGmuxj89H4Xu0R9d6Yus9FtY9k+p2yqD7WHmS7X/A5d3cpn
LIa/NWTekQDXuEoSUv8kOr6bi/RfovdQpDleEYhNmQk321bt4GDU/yp1CisQltVYyebfRuz7cp6j
YEV0/+Eh4XhW9edNiXHK5WMRfFIb/3GJdQlwTP0o36WSpAAA71bj1xNOdog6ji65E+9fGOC3UlQd
DfYSL0klTUTbmC/nBj6cngTSYzxG77ni9TpqJBiW62g7TSm+0O8CaEd/fni6x2JJoPzkHm9gmDv9
UVx4I8BFfmC+VfOiLnOGR7qsxxAup7aXxfudYcl/FvFnjGnS69FwQgdHqOwdN2fzFTezStU3cmWi
zSzSwV1293zYh1ASESmi7MPO4/4fjJweSYjF6cBH49ynhJlv4Yb8IF7ZI0oe04onT84n1Cfal8Pl
bJivrtUVomdKHkS2eQoDpZW9yoIotXVw9NSuUK1GKKMDm10FLjqajEbn/SpnIH74qHWiUK4WhVM0
O30ytMuhqxeyWoUFvVyE/tsSRKY/N3rM8uzRxDZ/gGnt2or2+HRRZMcntN714Y4lz9vKrbpf6KiR
2ZmKNP7Cmvyr2HwOq+ii24EI5fdk9egt0p54GnEgIRx4mpqe9fbTvoh/moFl7Dcum5UbueasgnyI
UaZrFwq98ym/0ScMpQ+yoDJNpFbZ6/T20xD+z497Qe91lSEdAc0k4g/Jf/HdQkUxyJdxMO01djHE
OVCDMqkf1IQpTBCUe2my/347UMxnd/fH032ffzA1JALBjYV1AoylN8c0FaXuzOllDVtZo7mcAxZ0
wlkS+kE99eIRRui7IhQ5dmYFoSx5Voxpdv9lHLabbJNiUZQcodZY6/gzuX5sWb8IP919E602D545
yLrG7FF1FrOuSUNK3kAv33IUFxKLoTFQIh60hhgG9WvF/T+ZwqX15Dg6wEutyRLuHTGpEFRtUwoY
elvsvVMIPGIwuIeTv8p314J/AoivpYwCEvBpdGseNVRbRKURMqg88b6QVvLrqDG90NuvbMDqiDpB
HyRvTfSJdfr6dMelNl4dIHh2UYZhrtaDVEOWH19r+zyrXgdEzSq+8kXNafq21S3S2TX72jwj7AX+
HZozdf74HIhMyewbvkvGKnqY1GpuNhuRNlnL8h8GngLLO/E6k9dxvG4CABdziITiv1/J5FwiQ/pi
5tZS02DbUoK1IJhqGzDjscEoIKoSyq9gWNEIK/eNgZtPSNtmHPyt0ZBvHsGr7bjjYH7VeZRW2n//
QKuNJer+k3ABydTPZaYaSyF6wOq0z3RFfk8iz4WFk6Ri4yy3Bq021NEkbFXGey9eBCar/m9k5VMM
+WrllmnEUc+sAdYceo34F2wDQ+YIc87L2yTerVbLwGq9c6LWW9Uo0SkjQ3x6dm4UeF1nzMWIPNDC
QgZhjD/CpS2xSxo+spCj+uqKNnnKY2dGCUkTHcnGxCwsms8gSFrPZhk7QU4A+dM3R355y4cCymZq
i67SytlBI/o1yoaO+b0FPd1MqIIJVr+yoGfVkE/9ls2KgYJ5PK/1KQX5g049m2SC9rqpJmw7yIEp
sPkf+2SOxZOYy10InWYC5+lWNyuT2HOn0N+QpbBbgexfFI4zN8fCXvFU67bCXAt734GdArRiWN0a
FZF+/qaodNn7EmOWcTuIEuC0J5P/itnFLYTyU/LpYgDcYo1bkQeqmtzKWBilB/bMuhabFl+7mwWl
d8N8tyZuH6cumEOG2TsAjkrrcFPpmccKJmS0HXIEw9tC/olvDm4UcwDqt9HQIOzLh2j3OA4chD7u
aLQYwfqI6h6yvJdF4SESwcjafKYt5LZc2YwATpmhHLrZANR6+4dBj+gzC/2FeIOEgpY3nSWlHi2R
4IPuAxoHcKmq9VywgV58xP/RWbVH33QpB2DlHOa6AbhwSr5SF9jDm+LBjqB2kG1wj6gY6qYUwjmh
Kfqnzq4lrQ3picFvSGH/Zsd3/SeJlcHFeZxom2F0uj+HZpa73hEMNjLOfaTC9TWTKQ9EjkcQBrKv
EHZFGOiwY/w1d1mz9gc1kVkD1UoNXOfVTEiSVZ4YzByK/034gsPQ5oT/QYe2IT9Et5r4P5nbiPcF
MJdc18S4avPHlys3Yy8hkMPxwz33DgB9yu0KxTLd1VuA1aGcpyYVU+37ff+s26KRDc3B8z/Ut7zf
1L11TqaF2RHCR+LLKbWjP1FRBWePmATuYPsgn1nQhkw0ymV1dJIzvxvaN18wBTaR44X90eybbfwI
vNqyQviLtF+uZDV0MpKkqHQJ8EGI4PAHw2XxxEsu6EKrJQkIP29cMgz0D3oeEijl8Hy1+N1Eudld
W2TfPd1fc+IZ/0AfyqtgYxhsQBMFYQba1DX7o97CVYOX3MEQoLoHI3y/qxyhN4FOU6qZvZ+Y4l12
UoTv63uaPU131FuF2kzui5cOWhf/EMA0LnCGjgQ8oLGJa/P3ie4xBDasD94XHfRTy6tacI7TdM+3
qXMFplo/CLV4pRP27yI9oFfnRzM6oSCMeQA5H8+MdmYuLbf8Ey/eQvVAOHtFSHOJDEOu8PReCWIf
vrfSf3LnRUeMoC3ae8CjZCn77siCPbuEXa5R7HASpWM+bnLMVuiqkUDHGeXCELcSLGrw5t2WHNNV
E5tdMWcNmfAGQQrmBFizKrPnBL2N0NYVebaNjMC0xofksQWWJoNpMPvdegEvPDl9T1t1MFqW4Y1V
x3fbAdAZ4beYy2MbtlQrgE4HtauHy1a4MLfaOufVHtk5wHK7YXc94zLODyDzxaWaMgwpPSC4hjJA
Rl5YDf17rvyQvlhu4k4m+2Tdx2bWlZuEYcz+KDnuKNL8B/NCRhCto0lcOfBGbIMV2SdKRmxWMwIf
QfQyoL+rH+p/r5HqHYKfja8+7kWiup346hXn4Qe2lDZfSGAfPRHPgq2LlJ4DaInbZPE8JDpSN1CZ
yST/fwow0Gi9De+UGLtDhs9gP55+RGYTOWxRhgJN4oYYOi+klCCVSal2uLQBaUkfHmBmrRobukzT
7Xp0rzgurA/+Iry0u52vZWMRzSSc7pmTMl+o6vLEvsedXJgRPvidWrv1w4eFQML0dRRgzTFjVg8u
ZZp8vIb/ebsUkwZ2BZeuzpZjP26KWjhD/XErVKV6sPpikvyqVACXS52tjYw3A5QVJnCF6WOPlQkP
c5zvKE3TrRntKGft2ct/4NQxEfc1ztWs7SH5Y+u6ATq1FDH6NIbdtN5hTmtibtHET69mzzvVb+Ar
jNHAmPwpzMpXm1ynH2QPnzQrbrAQK41yN4aAE5Br7/qi778Dfp7BYJprlUfz8ONyHW/dhb2AxGfP
E8gCn1+OIyWIfR+ap3G09RyQNyXDFxucqw4Q16ISfjuKp/auEM7vHtd5UJyUxwipYwrYCwt0jK3O
blJMyRerXXr7IGSeiJ1ZCL3DBlTcY5cBb6qQgw9N7Z8l2VhNcHx6c2TZ22D/o7l7difhtz5hDH58
a066Zpurow4oQvOi8LIY4GLP3gwteEamfUYn1vb/a8xuvh5TzDdCqEcCnOnGsEfjbTL12GvqosES
3VVcaqDNIIThJLDCvccaSWnw1O2SaIVTTKwPRjvZlci0av2peHmklm+lP1xH7KGuX5srYrtXDzMh
9V5tEs8vfEHBWN2nwIJLxgIBkWyNUCWQ+/hHj70LomShF7dI+00ZgQObJQoIuV/uTvcRjMI09JBr
5xkJ7wtV5leEN4Q8sGFl+ZRRnw3uS7CleAg+5TjdXPFxR7T/zuhU+kwgVd+Xh4T+MRMrFcIGlqIw
dkRBNEEBOuhqIU+n//nl0Uk907gBFvLVpj7tyihjdwi57lbjHBTTyRxvMQ2ZxpnNu8U68N/7czqY
bk6FfNch4q5ki+xXJqsInlYL6CbJ4vvbFFOnxVX/DyR0AxIqjmwuvFO0JHY5co78+39+HcV6j+Ez
BIHUafNx3ZDyGXHG6C8uuwJhXwGKZVuyxKtUkBjDTJXM5kTnLGJuoshhGsipjnnLidqo9oyXKKGx
G4repTFAZIcFsWQvXrmwe+r/YEhUcyk3nBESAnTtGjdplaru8RYYCXCvcd+4KYYlcFeU8dGb3VoR
h3LUYdF9U2FddW0cCUreABDRL8x8ucoZ0YQb/pOHO+Mcw82fA7EOB0QP0oQcEcVFp3yOxdR1XE0S
2dNSzGl7thhd3OxIAts/SPJHq5C8h/agf0wM9SidH5ks0Y4EWGuK6Kl/z4RL63wBBUz8RFXRxkLm
5HCnKiW8jNTF1TVVK27+hh5InsizryItqUpNv93Bws7INecCTip2reVkKRbsHVZUCJ2RZ/0Ssg5i
xnkQ9GFhFvr2Yehu9J4f51he6+kMZD2DE11lQgGTDvWAFvuE+m/RY9Ri7BrWNNextE5ApYQ/FWFu
g5UKeY7G/w568v8slepdrDwTDn896rgX5WbA6SbcDyh59e0HT57DzfcFujoXXR65pNM4AnY73W6Q
U7fBkqPOf0Y4MlRR3MxZ67dxbA0bJnZH+mq9KaL7vUuHQMApxOJRn0Sn9AFxd7z9m6aonnPl6oe5
fGNQelu/uTJWO1ymyhiY6b3/Sg+DrwwTIsCtoFtRYuQ66YBqDigOPhn8AHKPfSD8w5+KvYDO+Vow
0uOOdei7BQB/3b+9DLANkwETQnnEYwUHS5ZTF+Vi/Nwl4gfAt3FF5hfkTBdcvgtXEENES+LpVoCg
jP6Xc5/i7nZ8l3TO574zOB2j71UAaTtBAHVN16s8YGdENYM6I0tjCZsHAHh7zYat/lP907W8HDgl
MRuQ6OKlS80hiskDJaIMRMFMYaEtE/h5StPMzoeKOMAjNUp0TnPDARvFMWuvLLh/b+2qLPGI8Mw4
0VZRJSjf1xi5pXLjeOEYFo+prQ64HrzWFqf6pHRoucKH2nlbICjliGt0izA3F4UTrJMt2iYU0dLl
CEGVirWCKi4CcD4uuj/Yz8MFvYGXAQpHWyHQQfFxe1kk64F8CfiwF5e+TavM1oQypqP0ZoWE2TGD
9/t596O9Mf5goimb5AdouC0vJnqjbTS6ugJsSR2GXd64PPWba2xoaFI7/JHBeVP2lef/AyQDT6Z4
Qq/CyuNI4YVgKP4qdRLSu6gRk14/r45rDGLGr4f2I+eG9liJLkVQ3NV4lAdRfedsK6MxFeK6wUNf
MpL2zMt+uGa/p4dMhsPOozo3k/DcfieUHEOoV4XytYb5H+d2kzH5ypHcB6abpwZhqCGRV1XAlXt1
jCVNP1EElgcLQRc0LDta1L/5oMelqcWzj99eCNB/r0z4KUecGmzv//NaPId9K9k1jkwCC8NMe2bY
vq/yVaPOzNiG3zkuc88vEgsW6pZArV0Xn8chliVOmWOXSmfgWc1kwM1LQ3DNduLK6Wlk4ZRy8OLj
Yu0NUFdQK4iivHgXcPhBfC5sl0ecX4+/9zrCPnxUs/KtluHezlR+ecd03wHuCvnFQ/PvP6sLqA2d
JcfUAgNiBxGn+wHy7OEtcBwZnlAWlLiUj3QxuLmfm/p65F76qx0TTW9PgrB0ZJhwVHnM+0iGuABK
3j7tEE07AsB2wZyV8vZA+ZTeok4i2vCNDcTMnuArk0GwCad21macELi4/idJo0d9CzY9lpRREQJQ
A/EjCDBLT25MT8F/TMsGWTLsoHTwwdmaHJ87bEog+OCCwmuSh+Ns3mw+MO8ZHknn+4Rsky9ZGzn0
LlhsQDRr9iDuv/OGbVpNZUOd7SRP4AACDj3OVNtyoQoTak83bp17EgkU6Td91wjdxRwwY2VDODKX
ZgNTpmh5JmtD4NBB6/CGjulTTxsZnlBavE4UTvXoaihuIVY66TkzfANfcppGBF7+WhZjhg+r+V+J
hePR2tuLAQ+qXsTi3/xCwx1K1NHyabGSY7mXII3o7ri2ldwSE0abHqHKkWEdKi2TX9SR7C6cnRHU
15pLGPeoc6LbsK3UZKze49dLFQWfX/2xuzreBUBs11nxosOwhw7GYoZ93yaxoyez882lKDXjhBZJ
b8ZO1PRxxY+fmRdbnb0NS6t/7kIZgp54Dz7P2+89xyjYqs03qyGcLb7Xzg8qUu+GZMskEYh0c4QZ
6GtKXaHt7qN7NiWFPBdvtmFOnmz0bFTekDhIni8jIBugeZgkuXngvJs48q+xmsXIyzwSa+hYhn98
1fKiOte5H5azMGfO1AUySkr0teAVuFbOxIRf4On9SfV0F7kZNldi+1+FvPn3CJagK7wyj275/fqL
4dWIF1EWP4Bj7MrRA31VHYyWxm4qiXl0/qVNJcsHE63Zl9gBEEthOBLEpwCCzvHmhD7qOVRpHRfw
etWVI7Og++OfIb1UkOTUoosAbbuSTyxhmSHDZ2DQ/rORVJn/QFHk3BR38zxHRtOsNSUXelgRWGHw
Ob4BLzi5FtSLYFMdsS3xBIwvzNLFtfuHi5ZbO+8i+6LoYUm9lRa0YmVJvCUpDr09f72XOXEWi1AE
lefIIzh7Z9OtnX6o3dH1VkdL7vlG8p3DYFQ9kyX3DKKXxDy5V766HrlhQWFatkhn5ORPJTe1WZWF
BV81ipDz3p5Sv0alTsDiYey3kXd/l5gX33vHN+33DmmJMj26EJJ94gMcYF3aZ4wOUQlnmeyCNPiQ
kvTbX0Jm74WQiGqXXivV2ObcJCc3LiESNXmI9erRHQnWV2GG1O4NauqczH3Ijrk4QFKIZmuGp4vY
6Os4TNSupUjSZYnGzx98LwhjazEFXNjbvhsQqBBjHCNzqKmihDNesKU7beoMbTlKJ3HHKznmSh8d
/pbYVkP3zk7bt91ue3DjLg81mDoNv6NPTW33RHqlb9P4MDHDX7hgpMJ+EgSpkgHkz6HjMfqUdxwJ
JaTzLiU+XVZMNXN7tnjfEQ3sGEHKXoIk+rxPetcSFa5DWwCYlfBGxm0vRSfCI9yHutNtcBiBmwHI
sCyIspmESsr3CA7a1p9J+AyJ3JT8Mq9zB8Dku3WTZ+l08WcPsgDk4gdt2+LBnw4QAhGrVxbll0+O
NkQPeuCxn32rI3dfMvDHn/edrPlS1MtpvNpfvh/n5cWIrQtWTiNxW6bmMPAKuR2reobdBfTYAfPS
Uf0pPcqWfpGeTtWWQbw2TWaEC8/BcxZtHfpmc8aR6fwmokXiIUR6PWDKr4/Mwc176IbuK/aE6cK0
it59wUrUjgIdjbs3RmKkG1h/1m+wrXnMvk7ZzPY+xeNunXtCpS+BCrYvw0qS5MeKvd/ZpgHBKMdE
koDY8pVd+xg+qxZMkrlvcS0Xbe0LwtMqUq8ich1ta/yXs1oQObkzZ/C3TaU7UCs+FvzDqnEIszUE
3/M8ONqtAZsoanG6i46avdm9qOOQmjMHdCFZ5ulYXwBqpUVFXjDiu33L7pe48tN10v7v5DUtZnUM
qt3ej0ubcGiGBSZ2VYju0krnxppRDhloA+Oxww00eT9ihqpqHtZPetYH3E8RH86tT7vfGWGxk8m8
jvmAl2oMIuHCsToXOxvlihLMiZl4KSzF7B/3Vbe1kbAf+Uh3vEc7qB1GoFsb1fCjoEe2DPq6bRSX
Qy+agAumriGk6KSzG25rOlRBtSER6wrR7qZoZ8azoiUGSVET3IvJ9fQG60PjM3czHQ4QanQNG5bC
aOBj7NLqtpNvvzKnXXqHy/qqA6InGRlfQ8XvYhjdlADhygrrNOrRDBHXq7/QoqmA7OKpb2t/Wvc3
sykjMId6f/kljNRMm2vbDVd7vBNjomkHpfIPtMi7UGV/7ukP9gYIsSss+D3drfI65ncsit/PVg2O
ybTNf+4GMYjzPkxWSJF7JnRpwYc5lxUgiY/Jk29VGFsK65Wgjo9u+pIxkJZ5rRI5coXLmK88/ThH
BFPBv0pAVyy8l+oS+F4jFh/A8cmTphyxatcEIxupxBL9vS3pkJLCMj1iYDol8MM6dNtdfSN3pwCG
xBFoDHdazE4EkEuE6LL2jMdFijIdIWDalcgMXEzkaHd5TenDdpNQfzrgA09zK+l69EhJgqEBrkGA
YxR8gHxpaTMFrIS6rYn/zyOxNvDyWqYN//HJ0Auepl87s/LWN5UjYgZM5woz7ANsb3htVXLoOOcP
7ShkC2L0QgeVR2VDht8IlrwGUDZpaxERtDKoXYn68LQIWoIWvUOBgnwO0TufKSsgGs8edVohFXhg
PwWedoSi+njuY1HZEBoq4w4kO+Z3HWtZ/7KCcS2lBzXC7p4LnbgDpPTBnwuSALIJrhjbqedyntWa
J/eJyRy1+SsvAgPtisMYv8cxLJyCbhqN2SHOOi+hHfEptf8HXAPaPrWQxCZkUBDI3ttL0iRbUjcI
ychEI7a+Yl3s3Lyths0qUpX7b03hbxirRpMalmT/WNciOY8XBzMn+PsxoCRMI9IySCynLJ6pxdIh
WRCt6nLsKn/iYutQnDtD4fJfmGhzElFiedzi0LB81l+n9p99SVxe0b61z+uIOZWo1JDcmz4lvx14
bWYV64UTFsiWI+Aqhiw3EkBc6Wb1ZoCZfR5dCKYcpqDSisL+QTgoG8QsCmgQVUYpmO06GTNNVXsq
P7u3e5FqCmIzYto+hRZ53C2P4E/iNdF9m10rqdOGHk/KI4/6FopxU68afFZGSFK6qgVlOqhdmmo9
sEamb5tamTxP2uw5Dj6zYOJhublc6oIdpzHy7MtVKfyiH+XVSO49RDt/Xib5G9D8Zj6dikEL+KU3
DZvZMR6MQq4ko8Fxpb5JSWkMLO6qHS1PYfmVeBECv214+pSubzZH7Kz3C112Yhbw3XHgleQbY7Dx
e3jgj0P/xxTt5flcauYmVCVXg3bCHYwdUtp6/hhz7Fa/4r/JFVqy/7RM1V+vhBYqPvw3EhKvntxt
FzUKvER7SRtsX83a6ZTog9I0i2WtvaJSQt4V9V3Jg4UROlumEOcIvellNqgxosm3G2tQ+XSyu15r
L9ETaFS2P7VT/jIM9sBgjA+gMqq/4KKNjv/TKlorfm7yJmgaD2ShH8SKLjVc9ab4HImAx7K7GI8h
sMmYQm0EXOCgDgTEVWGqbmOZGi1KgfhmAQKJT5lQio9NPrvW3Mpn3L+z2Fhpy3sapIzPeXKFmHmv
YJcO5JMtfqqwuGKY3jmuKbMUq/88GIHCo3OoUEgvVS05Syz3jPIlaLGy2Q5sdj/r9BLdzHhFaLvd
l+Sr8af+vnfvn3pqmrFMPg4hNFkkcS3LhimtIDQNGFDgFiapT6BqlPN36XWq/XM0iyEuhgUcAWAF
saVedb2zR/CoKa12Pyx2fzg37Rj11MM6FpdtsmHBObJgTG20+6eKYvhSBHr9/WgzTTJcgRe2SYhB
hh2H0mVymmLhbxXB5jAhP4c7HGUzcj5YtkdAVEes+mCVnPhK2ffGdJwPE1A2vKnjQcdo9P7Oyu/s
AqsscjoQzwUYpUDDUdW9CQuXZqebySFBKx49bIHz8uw+iYTZ3Zy+uSdp2kAAj+hIJAhF/i6rBhG7
70WSUkQ6hsgLEcLRp2/W2NXfGLNlklChnB0CrqzyVI+8dw9BZEzfFwFhBSGgvxNvk8XN2IE8AZpf
bWklghz0DbIyNS8OpSkfaq16TyA6IpCQKidWpI0lEsimVd2yihEcR0fNGQLGhUphnMYp0JGR9xqB
hPQIaIWbEAQ3gruVxHG+JEmOa1QBWEpR8EeWpXKWyehy/k2E2NOKPSa0sFGpmGgl9IOmV45owBa4
KNF7ljuc/8q5r0LBDvOSHWXwvx9/lIsCgR4aOpwpW7743cD1E4vvlqqeMQu9bRgaZ4EfFTo7WuSq
VFPfkMAGLXoDs1S54OvBp8P9WVl+SxLcgH8xulW1SjdUHWEk4asFZbkhoILzTjw1KqcYmn6Pq+Xk
72+u5kgDmT6eLlPyv1pX9eYUoogAm2TKsOcGwpxNFpXd3ugma3svNAqHt5cuMpoDNRIFneIpjZYg
j1ecIZr1zrsTY9zyfnHSJqq2D7zHSNVMlCgwCMSAEl0QAejLk8imBNy57VwZ3d7A2pXwv9H4W1n8
hzGh5kT2+6B4RK1wWNhdifK4IIl5bWQuEmc5ZMH4kb2vPKTiFqLor3yPhdvqhPxJlJwnAduZOa5Z
4d0E1HhYuY4NrDYVIY4Y3TV6HWEVdwoW+JLlriqLb2KIddIXIysWIbBujUUnm/+hOB9ZiL6Hp9cB
pizNqqoQBWCdP7CUuaVEggSZlX/3PzVkxFgcDO0BV7GWFqsmwqf4drZgxjK9TarWJPorJ5fv67WA
rl6UHNWBoMsYj0Oa3ydajUTe4wh0xFTfopf/jUXmZp/PgKIGOfX+KwPXHiixHv/bFpy2M9CRO2nC
oyu+y067vmMslkyeBh0zjIg7rP56zVXiJ3+aYt4loydA/7B60K/0OWTbxhelVxT1HoWUd20GVHAt
+GG+dQhJx21/38BH0MWzE33daRPZBMS3/UBxWAKQtPh3eZJo3aVDtuhRBivWwcIhVl4tVoaJFAlA
AYrg6wG4FV+P7wvIHJ/yE9pwZSWwLr7qr6xtrNs1KXvo8hBIgrxfkVLePnMS6UopTdpc1ejeh0jj
LRhzbAm2T1nGii0+ZpU4nCJwmxuYdMUYOMj5VKaxRcGAR+gEzavR3TD/Os4qAdS6Vjqno76hrmZZ
LtqBj3X+bltFi/0+9hzivOLmpPFLGT9HJu46lkkY98fhSz1vAXVPHow02xhl4bt7PI3z6ImDkqqT
ntq9xjlZhYRbsM9xs1y+E1e/v0FbOj+mZmVSt0B7ZfS22iYYKTPj08Gu1LCqCed3d/KW3t3zgnuJ
PiDvL93Uj3DHtaRo0J401jEGjQ1b9TNBkWDSqKE84XmWdjgvvhSu644BTDBAysO9j73gYbbfe2dx
GVz3gSl4NaAI4ZrTfluLxvLoqlEcAjs94ujYVS2gh2ykB0mz/pOyf55Wbr/poB2B7Br2WV3lvkfj
aRDz4Q1FhWkEpfcUXQJ2MeHp/tnaYMB/Wwiy65sR1SUCNiWp4BZYiUUwtQgHrT1Nh9HxysOxQqfS
XcTh5k+tBn80dvpdefmuBLyDKqC1y5hKLJQTvSeu3ekz3lG0bjrW27w5ke5FbfGwJ3sI5SalDpZF
qgt6v1KxyGQhgrsxcuxIngACsUIe/ISJ+TO/V/0jxql3sPg2T3NWtT9IgmMt1KGYC7s6mM6UI41i
1pON/3BocZiqI4Ok2dcuXkwFj3i8GbrvZR4ojaw6iN+Vj20+HwvHrZuW+ZGHHcCJinWY2g4XYAA6
BFERZnLNAZE2juPSuFku9DZLwo4svEjRLW3x/OsAXiSzci/Y0jFKJHGogyvA1yk7kiJgZId+Is2a
coO2p4Kzk5vYOk1VAM/JhkVEMqfPSLP5FD3/D1bZT2gYD+Q02JmyHKIAjlJVR0HMdHZ4oOj1XrQI
94nVHdeDkJYGiHSSkixFa3grNzBqpdADnyrmbbmipz2P8EkzrlNVpPKTN+54/+Qn93JWLmuIPWk4
O3BMg8VHPAEMPp9e2+4kE3dKvxhh97JwX/WhSUQNRREYWOM0IENXnfb3lY5RCpQeAWc1Syffe08Z
NqBpg0ANFckMlqucx0MpX+IhYz8In2uGRycu6D1HK/SdWdozvUbvEj5ExBBaVWNlq98KlF8fwF0y
Km08fZgr372RdYKVpbl2s65vSFNpTF+z+j8dMuzHwL5LDUbjF3V2wiYiSWcVu4ncYd78/XpxfVqP
ADtCMv6Q80o0tB8e7GRqpw8jA2MbwDgN3v2mVO6lU01IkTaKB44NjUt73OT+QqKseWQOKoTE8qcM
gFRv88oDlTOuH4DKKlUnF3+H+4f3yq6XbQMAO4wOIeZ+jMTzjYZ7+hHsQm+O8rSaE4/pjYH86sBq
agik8dLqmBofv4YRO5YIxWI9MyHRH2Cg4ZsO1PVv+WydxDxbSaOEnZICnUew3AgMTsjeo+xG3EJx
f3E6hczCHkw4jfHcwAEDWpOdH+LzoKKybguzmF6oNybAUUxhrAcBW0jcHTC2+1A0sbWj83m5fmSV
wwVauo8fAaa3LsjrD+HLPA02MxZzxTTg5hxnIkE43PNiBuIa2ILSNY9DvQJtbg0tCZuEGYNKrZwZ
NctVYMpKvd47MmTdYtv4YiReCdeeNz4GcylwSpDQyxkWBekkTy0Yexa9s/uXnxo/tVWbNfrwQi4m
4k/OsCPpGmihkcfZ0Lx4fE29MI0/aEQW0On6XeYU+/F5SpajzTKJnNr+Yo1PqTYxck/FMN4nsP5w
1DwagSxouJfe4LoSD4rNZGunhui6X7mrfCnQm2Mqa3N2biSTLHgjPY3mSRgJN72RZEq7gqvqytdT
xZcnuPvRnhgqaP2V422SRwlRVNQjy4gvOJqdBhOP2z/mCBx+R3FLlClpsHANdYEZS6djPRyTWG1z
zWdvZCaOFuVMnNcpwh6eJ69zhUYoP99NvsFPfRwkKaTNFF9/hLw43+G2qfV2RaKK6Ecd4gpHKfO/
fglZHcE8O8+Vvdd8dUdYdFbV0z6Bw+PiVdNXBx3D/SvG2GG01PLpndUndAhhb6QnSK1O4YfSUNgY
yB+TvfejFeFIDLQAjeNhcltu66yCn7gEhqBkv9FCvWKV8F3tuNE3nuds99I7xTRCPSTdFoSBdFW3
iUdWqCBz9GcBdgcJhAVvHk9HAOWCBWir3+/GjDEW35/JWRxJkhm0Kd1pE4rmwJwFqQ/m1G3S07+5
NNQlMewOmDdeweR8bLNd7udfB7eLKyVb8lWIOJWH7Eba1QWJ1/o0r8BsUhefkBhZaFEGsgQCVY4R
9U7ZKYa4jNFNzwVeXansNU/JSDXRzfZK/HDwy+jmKXJ4BYQx9TDSF2Y1u/JunOrcwpM1zUgjNhdu
3O0x7hrlX4sBa+1KMwKrvLQvxrq8QNGTBdle0Vr10fYfAOivBvUT5tWbdT0VH0VdPC2Brpd3MX8a
WpGWYqw5S9rgYeRwEQtRJuwG/jqyB3Mx72xmU6BoDvw968pobUReOvZwkwGBGW4pTIu1mJR35yEb
95zoUqKBkfjnyymMwI8DRSG5HR1HpVoAx10SHHOVUSagBVFtNK+oDumdSxRZ9IbFIyDJ5aeAbOGe
rnz9FzSFzKoZLvaKojLySz6xTYacqVR/o9Fqcni4uDTyKKhydBj04xNlUxQKrwfmrFKODIdCZf4h
voExBIHiZ/w906OB+6SfFHrW+wwWwg+8Yz0iRx+i9LK0O8+GKDP0NPagscW6PiifvkPlxTuTdjxb
Dk9zxjmXPgnCs/ud4GEAqPtE5SmgWNZ5xlbJ277zQTETDs5Dl4qG0XTc2jXj8/rDt7YHuejmjmvG
ceMduXL2zKVmuiMQeYcDy6YSYYcD9JAPZ/F3+98s+V6OaqhznwHvQakf4Dm1iyVRrH4M/DayjtJj
Ci3wMo46Puwz4f52b+jCo9dnDfP8h4z+0EiZJCFCnhJap6gZQ4DW5GmhrlNQDHJGwvjCeTYZjxz4
lTnbIiIarA75YNfGenjpPdz86iGNH8a33jyJK5UT4n4yLIaMHOV5gfczjspqA+JWm6+1yVFfeJCh
h/z0/EBfM8Od28xnA38FGx4KD3HDT2xxRXEga9TQzGJdghoEpab1mca7JbsyoWGE7dpwobiNOU9L
tdh9BUXIhDlbzAtvSM6aLFMJsxjc2d5KJEDkWEu7bolUGoTl9uYcSfE8noO1R18H9ibFuayCQXHW
nUA0UrTb5VgjFGLrYmbthFM0FK3UZFLMc2xUWD+fHLZyfvVyAcgQWfKi/R90TG0FuKhdi95KEX88
hUhzdlV6HavoD9r/Ckz5X1mZbARy9mNeaidrQUX434/aF5M/TuizAXNwEDAH2EWujhmqhgWryASH
vk6rLLHTaBkvzhrRmcv7wW7AxEKsMBxGzxnm5FiVEjrM0V0hMo5P/2CzaguxMZ2tQVzswHBntuvY
Wdjpi7lJD44R55L3OU0UuWgmdrEgbLrZydoAcNOnYdLJHK8V2fpmyaB6r8eiBzrnTJC49RVo9//m
B+I4ChDXyte71zkMniWuO7nmhQFqAebOffVycmr8DzUEMca5pMl5WuCOanhxSFYzdhhV1IYY/rYF
8B10qytoz9htYpcik598GEYL9z4hokwArK0uckQCMdqbXE6EOdJUvLOdpyZI6p/MuMZ7Moxt0PHz
e7UHb3k1+D5l+W5gmZmilFGsQld9XbfIXqnxavTJe692lWMFgm/stEfttWYgWTw4sxlfBP8R9Ush
94yTuxuFqQA/S0x7p/rSMrGBXxZpZJHowziIyc04u+z7u0T5dcEPDpp5evAz/0eU6VOsnV/wdp2R
2f+N80LquPlLGd/OfFW16J1nkWVD6bZoVwliAu4N54a28PSLprXHgHspApNI9nQPs35tsbjS84ah
U9Xd3fbgdf100XMXsJpaQwpmmuau2waMPT/MXgctAbqsM+ygS4A8XOiXLMEqne8iU1lDN+sqoXHW
dztADF4JNN8f5lSDyFMeMUyNX2lU0Ia/FaVu7zuKppSIiQjkT2QiTAmeocqmWfIe0zQjSBskM0Mk
WiI8AxzNwwMUm9jRT6rna33c4Dgv4I2o0Hh8jm/JbGG34IuzSk1I5hCc+dQlxjeJiyFaf2FxExaP
OWY5aBeKXVIHENqdAPsEx9IYF2nxSwKuT0a96zG96x/QYfOJvdlEu59Zm7wbleGj9Uxp99QKkatj
dYcWqqo2Cp1FnbH/obpzzXKMdQxQEu+NusWoED0d52G8Ru+HULGGcjRdeDh3us6HI19Rmh8h48C1
PMsrAPpkFRtWuWXCv+7g1fScSIwO/suyNnM0muadBXgh9kMC1DVKhmnXUgV/XgtyPD/wSIocsSWk
b13zCpHfaPWMob0nv6kB1Goz9pEWb5UdQ/gjZ/OcuExBcHUhXlEEnxVxqxr7SUbweP+KyARBXdGH
VyH1+fSPoLUiFlUXlx3mAq4ml7fV9A7NyyFa/0NTfYDKin8/frGAI8hb3Q5JJrRs/R2Xwv5o+3Ke
8QfHLUw9CC9P74VzHMbrGUIKoK47JSIR9nBzr7zXjZekbYWtXnjCQkEz6oYYXXkY9RVyMXfS/UE7
kHN/CfHcR3fHbSCj8ihHm8UbhgyDZuQc7tfh8AAcEvWEF73K+HI7GVS28OtPDVJSrzWHpkOU8eWx
66CMZf5D3ODhvwAdO+2Xqp/AzSDC/BUbAzhHsEwBCQeCagSupFTwiccEmbslMW2pp8LZ5pI6Vw64
ukNh/enAuMVGpLPvtwSfLAHORk3v8TYsdcoklAHyYER4jqozMbb5DnsVIAUSTqZDhQgJd4lUgtDt
DgUQONU5gv6Z7YZw3JVd3anZIgplXETe662cnU/vx1oxtdk0aWn5aLgIciMLfVOgGvgse+bdmWyp
bmJVctE2NUVi1LBt18JChBHqOE/SARBVr2KrY28S9lUEqQTvySNl0QhkbK33TSVw00mieWRTLVqy
HHhJFV/c8NT8CD+n9nEN5Zp7j8Sa2U0L3DprV4x9REMN26ypJgk1s7eva9a2gXrpfSorCEZA5mdJ
0n6xVyvtkbQZRL8VeZhvn2jaN5nZo2fgghk/WCh2zBP3jcwEdACjqId2sDzNesHijFvjcGlpCF75
xHMnBznLMuTReNJ+yx/+3Z/WPol01p2ynvk1oHbiFmySOPgctedninSTiwlSrMhxrfwEvKiqRH0g
Qb6Til026fl1PdMfTXzVEGGEkJgTmd9kWuTU64GjcJvN2RqmnIr809Vpvb7dgS0m1K8R6qUSxg4U
Yqz2i0kXfY8r6axfskbvUld+F/l+KWNqEb7Cuy0yMEoi4E1kfitG7/eeQEirRXiK0B36ytSdeGR9
kDaX6Z0SZ41kwGFmrmt28pDTF167QBafH9fzO0Voyhf5fyHmCdj21mLQhWiS3tvtpW/MnQCCGhES
U3SzB/cHm0ydH1nxj/aPaTy+DZEGxuwUl5BGV9gdmRaHnsiRXXkYrKM7WIXKpmwHktMPcpzMJ5gM
wcgv6myVJVTDQsPZo+WD46vIV/5t/dRWhm8F1wEg4DnIw+Tv7lxYJn7OmKT7QbHWpo/SFQCHs+Wm
QIWyWCGHEt5DfyUdpbvAOtMM6QEhYevJS5DFjHy5LcxIPScdnHAvq1WsAYarw5DbvCRqBxHF4+Ja
gK8icRr1v0qLY8VjJUWXWF4fow32b2mkixWcIbYZDh6612Hbf2thMpgWZmmP7h38rFMo05QA32ln
Xu+ac0rL5UTogCBBPn66mHxhvNFCSbPLp0ZZiLKK3Yk3Gb2syNWm/Ley5zqGqDb7YcTmtceG6L/6
nhYHSIObccS0KFLCM8+bllZNtRyzgaxWYt+ws2cPkSmHDws7XvnVH59A7KJU7uB9dEPcftGq0gYX
Ypg90XLD3ItKZQgpAbRzmg523MOVzbG/fW9MXbXpZgB43JqvE8t+41GvS9iqP/mEtPxMnpRZqW/Q
Ndw3Awg8jZ58SwAwlA5oS+yMsqJ0UBOPzBJ8bXv1qO5CRJxVxR4a1CzGsDaOfvIVKdYR/bGxV0PR
6vHzu82IAEDS1mwRoyhgpUYgNJQwUyM9BPSTTCJGTm7qpa3id6upSqU+dv8iQ/Ka+MrAntsSg56f
+03WToriq/1jyF8UrnRM8rKhUNm+cHSKhfv7GLsxDeex7fCet3Klh3IbFdu7tAtSKB1EPefx9yKe
lwj+s+St+K29RvAIhcejWVNqYDxB/EQoHV//fqPCGpoOBqk6BWyb1bmXlikVvqETPho237nUflVS
UzuoyKxtujIv90mMIcNmcImhVGWBMB2h/T40W48YehivCGqQb0OvPNzsJddh5ujiPEEQtU3+i2yi
B+py+7EXqCbrodVFy2mml58dJmDVrZgbfaAkoapZjTLMJCvwu2iztQ9QqUiy91lSOAwSKDEhLn4F
bhf1h1Xh/+ti4X7PgI3MeNslcfOxXUueqWorKqAly9KmHSCHyHkDQ6Mm490ZG9MVy1RX/bPiHwLK
qciWtA6hZIE9WlGi0UEfdtaB1xDCrOZ0vroiCr1+xGTzIV3t6zSA60HJXkU1g9WD9s0W57sQGDOO
tmNsTCSwZ3SQ96cfLMmqscItONOGOi65GX4TGl7s8/w16G/kSGnuRFeJ99Mkoxb41FPVjE0hBsss
44yPUYLaTxfcQKhis8txEfGo5dBEtza5OSkedVYicZ32C99s7nrdwvXzYhjM6OV1UZfz7hcSgNtP
FdHtyHCpkZCqvwtnyEOOwARkCh9qg1Cej4imatYlp3gKRGHx6grWNYseqdHK76o5bJ5i8OSaflSM
ulHMv+jglHyikNuJ7wORvFXoGXVJKoWDJwH1QGTrtw4yzKCZtdPp/KcY1WcTbEU7tLZXKYR/C1os
dNHYCUSAsY2x7Xz9vA5JZLI/LQNuY1s1ECUq8tPhMcBaZi1RUffO6wnt35vwh/R7n097208An8Ir
K9D3C8d+mC8eSwTDCBU9mMDkgPJ7Wo8+l+k5/iI7p0epnoqgG39izIke2+8X/e84ftcDES0qWDq5
7S/jD0TXHq2hBIxrdm8NXkxteYaL3ZmivDzk4FLLCySiTJda4697QbYRqU0OYznHWnJ7HkV6nyVM
T++FtL2E3aUt17kiKVkWhgXdzCTHOlhfINRkGynk/4xNOlU46blpwLCGFBXL2bbxnL66GQX2gTmK
1YJ5n1XhUmNoq20KOXaHq/qsieODVxSu4cD7UFfNR0iQcOsJJQohT3cjyj1JqOrmF+E6uBEvaBb7
58wrqKDo5WQxr0/zPLGz2dg6tL71zEHk3CLMTL69PfKzgamMEcspNYmAqU/LpH3W0B9po6+upTLx
pnqFY2rH/PxBX4UWdl2wEtZyfiEH/VyBG0uhEW70uwj+uErdKJr6WJ4caNHQARvzGlQXflSLH9kQ
DLJM5GOsiXx+rnrQW8pUgf10OVtVyMNnP6scWAEcl51m5IkqpQz82i6wfpUfAccJ4h99HA7f8g/4
Ojp2hU08E0rw2K62OCUzHIw3RmfmpVdm5xjpy04uDuT/xqvezZy2fAFlaTFoNgxDF03cHyE3eVi5
1/i/mYP16AUB3Xuswwee5ldxqBmHtZHBjYzCq9eZQSBFqiCG2HAbxZKRrHiq63mXLRxUig7bB5Bs
2hg7KoyLVLW0/N7sq2YnRIIW1A6I3YQ9PxnVt6b4CWMeXVqIXQU0z1bMNeJbppm0JXOeJMpmT7y5
gVmtKowsrhgCQWy5KvwY6WCb8wkMSTpwyNpFrtT5jvrtUXSq2AuuPxUsqOxBmhowvByzOzdkR5gg
FLb+E7AoXOYlFz6aUDPMNVzyFZWFyCsG+5/0gojCixLGD94OLt11zCc5fJD/8ILQEABNgooVgXHN
Qo/RDqrzqSkorCWmEbK6+XzA/zjYSZRityYn32pSGZ0cDlvAEPScehgD5Y9nPaTav11Ee/cvlKew
Fu20pL24Pc1L5JsVRecIInzUjuYtGdLB/S2sjMH9qRiHrDz7dtEJhOK314hQBRnngZogBBYyyYP+
bEbFlxaZGzk2EIG63G7pKS4lI8sN3Fs2jYGD59i3PG2U0pIFOR7Ob3knb/g1RhRsFfcZcoK+BBw0
6iMysVGgsDmhmnKQaUDzj4e/wMLlGzpoqLMJnlWNZ3meoAAMOrebvUNK/76pdx+s5wN73WVPUnxm
tzqfxQqzWKJh/Lq7UfUiWegjl6xsN6V34V/DwK2G+9yDsWtWlRX8Lj9Q/aujPE8EvcVHBq93Oxbh
0xNh8N9BcLdO80UnhHFX4S12WojfcvAvRnlXAjahIUN7H7Wz93Kihe2Mbr4Ija9fwQnV7Tma8SiZ
sQE8BvrCtQ/DdT0oMJ7h7+75xVs/LLKiCOyV1iopSVeCR9YOjoikbjaagcmGQEGbGeqBVG/37QAa
Ugr5Hj3LxT52tjnYgTusiHVnJ/5sngryGwL0Rid1CR+H4VcVMMSprdcYYT8m/0Y+phhHX35KltA2
+8HqiFbWNlPtqxRl8MXN8SplmUZqpy64Qcs+g1d9oS5taaD+rM/q7uWUPRE/g9V/y98Qz7r8Y7fb
qFApxMUJiq8J7FypMfq3Loa/D9eDVdPhQQxtKBNwWJwG1aLuap/NnPbSZNZ2G0F6kWnB4j7tA1mV
N+ncX2pur26h0PpPVo92zDXny7CZ2RXfEFOzIfrcWcFag/E9UPFUshDBvgX55Tk+heAgOcHSsQhy
hInHijURRW5TYcNtaQ3hmvgzHbpkmQwMescm7u9LWKQkeSXVbVFrP5ubCq/2DgjhEIG/NWeepw8+
SI4RQPZB4EgrqZrMiTtOBCgKOXNHddQa6XonE5J2rxv92ZQ27un9+djD1dSbP2OBex5Hoql/1lCm
K3vRVH3+PZZqx8NaHV6TXtaMXb6Gdo8OZKvzG50bjukoL6Ds1GSQEXG0GxHiftMwsuSAGpqvQH0X
EUTnhZ+ZOfj+c1F3gK2+tpPY7basxXssymCWdCezviTmdZ9xNH5LLB9ZbeLaAe5eat0wCeTK6jgr
l3xtsH2GaTqfAI+xiSecrw65i8bGj/mr7LCgP0ExEteQdDTF7K14A2n1tzVU4/ZkcFl9Xbz0Tlvw
gAAna0sF86+dhK/HzZuyFwzFJDnqLjeNuFmZV3lE+KAWTwT8kJh2HrIkqKrse2u+LYOqCjhg10+E
kMguF4pU+x5mzxFbUmGUfK9X194oGyPEyT7kxFq8RAQNfwq7+H0kI7cRUrqV6fmsCajwrpcGxWDn
AsKZrkjeS4JWbWuOe/HSz0/nyk10rWCXhpCEZIlx4ugmytuBEmDEfsgQlc3PbL/JvHpt71wf3v1B
IXJix/qE0IawlLCHkdtUm14+wadxFy0MuFypmdj1aXqE81SRmyoyxkCW27CIzfyymafdiKxCBCOG
IMpz4fGE37v6C91yVauzFz6KIE353XK9I1OpLWeMTB7AeRVmoQc5X6TVrCXjKokWW970Lw6XN8+f
26fkkfrZi7Aopo48uy29bc4BtJkRp/BCUgUou8SNNpaAbVMiqBBsWFwO81bUDjX24QAbwGgcjgzy
byhh9ydhm/+A7SM3Hgnvsm7PI//coTISJ1BzP6KUpIKlD+Tbv86WhoGkYbKa/seUEDCBILxulP6n
nkltyDuiKE0pU5Ps0LHvWLEN6R18Znzad+7OtV88rVArPapS9QKKwGC4U9Jruy7YeOAEmeyrOUs4
IxHXW8WlSJZ3gmnMhr8+H34YS7isTKxFA2RrDNAfgI7oQPDrALjcstru4PQUxXf/+pmXDlhQ4Eyc
o1APJu/Yt4RnExw3PR+LMbsSfiEZkIlX+czT+/7DaS5+lVbkFU8OtXYFbFlHOD0s9JCSo3VM9X8D
azafzaEKlTzod+XYK+7e4tTQtWEWBf+qcVp5TPAA+1P9IbXaQD3iVGiYLX0dD8+NE6HgzTadfU2O
qN5arwmAkWBWrnAQVqZBtLQJk1OIlf6c+1CAGdB2aPykGssgg8Yhcjds9DhaFMFsu+LbDZLflO7P
U1jEtMJopcgAxKTbK/ttqW4raVLLHsNrvZXDVUCBNA1P+BOF1+nmtBAGvjPbxsuIBukm/FBGLQ0q
ZP+ucQInEzUSiA8Bc6VDtikQTm5SlRo696ZdKu/QRY49Qz34GhYKoM48aZIYx8mrS8XqKNv65sKS
l1K3JXdJMWev4DAA3vTIzzZy93XQdVrXFdEDb8IKo2g/eTaJfX2B5F4HIrGmwc9x2trVneEQkPv0
jXu2NkmAIYYlisbLyAuaYJJqBzS2ftQEg26fN+MVAD1lbuGPfMWXHr6pa1nIWrEIWSpV/qj2Abjt
ycjud7ii1EYxlHmxW8s6G77sjw8ENq9lpI7zvLdyi/bCLHXqrw5SCY1e4gdsy6WbI+GES92a5bEz
1zkSbf+NmG5jr9eTkgo3Y6Fm0j4M1oJYXu+bp9dlJ7nYZqTKuyXLA4Tg8TM45f1Pk5xPnkKlSdi6
TreCIl/VxHg/S+sPj+vaOoJi1TsbnAfQHpt44Obb2+D4F/PnRPURfOHs+cCHMK95FO01wu0YeEhb
eAyLGo6wj68hPa1/gvCsoKtNhm4+vZsnNmC2/ePLNoQTEDjZf2RXCbGwP07pVbkTDGNvOuyZ6AZq
ceY41rRgE6ydlCczT2ogzmSjMJU4TmDvon4U+p4bt999Nle+OzuJzIMIrepv3zBM0bd/juA91laZ
V+g668vSK8BvYsRnjtyOmA+DQRleTjPEKelSwq6OItj0ptANuSt0ydC/Szyusz/g7FgAkqY82RgS
IiOjCf+mrmPltVsjFtUhpf9dyjwekfthX5GQnLxEwlGiGI/IapBKCi0SyA/SGdYxCsqvO9lvhjML
ba0szvKr+SFO85RUE6NW5/cuJoMbDxSqCZIiw61ktnXIn44jTNUpmmvGxu6cuoyVICzB/ewucnQX
jkH3GKz0g3hHq3qLmEMCDCpqWhshmfJwJB0iTf/mq7xJhe06Tke3POn+S7U/vkT8q7yavAj3o7Hf
/DHrYgP6+5aX/7hcRHopcO7YSIJMIszpr2Eq75m9GkCZ5ErZjZVYdNRP0ExyRl20b1B9WOPd1BF3
2ReLLfDaIucrUvKFWi41NOS6Ulh4y9eqimL7PWRpycjsOIOhWy4hIrTRoYs+HpPm6ex71Pw9drN8
MxFf3WI5No2aPAieYku7ZfXAOxKUWRhIxPC4R5q1O5w3HW8TwdolfecrBR7ylGiG7SgoEaztsVlC
kkuwfehXEMhrpbEBu3G//aasE0Au0P5zib4J7WAw77Kd94XIbF1Qpp8DU36vBjLRnj9CT0mzjLul
X23iOQtMRTiE9tZIcq97HjzvYteXjPSXvbtbvIc6qICMj3NZ626CjQhBIAqFMwGaQtWQq2xpZt9n
PzEX1i34YKQ85NgNEVaoD2mYTEEyyanJgBZR4BYegot6+nJAedGkRhFtpMO1CA2TzgzSE1QdixKl
8MIFt0xbdLm0yK2XZyjm6VyRmoGoc3TXLecfK2Pw1ate/0CIzsWfC11tEJSFbGWybSSi2Ku6ejUU
VpkND1AZzbxGJoDjHOm494h3eeyQGVfrhPvFD0YAN5CGED140CCqvyHzWG2sKcizZRbOGjgp3rFh
1duTpC+MKnlRPCEHd0jAqm69ADDiPRtBc+99D9Q60XvJD6SoJDHE0fLlyy/vaekaNIJ7xlY8WYJu
nc1bNRef4LfXQoRiafdLQTE+7KDvI4Y3cT7nhB1qhmayqxObi6QcNke/b4b60WI9r/SFHzt3bsjT
it8BDYFwQ/afWxUvRICBKGwrIJXIe0ZdYFa1NQP6NQk0B8RJHmezvYfPAb/HQgPmGVBOV8v3sLWW
3RV/U2p3/BpQfCPNHu/NVWmB8dU0JxljMUdCSmqopu6YYQC7h8vETN+TacwASsxJ9tZXgPxxpZDQ
jo86xZCq/BxjqyOtwEvgDqsvz6X74CH27MRI5TJq/uYjFKDaQNxTE2ul4i/eTT3mmEFh1OmregUJ
89bgwED3P6gZZEK6ZNOr+fj+EjWQw4FZ4Jm64YKBCbvn2j6S0866Af5zDM+pJKO4Bv59OjwIfk7Z
dIn4pVxW3qKO4WvLN14RRcHYeO8l4gTmQhmSiMvdR+l9m6mmccZpT6UT0IEbX5v/IdJWZvtcWDt0
qqt8LjzgU3dwBkKiP/7ubZ2MXWJgoWQb8cHgNPanRTJreW/j4rsE7Ol+W1BGn7FBQNhltM/x6DcB
CfcYW1jW9ZXiOYug0PFaEiUA0xDmvZNEuLFD6g4bqsIo3woy+d5IEmEOzj2GF0e2Q10d3BqfvDgK
Y6DDBLZ/nnXS3JJfhSoT3XjS0yA8GDebuevB3VFDPhmET2lK8DgxxxJKVftC19SqO9k6il71zWeQ
t734IqR2qakD/GHwpWmx/tkUzWWoG1dhJl9qFQ0wwHMRI+YF3z11Bx6yO0DFJsaijhLVXsH2wlgx
VOTczA0Cx5zAC4zUJZLMYxI5s0slvelnJrw8kGRbDMSPzzZZiPeOVxFLD7mMlW6dRT2wLJa9oKRw
gg9pIITevPFuWpeEGa8gADwanomIx6DwWj34g7DcrBmFipC6ik/dhQjO6PbHllcCskDJ5x58DqIY
Ium6svTR5wRBJfWFkcpvtIanH9tZpFJC6c8eT3C8/qbPWB2GNTvXowOPyD2r86S6H4ZRGhuGZc+O
6Zw+PBF3iMl6RdwOGSaza2W6APUmnsg63YTDX0uATQw8rBDSyp53ikIg2VwAnWu/N13WQz+DsBea
2EC0tlj6u8ZMpxqgcKIbhAZDx8BBonzpVtsm6SN44lnCwn5MwvujQ9nqGsVNrXxna8TOYqkoivQK
L4o4eg9u6Lty2P94UwLfmh1HxepNghImOLYaZ08zQu/gEk7XL7oOMsKmcyLnPW7qldyG0pykY5h9
m76uGRCgpAeYBPHVbW8vpUCOtoCFhlEvl987KJ0I9iQehiZuFE2YEvDA6ytLW5xwM8ovOudw7WmJ
U1hDBrCqwNTYpUdvH1kAPIBNqodVNmCEwDMF8RUrhRFJ4treNldaYVjuHkvufkxrji2CpH5i1kds
IUPGpgkawAUczT/yOYxMU7Jzq39c3OD+yod6lWck5Nd7QszVRmXhEhwOL7EdMDqlwakFmnqQ22gB
vYkRABRoxQhLCqhmxnEALJ9tS3u+vhr24i76AHWUQnyA87j6a6bwhMQo4crRQhFm31Xq7D4C82W/
QLfJ7PU8abjW+g5wRMlVUZ7rnJq0sAddTAB8dJ8QHROIr379HpnHGKmdvPP66bNjMT0iuJU1DmUW
q/3DG803i/b3W37eJ/HoOPh9+VSq/xTwUw64QG+pk4w77Ig8GTW1geqK3WvFck8gvOc8tR9F5nWG
TjIt5eZZfZ5BClg63eXhFEDRKq9oj0D0q7SkE6WerPr4IKTeXkYOoy/sVk0Ul8JbN+JO1OIk161t
Fy8JMh2i8Q3yI14imESPL+Yxr1yWkAI+FwiZJjqpaeALnDFqsesXapLHjKLT0AakDlhc8VQohprF
T/x8l8fmktulwm78cIoWVDVpQirdeEQ61emF6jE9AfsLn4cTa7BKawe5PrrPPE3H1zUofz12hsjT
RiMW3pKAm75qK3jxc8EtFCAIyjcTK6lqVDBpE/cC6yX+6U+MXvl+KJnlOXc+Y3+giXRjJjZwajYh
Q4+Ip39YmYPhwM6WKIkCmDntDCYVqQ+7yY8g1Fb5jwzcjdqcKiOld5j849MtGMNrmLcS0bDUluSL
+JQnT4a8rxr4k5m048zPMeSfbf/dOz72+TVxxmDSGHBl+HB4b220qfvT+9kUKg0UBqkKdk9oT5cm
EVNHAGv6Yzca7/1GoXfHj71HGTGXQwYIHiQumGkGeuDdVE5CkDvWAAZMgUTNxhs5evDhCdLACx0u
OiDIqq3Cmoet0M2oCw2+5JxWcxYOnsh9sO7ItamFCTZhYHuGf++mz67brSywXSzAaAAMeNA5FmZ/
0b5x98tvXIz3Y2AQyMwb6CYSGZOpkqWMxFBUlcD9N54Nc51q2iqrcuVIrfjdUCz2+eeoWOiZfn3Y
RsQWJu8m8N+duVTIEvJmhtXZAJAxcAHFJLLsKMbXOBqu0QGIqNqza1ZXSQXet6phMihW/xe0S3Cg
6Xw22ggIcD7r1kTdNVHBq1UHMUm13T5vhiC0DJbRGAPYk9nZJiGL85vbMscMi9EL6/NCCbzl4/WD
HC/kQFKj0WWL1XABW19/cg3PwOXj6QLoZXLlqRk3daQcq+6M4fbNR3advtbgAQx5xIpyb6JyJfDY
+rnbBFJx92qT7zf3GZ6TKoFZC2og885wIHsG7Zej99ZRZaEKqiyInJaTr25GEYmYAFZ1lwUPtna9
FYogSTo5psG3MKd0ltTptA4g6j85A1pvmBnsvZ3OJ4FRd6yiofhm1mZFrz1rTmUFQgTMKspnr4u4
8MCiUgRHvprLCN9u/Qhiz2XeuQdCTdnARPmOMwYULiPcKpGTeGKYUPQ2p5W50iTihLO5CUQg1lBy
D9RGpzWnfVN8m5vlJm4+L0igI3G7F2q+S6esYHsYVqv9U+G/9qR4pRL2TB7IAEW2x6S67jZPo4k5
LprWEoYBa8fRY4VNW2z87bvtjcKoRmztn2htxm9gp7H4WViuk8jeFtoGQXi9O2rRDXYsRQ5cCybP
n0FoqXn0S8z/XgtQEoAJB6xlIqTyCVDH1353qPog1v/eop6PQ2BbKoR9T7srsAlnSrbqIYzu/Kol
3gRu/QtPnhmJVPCHVJqVVXcoU9+6MbOQyWtfSVF2VNgHE7PVw6MPGACFul5IQqbVtJQ1Pq4CfLrZ
1nQXWQe1aEC13sE4wc63/AYJ3rNAtSkdZ6f/i9MSxZ3R+VI9uvz1ILG2QmoQaEM+f+XFaGRBpYiE
3yByxvS5MEi+4g2kgx2yp7RsXyHp5+D8RGqnAXH0gWOC1RU3ZCK63WfzPFZPR52hH15raXUIWVMj
Oihtrvo+RQq7XD13NXJGeaJIa2Rg6n3e9bT87QcQF0oiaU5ldekCAs+DASgkUbzHMWtzJ5Z0H58I
ZRBl7N4Wal0kdRkCAWcxw4M6X2cGDV/Qm17zI0nPRNxoAtrEKiGfh8KSx/cXQKMMoLO7LKia5LHs
7m/4Lh3MxW2VtWvEiNL5LK3gt7Cqwun9PbRCzLz8ETh45X3nYyIDHsyFhHfJ0jSdLO0G7NRcHFm4
dGNV/oxnvlCxZx86DyXNXCUrlRsZw8FEcXT5j5bQvq+5c19UIEqkJtyZ6iRbrADHYiqrkCUNTN/g
h2SRwzZr/a6SGl75VJSo7qxgtbQUZdO7Q1uf9b5LsTnb0T4k5CKUh4z0jQoUp30kX6M6gh0qbPo0
pAapYZkcCeetv2E68F0WX+DuwZ0k6nfhaqpp1Wb2BAgI8PaWRJ1WCJJ7iZeXHAD7KhrNG8RLtWsG
hZlVECIT8DII5AEaDpifgY0NT1nX1/RFJQ2BpZwI7R55xoQoom8UiQJFFdTBAsluuwL8DuYkHcG+
Y04JRQuuMcGIVTzOFm+4QBYvgzUrj+HpE46QodWGr8sRzU2bd9nRRVFGxiIiWyiLTwv466BvVTwv
cTJJBaI4haxDkB29ddeecipDy9Y5ErnpaUzAiSX1FATfzvmJkS4uG23ZFWmpaicaXl7CS8R48UIi
jH1BM3jQ8jl+I9st61JpjhZhbDea0lGb2wc4ESW0glPaCueHuH+mSeJeN0tqcdxmxpRFU1oA+jbJ
GDRDy4yohOHep7LH/Ss/tNPTVE4AXCAaOCT8EcxvMlChnkX2VTRvGgI0ksGCRUeWCdHPuzvQic7G
K7C8pDPlkB3i2zTguYo3SVxDDxivT6uUQy3BRjMOSJMHXFWJ3neJAXHEHeYPBviIyB61znEb8kdh
I7x8WaAbNgpGuGtenqLOADmKlHUEhSK/GQYpg/skvl0yqHZiTzSYB90T9DMuV4fij6slnmixLVlr
dFeG/xh/LvLJOKlr0U3Ag7TYU6Srg2CaEsINRBhOuGbIpow90S3NUkLylESaNElvYra1yeReZHC5
6c6/k7/FoSJSplu8OtQTTrZG2SWyqT2qK0smkHs8JS9iBeFUvg73cx++0rWMDjpa/b2eHlj/BTLz
dGzBZk9sfOwXsW2NQRCZMhEj7k/BucMhyMH5KgakuJDjIbXaddJYKmIroWGAUVwbCkZUkoa9i47b
EVBTOZ5QQwApKbAq4ozK9/AHOVZdUs1GbbuWmtclNtvGmFCMEiMzil3ibjSV4DI64NwZGwdH7kly
YK8Hkh0oS0k84qmE+PeWEaU897z1FN/OXCr69Jljgw4atWga7eL3vb3F+kvmMX085LKZXBzZplM4
XN2sHi3zDrsV8e0fLegZUUmRav0V7uy5eyNK124C2D/ERgLtrjor1gxb/Be89yiFL1uTPoC6fdt4
7gftngoLiwJa43DmckSmd1rJlcVEJ6nMkGVH00Domv9rp68A1laFjEFboNMstIEg30tufd+05KrN
6mG+XIEbPw4C2nw2lsLtk+9Fkk2KnCDY/LRn2RR5NDNR4ywBFYmotK7muNbTet9SxPiaq9PGqD9m
tt0n/YkbFB/si4S3Bm/IEbHGWBrLSH/e8kKy2/9eGoGVBV1cwX70fw1dLI5Kqs5Ae+V0uOByVrcl
IPO196cZflXFXYOoHqyKoO9wn9QD9a9FHBu2+wztgcx68KI8iBgK07HV2xEwKKdxxS1x46PhkZyn
dKJ2tKpQdi4g0fahDg41WqYuCTK9IhZj79Ku1mtVnASs05t7v4Rs8bDUC+KVu327x89T9JTe0oCy
ygxBwkf5Yf3WZy6R1FPs6rLopazJAApEzxdFLNAojyfWrg+kTfQ2EhXxcV3I1+j/3o/Aynmw4q5n
gjr4cstK0l8bzUmRd+znMH1bdoziLWaGa10qmk+gulFqyj6Eb3Pfzi+IBIkImlKt+EvStDUhHAvc
0VJRhG2+JEYOK66H61QX+KEd/26KO8pZ9yt6khxWBT6WssWEUm2jos/SAI/ugEKYdsUrgpjKmpJo
/GYvmXzPW5jzDqYTJu+iuxhxG8zxKEPf0WXEtKMcLSF2RbMuYVYm8kbamsb6nFFYiRaV5IcZuYy8
osTF6WMnbVxqmb6hEHu7pwnfoNrzwL5m/sbGF7/3Ju01ihu92oDKrGh4TfPx7XnBR9oiFzknzz3d
WhVD/JgFy0KVe5vGzjpz4FFseuTnP3XMjQdpThNscE8Ccdb8+nZdHSo7MmGGclGkqscMF5w9VKhg
mSyO1emFvw13n3/FSxe5eYZIDjmZoBoSVyuGN4WUtVIOOVtfaH4WrMdmw5peCKG5s0VlKxx/OtUu
nz5rYsaJ40420Jfmp58x4FEbwURdyn3v6PqCKY3sh4o+E+2YJzpCinpDHX5jzK5MOroYwydX6VY7
eGp+Xm/ddocv7nkpGtbOD2PZZzoZlYgDScCWMKgvthRJ7kK3qDuXzoxpwUdLeo1S2ejDNOKaWXLh
2kWuhatwZYakc183O1IAPVPNBS2GBhZoNb8f28pnCN//Z5lt898xDEAO5fw4EyimaX/YI43sRDgG
4jeChEciaU45FkaylaOLtUnBSXDe47t/4WjW3s/2mp/JQU5Ifq+2TYdrqaEUrdUTHsopccH4tDbc
I67nx6eAB8M4ghPI8I/qJppPqER7dKE9WVEiKD/E79OPuj8ysGMeLbnDZ9Dhfa1F1Q0wqizv2nnr
xho2RUDIt6ycq8B4hjB/fTZcW9Tc85XJnsV4oJrdZrqtaCgBVMV7vrap216/ByWnHMd8oLGwosHX
TVSPJVjnVUuHDR95V3BpwKmTI3cE/ecq8QYcVgY4+29ZAC4AVlogul5XKYIGk9KAHcK4bZPQdjJG
EhDBw1nXRSXlDjGNMj4IGNk4jxeMYNkcDKGGmDEjCKrrh+rhdQLZDO60BfKO2ipuxRvXyuQJnGMb
Ihgee+ZCQIWD3uCBenW7YsNKi5OVSn6yRzOqN18drxPs1pbHi1mocb+NGemRG4bQ5z1RSenlsPFj
mT9nfu5iUMcV79wcZmXPqU2j9wCofUC/OuJtWSta3myXhGITc8FftB8y3/tjCduKbbAi4yu30sPx
ukf0OkdEyMk78GajXu4p654Y12fnrtfUGzxJAqZFAw5U4GnvZPtFO91L6m/6yn2sjlN2oCkH7xfi
4HqlytKhsO5GJfEzb1xUigGFUa5A3/F+TWnjCEueoE4cJBaK8+WMb7mRZ3FKXa/btpLx8QmUf0tW
ypcya5pIpWW6ffpBMIF3jCcn+zQdd9Eq4E6qMuxPkZXTBfsPQZQqyyLxEPV0tzATSQ0KaGz0Jzkq
SGYGeraUSee9elCTqiOuue1H5wJ7yxeTdIRKChz+0cVHlIGbomBI3cdqEXukFm3xew/UTY/6U68v
ATogUovgH2aMeUPAWQdKmDtFIdOODfa9iqp/aFDrmdNl/38CxyGmOBRifMVxiU+ZZLu3XGsKR6Bm
Tbk6nXdS5gxv0g5+j/aCtb4z7pKa9Op5cqYjIuJg/EMg+5q+D+Z1U32bXG4Uw/n5yd0qfDqRgoTY
NEfggKQLUHcmVIvEbYiDD8Jp5hYCVQmdmbbNuXIm9h1WzRoaGnxJEr6XDHc2kJZgX5Jp7Qdr7IbV
teRvjdtBDmamDpCVosQJIGeyzSRvdaNvyWdXoMtk3rW4XH3vul58FSBOhWek5LMtJATCVK2Ola9+
ABF2y3Puo+07/40TCztDWN/YASPxG/lQD7K1dNrR9mLzNCLgI6xyMf4rnjDzKCYAkKQsaKp5SWu8
G2v02lcHxOV0OMhTjD97QGNgvE0m9lwDObvWpekF40L7mhVSVhZtiDdFv2S2eZjPNV8N+XKlcsUJ
MLxN8akFh6WMGqydQcpOQbS1htXNWZ9lPrXussc8bulJ9n0mgndoSEV5/V3eD4WZSlP0GDMP5mvH
HxByeVzo0aTAQGOrxzZWorrmSFFOXjwzJ8jzIwhj8r6K+pyOXfyE6Q5dCDitMdhEBBbRE4nyES5E
9nWZniGJXXrd1A+j9kxHGBVvIBThsLJJ3oGwZHUQdORjsns+qkgzKv5rNo8kpmtCoAyFKqqEXo6M
Sf0cgFS2K4BicGZb+edomOueR9G2OTSmhqk9mMZjoI5OJ3k6b/D1liUX7FikGCToQOOYrXGoaAZ8
7R4mofSkPPoDmwOeSuw26sQhhQdDGc/qIGmknhBhvW6NXKH9I0TqpnAkgQlZS6GNyyXC8LyRp7hl
NyqlEwP+APnyfxOGxCJScy5haY6aBv0LaQD/lelXwvgg4UfGP6KqJ4akHWnbGO0Q1rwmT2doxaXY
CGptdQ6wuFh+k9M+6OjGTfnDyOWR4jKKa5d6Gj1tOOfj3Vyv1fo0zoxp4wKdkscQvvhULzUhYWYD
kk9qBd9G4uiRXSstBGdwQPSJShTWZcHSv0pQo4OhVMoxxX674T6icrrEivPBIo+nORJJLrvNBAbr
FgN78uiwZSlCn+1VlAw6CcGWygxCNezbo/yeZFJxyfIf2tiNyAqj7khdKuc2TrAehcblVOLCpytX
YLcQ3mogaY0Pc4tNDmUtsK/u5mcbBxd1mVvu5Esz2ZovCoduBHYc+kFPzduh3DU5+UpPGW1aEVC+
gaXXGsTVZT6L1d5TB2fnpId5hf30gBQvSGkObMNFKXr0xWDnkJsV/vPMwktWbsr1DtEIs1SuuHZ3
fouwy0+uxW8l6PUPVY1rVc7qoAhEcgc9Y+u2wWWi8iBOwvML13klDsbBUt/rPtBdSGWqtMrJeBN1
nB7awoBmwknSfTkOHNUnck7wXtLM2XmqV968QzjxpqeDQqjGUTjIPkBf5Nk5QEZyTHLatKF6qSkH
d00vIbalt2z5jMldOKaSMvdxayqf6DQ9TX9cJD54fQh0VZ2uxDuikUqdRVInovOjrAuvMvtq2wk2
0BEQmvNJ/a0tSlIKADSyIZlzunwC2g8ZHqS8yC65D2VZNskZ8NQRPR/9EEi1OgelwHu7mOlg+rrc
gfnSwexhmrT8AziasgqG6pl1hh3icfYT2/PAIeupOimz4yVFH5i9o90AqLfWQKMdNGspdoN5x5eV
39ZotDz5ZpqmwALSJT3umsdkCvgJ8pLx9dzQmWrqwzjWxh+0apgU5h6FWiZkBpyj0VnwMEMeK1zs
mwgdGLo3moVOC+FAbOp0tauQVdV8SDjY40slTdvjktK9v7ohgcBGCdgKYy5R+0v61pv9P9eNNglY
Gui1dkQB6D7zvzTIQsYGf15Ffni3bsfeb+5b6aeklwEVnh2EyOeHXytFI6UrSrD+CPiIOUKdBkiP
+uS6VN9C/7EPTdzooERAKW19fF6K0wghxRSY649zgcBuu6oZOr+UVA4qo3RjBR3/QUYqZlb6VbZD
GEJnBaO3FpEtAp8kdLKW5aREBpFSBL1rKPpi44MvEoeq1HvKaOWMI8VuYK95jMf88VZZg1thSIWm
Vlsjf8NA5kQCDkFEExUQi9aWZ/Z4S/gVaGrQWV3y5rUyDAoWIhIiecZ3+L6DKk/3CdEX4DzY9jmc
UN86lk4e15gvpPGmp6IH8dbooOVScdfVIpViPR0nvQ8uGVFspVcfU09UfWx1ci1Aj0UevOKl1jQ4
Kp+3BZLqDtBsTDS6zll07SrLFVro0FbBropzzrdCHlgvEiukLg7pCuWzkKjjMJ0LlAqThL0jIGCU
etWdE0upa2ARSnMfE44UYiU8m0zCvwO5JKtX96FiNTgAB0GPowgYEL5do/twpBa8zkY4v5xhVGl2
24cJ3kFcw7QCfaGXZJZwicRfCJdtXnpDaT9p0La0JBwWD5MRpluSehoY5FhZ2rb0FF3tHnLHxZ9i
YVu5v9KJouDP0tGxuISu8zboyayK9X+uhF4arux6LMtq+RAJrW4ZDycKIHW4IKtMawIkWGcLqv6R
mS90zzYB1/khKInSngs5IusEgZw9bm8AM/7YDanlbIMrV9TOQRzSFjJSei0mbHonLcYR0vYmTGnX
gvOPYRzj8lmfiqIhY2/bXyOUrtUVm9q3mlV0Np/Adfv7q2WL4/EhY/ZpW6hS4NNgoL5Nbhmfc5w2
4wlsLfes/UOqT/WI84zw5vj2aCa2QBnmRcfCHW4cJ7YNqkiw3+V5qzylTJVlehnJAergsv25Z4+N
0bDR/0KSJn/olKKCAQq+blRvWbq22kMr141USslIpyi065ke/IheqL326eUf8d/3tpG6nToC1MFy
CM1AjlCsrdGtWEt/znX92+RVC4LbJsGWb430C1aIvPLE0d0j27px9iNNpKAVaIjTKy9WejU3EJXf
QLHqsRz08GUz+nK43eYNSFiy6b9pjNz/I9Fl2pbci2im7R0mfi8swWWJPcDsfXmIaXjXnjw+jFDY
Da/G0CZ7Gstnh44VKS3O2ovbWqqOnVDMzpglYPNKz4SyV/pF+zpHQ0cBv/URRvsVzVxVzHepXZbf
l7t8KSq8/esgKKXtQyz5qjnFur2TRVxVNQW3wwZlK5+tR2He0nRErhid2FquZd+Zudzwpz0NY/8d
uYQ4CXbuR76umQuzs+XUIn+CJG1SdlkZ3aVLuMeP1xHueF50xjrWKIi5p2yOtVAWvIkcc1ltbExR
YuloBNiWEQqNT8YOUoybwHtqx9p9u0kVEl7uqemQlCDmzCP/B+U8a68O151fLACjEoPaot71vaoS
BAopi+jNovUs7r04YHHjJHf2gukgVBUYQ7OYEn7QmWwj1Gnh6zPbBxgJaoKa877jHq8NH9F4Wpd5
ge2A/Gltph8CMYDGFENDNOZN1HW04SsClzsVbHOv4yLB3PhFiB07fC114e3GcwU8aqHaR/sme8BE
lDaenEqeCaC0dfm4t3YMQObnrkxvOvYeRmWOHUKRhAJ5KhadlB0uvgehnqc4/VP3yOywJGC5dOfr
8pq9+V/N5AUrJGGw+3IMzFbhxBuyP8psPQ/NJv/GxJDUppLpQlhitHIqBx/J3sQuFr/3h0szMKd2
JvjMzGgW+0AEl4dQAKXzB7kmWZpIWCsACagK5oExg4wcZLE0ULC1iBZhA/swNdpvOYjiFVND/PFw
4YCQe4Vh3JlqwRglWqYJn0lUIYhH6HhZUmd/Q7oamxllxji/F2J5wPf8QecBReY3Lcy53K/fhcP5
aG/DZDq5bgoh2FmczlPLaSOF5KMB188fi22cV9u7H1464TBx/YOxbyLHjFKy0Az6SFEcGfHlivQ7
dkiNoFi0wrSxLhPW6spebqaxevMnwvlX7LqN9g5kuCcPphqB8y6jq9lEKa42XYPDv+tmJljvZd/p
HCM9Fm5W+/RuKbZGIpE3n7X+wm4OqOu0GtMlrLE14yxMpc6mBvVeo/lfLaR46RCO09OMQ39edYWM
m1Ahgt9IfvvM8ZTmLWfbxELPSim+GBpZsrQGTGhHUoyE0IxIKlg4x2QX5suj6MCsI27u68ByoSzU
2YLAXVSw2mqMZW6BvmKedVsSICoiEcD1qZCmfMMSYobEJdVpR0y9mTOWVjHVhb/RvYn/MCayXLiQ
KNGfBLn+zIyA6wZJvLzKO+GkXATEf1yfNAXWP2OG0+LM8ArAmO15pOPUEtaOi8wU8ZaADHcMD4u+
W4TX326ayQ4Kban+w8OH1u8lcpBj1zT5qvO3lQba1yL4U4qi9UZE/igdjfrve22+SHBVdNuBqqZj
85KsMSOJwArlBHnX7Eros1/h4WYDOnBYd8NQw/1+Xd39odCtP437DubTZ1K6OZYdEtfr9Gm9AJKs
bFrds/Op1XODzQO/cKc7fk9IW1IQHDnY3lVxOvw2ScEutvSjU+sTcuF4t/ZnstSqB4Zk+y1ZAa4U
mXLMdq4gPMpWLrZKWe723IEHYpmobSdoGckZlIhoYUxVi6XvE6iDfUTxZ4KTxrR4WE8fDJ5bCHtU
hBTIyu2HdijauqpexU1dLEnIDGd5bbSD1tiDJZ/QidMMJygfMbKAJEL24IjfDu94wO0tsXXjhT2X
olfWrqtmrHTxq9trvNd+Tmt9frEBKSN6wBgLdFFks88NwTLI3bz8lWlZdaT1FM4A8TWD7ZewAdVh
eNVNtE/oQht5W8SiiXjahNfZTVWpwvNxZGKlTy9SselOY19Jy90JT5cuYUOv8uhNoxbapxhsTmzM
H1YpROc96DahVKfRmUa4z8nciV9Wu3mLr+FWb1oGpPHfJG60h63ToSEuBYrhyKM0WCBHfZ14x9E7
E7CBS10OFZRzrhlPE34aL+qEMtsKo4d7kiARCXbOd26w098FgH2Z75vznY9hkTbKIvXO9VmiXwoF
xiMyBhGbvQAuUzIO2xNnye06m+xpilKKrJubVmjbwKqRRE6NDonauAujH83M/jRSu3XZfCd/i7VO
+DPZzPe4tFg3YepWdaEPs15d/hEFutYbYZ42ryXWBCS1uhXcpkcbTGIhnbVTLrnK5elZDqa8l+oB
GkC48g4GJykJ/5NJ31QQiJuOr1ocuJE/ZaCUXkmIgs/HHhkNXOHB3lJTbVoAzjv+HbzjxCsUtdXE
zhC9sho7okif/jWcHQFFyaULde2YKqAdm2fFSR/ai58OpkERGjyIw/hREbfxsFa52pI9SSlUc1ek
1uoRHOLLG5JlAyPjLVlKk64IUoL8pnmkyWHI56aI3Im7WtZYKJgAX/o45hyoG/SKRke1eGZEndm4
ZEQdE8NRFn9EHwkdawUNkQGAuaGzgiDFN5eMN4XU6kNC898IdLf0tM6iqOdaqQ3VRtQV0gkcNrzg
HcX729z+VSmj5C4mmU8zSDGxt8QG/2z7SdIad8vKyCu5VMgxemK8zyjvBYoCecRwiwAJpwDdNVqm
zPwJMLiL9kCQmEmbRTCLH5JOf+OfgaIYeMCi/++vbv1Fbq/ZpyN1ef+y/eaiYiqCtEN2gjB3Itv2
2kSiw8iSI3e5EHnb+UxFZN+YBUp9mqp5PIVGW7Np6Q+2Z+lJ7ZxIlSCusDf5pJbIRLlA8BZ02H33
6uA1TM6lgLn/j9CpIIvRVRt2EI/cL4e8q0+Rr9YMB9r5STly5LzOvFWPjQLhwP/+nrpeNEZkefbw
NcUUzPMw6E4Kr8bZsuEX8DCzJ6EgOJSVDRxHc5DC3D7uR/MVDfQQ+iuAtcweoZ21uMJA6qXz2K7h
i96nsrgVxE80OntLehFZSnkC4Hj5s0hZ/OkKPKCjZSm4ydlCB9tE73zywvShZerI5c0lM7YsamiB
lkMqnPOMMhQEs3O2NEfjS4QD48bwxyuByDh8l/zZEZzdye7A+AWPWOyrx3CEwca1gux94DDhKACK
pdD5p2MISNQ7FztJ+4VAhjzfupVcF4NrErlAepa9Ng9kwa0MGajETAq+4Q7TDZZySsYW1khCsHO7
r2R07/duGHDM4M0k3kFufBe71U0FhsgYEPMcrpt1O+4FRcK3754uTFtsiNZ983Nxv9//dX+Sz9X+
PYcLZU21/wFYU4RgoC7tTKB5SitSndYfrHhlJiEm/hPl5/lIp4/L/GOzQ0edS0lRj3dYNrK+n+jc
9eseivkKbbeQQjThUVs2kCVoA5NxInzvKigY7fg+ZBiDSpxr700fqy4ygVzArTRwJGFElONtJTW9
HD8CmqYgm0KfLjBJgR9OGcp7ymPTK53q3N1lqvqze/v3IvdTI0Jnclk5MndqcOM4d/2ny3vDM3bh
oSDmalJ5mc4uX6dLC+nB0R2b6IwiUxro2nDmrj5uy/Sc94HIQL7a5Dt62QQnCF4a5SbHhJwjQLJ8
kwE1aS4SP7yaf8NGIYhfNsP1cZvw6iGisXUn/bZ73TJLCLDThS2tnsW+B5LPk9z49rXeKWgy9JmK
VqzJZfBrVsp5z18gZO3+cS53torj65piSbJaN1qYShBVKtBpWIQ8a3gWc7tGxzp/vFCsjz4e+f/t
0BDu3ldru4dwID9+91241ctr0N04mMZ3Oqm48uspVVI4MzSMGPij/tPsi4RqqI1fcW9G3x9AgSR0
q9M7bG6WLG9CdbIA85NWY3xudiWFF31mjbF+j7GsNIdjec8KDStHSWFXK165PwtUzCGI/Vcmc8wU
QV6hflAVbnGEcVW5lH+1Ef3f1lIKIOON03F5JIYvBG0LKu6sOP6kSCcACHjctkjKWp7YV3VMfb3/
nLtq6xHV9yFlUCD5Bla68QG8letn7LATOXfSrunFZdFHGGA71iC16qczQOdyvJncve6Ijx82H9K+
+I4GFOSKQ1MPNG7j71y8JCNbpEEKdjYvtW3OtAKIdGbBzLTP640eQThCJadJpnAMLh/vl56CU3IM
/Q9zisCnGYM8gbTndaCYoTrY3cxP445YNrls0CNzTf7NGHswJTIDgVv/r2PWV5KIy/l6QFJ9J+7A
oZwPr0orRwlNDQ+BmS+x3dbDfiP0lXD0yHRN+PYGF3ID3G9MmknjWgG/KPvrXaW0aD8CLJiSMAFR
X4VsywJq8T6YpPbjZm4rNK/9YEm51rTghCPAxjCT006XU4giD3iw3zouBXQWcbeUuxEbH34IuAYO
gl4OmlvuCEXue4QZy/EYwCHUlOXnlD/YMZN/D5Em5LvXZ3B1fgEni/nShK4hF+tjYXkYb8bUW+0M
O7lT7c9Kf3j8H6T1z9Ytny14SP0XzGJt+drG9L1WZ7S3SqY5tS7nDyaH5RUnv0JWXJ1IJDYU0CcJ
Knt9AnZRmfNmVhLySe+Puh5eGV7A9OkFbAHDyftDDVcT/fVbilqLeJFSDH6c1VLaUBQlzBGnUUjS
o1rjHhL/vuaB8Sn6zk36N51J8PkkNtaJcgZSDjVy+TJ5TifL55SWLUVAb2PClw7Iq3YCK0wdLTkn
fN++jMQI8E4Mz/5UeyfaRqGMA3MFd1afxNVO7znP+lNQ7QRfCBaiR/b/+1wu0DLz2kOxPklss/LC
sZdhAtH6INONikhsAh3FKuGlGSs3/cJtdTJLebCUGh/Mo9ANejm01a21lFHPP7tEk33ueReBuxjk
YbcMvHnpZa8TGVOEYIw5kT/ev8lOt3qbB+1haJL/JMsvopqrb+WsOCf19wTehwPw1fRCAO+LltbU
QSAa01bxgo6vR/QPHP3wD2vaa4o2RM7eeSYIws07oeQ3YVvpKgp1WUAiwNagmea8/mRAakf0YQNI
jHkeyhYLVjSzeBhWlDH6FaqhHOLB6hbDLzDkQzioFlJStTPvsihKENQ07PhIr8EZvbUhbd4rQr94
+8Mz0aV9nOTf4se1VDxh7p1mh2Va1Z0pmZnGeBlXMFkjboOPka4IJxQckYrXf3XxrROzWFpvQfzU
ciId9+5SBuXcbSDDu5x3DCOkeKZapU/ncmtLPNKM5JUFsv+XCYNg0hPRLBBUj75/gGFFvBr/F2g+
6xDe5KPbYVtI1ji+T8mlvqqDYt1u1uUrhoV0LN/nn+xOKo0xlrCiZCTehDbLGb1Ct4ir5ntJmT0J
gcuPjbhlAwyGSQI9gTqtSqvYauUSXSAHdI8o98Qw2Kc5oht2kKpl/ZQd42VNkCwk5zQZsqrJJ13Y
U7l0C3AnIdKUR1TzM3R9B85NInODO462R0zIzEFd06hLYoAZRV85kdrTlhkRrP90Y3vKm+yC/5ys
SF3lUn/kINeE5Mgf5KyVv4gy2cFsjyaO4/Jkzai65AxvdVk0Sa01CfKYjrytdQzH1OKmk8EzDup6
s/Tku4DHeGnk3pO7H/84s3njWnEuW3Z/EdKXWq77e9xvG+CiJQH3OWpK52jkK6CbhdjL93557WOz
TSl5GHr+eP082+OaqHo3+nY83oFGCzMIa0Gml2aQk5AtGxThxumxPu45iRGuvo+AsqysdLmju5QW
lRiuvJ6Mq5M4d5gFMd6KNJPFXBVtFOZadWsnd4fieGrL8rNgRB/y8zYfBs7WLlLI1c04memX4AWD
1j+9J0RLCqYpSSCAGxvF+xPQIQFXmOGW6rvpjYo2JroN7wGAmoYfRKYsA732u5RBPPXW+JbrcmJN
SM4tp+OzkIpU/IbJs1qFFlpmociTnIhOESFo2VuuqpLlB41AMikwzOJ+WilbbIgAwF81iDrHHSt2
GX1IcXSBwECWfdXh8r+B7L9qpJDae20bh8wNzxd9hFWQkrhkGRSvaEMBIpUAb+UZXUQrEe1wBweD
ViQcbHDyPQeFCz5WSwIZdlYoos7H4RgPvKoYS6CDIS+dLRLuFaMHE++GaQHu0kwazF+E9Y1yN4Cc
ScZNMXf7SFL4/hZI/Z/EfEwN2j48OsLSx0HDZ48BfBOednNVFNsINKCVEMrOrTqFPqPTt+51cgGd
GpUaGCcFMNrRUGET2LkzvwNb3qIKcGFL9roJoeh0QSg960oKL8k0/OnWtl5mdxFZENIDCZtHHg9f
PeQ0Zbx59FpFYQGTOxEwKnWe48IezMII63widzjUqQW+yCxC8p0LszbhgnH9K3GbUaS3jrxP6bzi
bbxHKyPneIWqT+ui41HZN4jqww19DSHVoCu9OCBjG5GEOKstHmD3jUftjjyfFHIWuLRQ18kT+ygB
ZgkmjDmnNiLTR2fbr7bd3qxSsRCjEXV3Ee+WwY2x059cOqMWl5JgAj8dXb3znE9eifsDW9hoRdsX
H3w0IPSVEYqKMkxlRkd8qzeFAhRklyODtCAqUecthuMAPkN3zx3IYa3X3wGqDfT6Mt3vINInpBLG
qE++gXa1+RwaQHl6942BByB7aEXiQVy+C5wXF2UFitzIt6JkPKwzjC7oG+XxCT7WnNqpZpTvZIiI
iIUa6RhqXe4WWz9h2G4GiMyFfenHghKwovEK2GIqVlxuHjQdVGcSwveEl7wDWnIvI2AqNplcO+Vl
mCP/S+r17oYBINWenfkDgwPMDW/By/Ricm7e5lQBzOzjy+rZpQ8yN/OyvFIs5npfJnE5IzhPua9q
rOHAqGdWS9X38vq6aL6zgVs4S7nGcyZlTBpvxUhEef1GoIIZ6ortSPwQ4LERrZiywb6pvVCvAsB6
1MkuF+sV5AdqzpKvc8ad9RIoTLaB59VNNjqHYq1WUb+x1uXW8KOTTU/IW3wlrzkVt0nJgOmAiMTQ
3rQ3p2cHLqkp0arf5q0z0Wm0Q3NuvOIZnIPxsCGDQNc3Hpa6RKdmB5dp+DRH2Y47Mwrpd+z2BsDc
3gcBfqOZqLyAOjZvyEa5AWqGry7C66FZ2bSJ5JfOV2xgfWV84ltMP3fjVEsqg3n38ewJolWDjowi
1gS3wg4GHhQjNaK//E1ivf6SPuthO+/Qy9MbmcYlvsO+Slly6xYuodNM/RG0zjhUitNUt0QoFz9l
qVsExiRs9RayvPoPHne5VRAzAQbMhYTtyABMuqPRwC09Loxv4LRklIz/TbRGVL2ca7zkVX9APXXO
DfKwwZ3lCzjqCfkr4UTI5T8iCHaK7wtvc3md7qkKrkqxNS+h+3iO7N7HFkev8xgFmI3hX6me/9oH
6TPl01HXeNWmHpzGB7jAMx4vgX7LDhzEJGhZV/iRZPSGxtP11uTvIK7hLvi/f9hXqFD7rihFYY9l
r+ttx4uXnVaGhU3W3nU398Uz3DkldUfmG3LpFTisyzN1goI/79C/CDUjpjVKHVBAjsKR858MArb+
Z4aONLr4W1dNLFaXVS4XLc/JAEbu7KwlMAwtZLLMtBBh8i+mkLMEK+or+zHPU8wTIaOOzVn2fEjj
SaM4eXrIJd4vCKnpoAIm/3Z7Tb0szh+K/dyv0i3pSVd271W7L47qTiW1KfqGhPMLwNSn6EPlE3FV
3olO/3p59r5w+ZxMl66ZksT+G8wAA0Kmk4YLkuYbcP4I9v7nXIBYaMjR4zO9052gT8EbTXsAc0TR
mnWon795WD+SW5vo9dNGJdm+PJ/JDIkjoAsrivwRYfGwUwcXA44AvIdJbkJCJMtuVUjD9r/oOepo
9cL6uRcuCo0OAtVXq/E6nkYKHLW11DfrXKw1x6PrdNjtZ1h1hd+7pf5UCcM9ED6JwSyzTUvtikrW
BDKFgpJL9kophG7chDSSPISHR1CLSEKST+aE3T+V3CXHkF1mVVA4dlLb7FJ1asqHDYfuT9j0oeyi
CBOYe76nt5qL7BVYZ2L3YZzmVlGTO1cqTcZ4Ynjh0aNd/L71Wa1ZX8lZr7EOQNQrqlJ9VkL5BO1u
qSSB+nqY/uRo0CHjwxfHnG9ihRieSdDP9avG0lz+Nb6fWCVu48QwGLSlsRGa4RVuRbWpuNIf12hP
JNDlFOTNKVhiTyAM4JSmKinxKq6DQUH26iaNLw9OpvOoNnTJY3TpcrvrTYH/xgFI8D3Ht/bYwdRJ
08SQdlpjuYD2aSVhbuKRdnOUOCnhJOPXN9mkeEBrqcd/X5GF/0ENBZOeJ6kx2ep7NzKjgEF4TB1O
mQFvv7OrRt1TCTQo7pCdDmGdBxSK+b1kIqCWY/BQPdTb06Qv67va8/BTJwaM7roPfdw3lTiME/LM
ny/i31j5wjmrKqkY15icKX4n5YLWsktn0uh6fOQGraI6Lz+P6a78QLd2hE7F+QBxAwT3qKCMcgO/
RnmgGKtrSU5HH6iHhRlzPl3EFrpvhjQOJD1GDWSpuJ3edcOSI2+OASpjhBv+dR2e8tooRjZaWUp2
/73AjKIX3Je15Vo0wkZQn0kya0IaAHihLNGqmdPJqj+JxaadHhI0kheqmSzBpf2eGuqumFwtAIy5
SrUMOYWrT659cmNFATxoOJQN0/4emCqXrUb5T/UbEEigmqAsVDvlKde5Rfd4EYHolkVq1WJMG1e3
aZOSdHyHPyvM5Mld5Tx4X/k/hv2nKinlJ92mhW23e48kVBJjcWssW1tzCdraD1wN7ic/lFIOpLFi
TfSOvv7J8qsqiKw4CliIX8rdvzS/iWfg4xjNSDVv/ZLcosUdMujWlp0dldO3/1kdDUSPWV7zYhXr
GbeGj38TQcOiygTQUM6oztehDxfCNYsa5ZK/cmEFf+i055fgZUfiBptjfzJrCpIRwz6ZBb+v2tRW
TWiOwHSM1QWZoP4opV7mnEJRXsPcHD2yA4+LPAn8VE7NomJB629oNAh7onKxy7Y8VSZKe2Gyj4/E
PTmWgBe/r6rAkXnqx/YiWz7bIcEuZcUscTBHz4UFF2RMokOQHnpw204mPHO2ZtblTR6LUx/0oGgs
fZSh0M3i+9aMbtz3rFb+ex/opdIa5d7WLA8MX0cIYrUbDr9YWT5Jmnxvk2KDK53m0FrfoEeHEq9C
fIBLyky59Wl053EjtAae8f7Z4qILOyeKBsSbmA8docJ5l33zKq4JJFmAaeRRmJdrCGitOOFVu9Ud
10Z067/JOCHKqU9ncpKQWfIszkz1nAG0LTvHPrAKe0AFxkISKYsLamX+rb0q9A15/7yWnT0yuLZ2
B09q1K7r88w/XRSbhVOJLTbQ81/bDWGDhMdFCBVitonGqVmSKQBQBbdbhpMyBDgv4IieRt9gZJxz
SUA/kIj4ND00DWv3MSSaDIZ2Fqw9YjA5WVDi2GD9nr7c2UON9CYkUZHRw1LEdB6D8wMid8y7Zod/
KmJMGOhn3Ez+ml6U0cqISWgHzvNMHxdIezPZtl4ZB6GOXPjo5zOeEe3SEbkhnJ5Ww4/vGr11UkEH
Tyi+/r4p97O/MmMhip8O/d0k4PuCBmBBH24RKlMArlBQZa11tkG75j6OpqloyS1BZjfA4uXIORUy
ukjY5X6mSNp0sO3T5Ca6F9LlduGaUTpdusKYtT2V8F0nD20izUTd9VSIDvqtp1WLzTQhDvLtbga+
1sLfeeIxSu+wFurB5IucRvC9X/N/1bQqJDT8+wem4Qy/vuaDNaD9fZnT8YU4qwjurkDnsKPePKPB
0SIsfH7zU7Fx2N4lpSTPfcPCTiKBNNzlo/BkM1WjZ1LVYQYCFR4DaJ3DcbsRjsAU6EmCXOV0JPCR
Mf923GnYwo0C5OJc4bZMwt+XIhuiVPrebquXixJtolb82Iv/pVcQ8zOq258XakZUY16ve5+7nM2Q
c1YVNbaa9wrGWVf5fe2zYziHEQQ6yMFsMOEpoFQh7qnCXC+sh72Xp8JQJjHTJxwN9hIgLfXPlIQV
fWL9v6IK5nHfkBWYCq8h5Sby+vhV3OlQGMb4OfNdZ/f+JYZSVceKlRnK6cHpKAyVgpq/7VOfhwZQ
3LFqZPDvIyd72SYruEeuPQvLdcEhcfhUHYgsVC7A3NhdBZ/od/Xv6SNxhNh2BpOo2eYIvelQ6RAh
HiTPu64J2y7ZLNSjpUxqzj3mr3ulEKP8IgkR6h9ReavaIyfLNpi1t6syztIJq5zIwB0VfIQESx7r
zE5uU1B3iDwWSvVkVXjwSm565FG0UUh7M8AxL5aQryBS3NfV6tbnB5KfFeLA5A6IEGv4xOIUiruK
wAvCZyrfJ2xrqM5c4+My09v9N/Wvce2WNL/ZFByh9kJElg9ho8kgQdbm7jFAJ8AWORkIYRY/YWCa
UiCuoLbFVk9zxxLV68qNogn70WnRvmpjoP+NJDCDpFPEMidvTNk6m3NdyZ9FEnzRe18YQI2bLRNc
dbos/CASmcZyPDgrtEwDNDHmzMOf7VtANcmRX8uhr6KWr4U7R9RNv2hETTMYJksVT6/zHSgfZ1WP
f2evD7Djp7DVgM6NG1RmZ9jRTP4ga+rlGuIA2/RBaeThJ5HnS38GG0jRrZrm/96Vz6mwOyQ7agtV
UI6FkKM52iPv8RmTnQusCzMk9XKNYfwzbpdpbGsG6IwWjegi7fvuu6NHm8w2oWI0iXP5WPYeBpBX
lFke+JJLLYtN9HG1SW15VdB71TTKijOo5sjcdUfUMCubPrC4espzmYKRFLRemHfwoHlX45586Aon
O9+DCQEUACSAZyLchMua4v/YMjr8RwE9oXYuhwxrYtsZ5q/o9iWqcm0dzlBgn8Y0ctiazh10SUou
EdBNyPhQLi9qIBYHBbHTNwmhxI5Un0onNEKQgkBIc9L5TxJwM/JMSnt8X5NwLphVfvx2tDDrYZbQ
+OaCFe65jNfZ6wSKFig3a9XGTsuB8/tVu7bINYV9RZNsCed+RC9tc1LHsFZKplp1hAmXIrqtmBAb
DygX3TqmjAcl09aSDPWDhteWdrJehc1gjn/4XMmGIOL+Nx0RwpKdUtW5RW7k187e9iIvTu1BiXUE
4ZiUmgdaHLItMNv8LrRE8ny4d81GYlrxNbAgH5dRcYIfGzJVsdDdsXxrFuNIrjSgZNco/dkqp2in
guSx+02gwo6dYbjRtG/ugf9Fpsh1w0KwCEotY16mKjUgKIyI0m5gpEoBuJs/tSOVVwQqHAPYdSce
OBB8zfbtT41//Rsgr20byJFrne9NfRYGE4UdjHaYnn439YDOEtRBG0a+u0FvaUgMevlIR9ekX3FI
KdpYnATx6qnlRb5V7DXsGc33WU66LoZmd6rmes49KHOPOYAHXqhXTfNz1wObHZ81peecfHq0hXRk
vHe9TqwO1TGLyRo4dbcngoGrRLSL/WLCPIIhcwCRyCMoACGS5q0UTlICoV+i6giwmGHCWncDSIsk
KuRHKWFUF61/Q4W1noTGi4mTSU6uwzYHdX2KN1dYPysJ+UtDpsd3OzQtcznMy98E3+AIRxywdu0d
5Mea5t6MgdJmv8vW/t9/5+6cxffEgzR5gOcwK2fqO+oimqHWzcK9AMtMegX13D+TzMNsMUIbp2n0
tTATYU6KOYGIYzdvMHbGWsELmdlHIecnZIIPPDqYz6KSWpM56g45l75vvE+b63O9MpEait00rHXs
B3b4yPzkDZxATaIDGn18Rz/lx74fSu36aTdr4OU5yP72SZMISyk7b6lQvPqTnP3Wg3LRHB3Mj35D
96rjeb+kEu4qj+GVt1NvKr5Day0U4sOdsKS0tXGeFg7+L93tzzSMj0BRGVJzAbSuV6t94nS/gmyz
p0s/uM/U4cIVoq0ObUuQrry6JNkiSY5f10WKYbmMu/kSL9FsJSZCKIoyBE9BKjHkos7LH2miWTxc
XhY0CbaqKC06De7qhjXPC3YoFNFeZ984/pSStsB4O2SlIVhL/63ZNOsL0Br22kunMTwy92TmxrGg
wSofkQzwRV8NO7CQk1MfSluSAXhrl+I2M2vLzHtXN3kceL9zbMSJEISnI1GdwtNtce4NLQTzAqWY
Wp2m38DkCuSU0l81jZ47mc9b1n9bguuS0vkJwCD6HG0moj2AFCOw/oGtVz9wOZbHB6Z2fOBx/mOt
CG/BA908xWU2NKtZqFNdYiqdvyWmTtpy+8UQCI2v9y50SDZxOCQxeMIx3NhfLofiq3SMJxeb7Rij
uTp9zyk+WoO87wCgaJuPNaT5xkNXCQwX2esYB8Jf1j7lhpbBB+LePa8BAnTsygnbc08BqOxvFYv0
dfVucpE4yBBi/jJRhGFKw8mEmVO0qzrHSwpDhz1zxz2JuhsvIE7Jw9aKq748lPmhPbVw46c7MnCJ
Kx4uqRyy4bN+NOluWR663MH2uUhwllfbQFjOdwGhXiey0xj/T0f2x/Sx5g4Y7wIZorJ3S7P9jCfz
gEdfWKgxb7+kAox1cxNQWXLW41thZQgY74XXW3rgqNIIL6Gi4lSzTw9Av1ngLUuxn54ahx5p7sVB
2YNRGC2plrZ6sRfBpzwcWLgSe6rVUBkxHK3TfTdjqe1rEyCcqWIgqLn3f0rtDipQVtdWmjJc7zKZ
YXpgob09Y4AG4xrAn9hAwsS+uA+dzXow3T57AntUR/NFyp6IG+xTLRFKxpUBn3LfV8H1yGF7+29s
9F7MSnEbKibBRAutL4ErnZKY7+kiIXQZkmfmGkQqcP2jv31WXkBIgL3/5cQX8+WpHUR6imqgvaAr
iRwLm8wCpDsOiANkARwXIUYekLHuI2xZuFGpOf9TcDrkkjftSIacvcDDfIRA6BUFNHfh/axy1skE
RZwaIWwQVVqe8YoyxyRiS8gQKhSFtNXr3piQI3wot67W3EZv3a+m9jSlEBzJtZGYvqgrhH/q9jJ8
gVFE+Mdum6Hr25+5xX4L421gh7JOlRQ49k/5rT7GeL/eHlriWUMjRNSMI4UGFscVDREQCYXhUcRi
4Owr5VE5JcryRD515v0tsFaMGLH5MuXzMjIYxXhADvp6ScOlJZgT1MGwkLr2eZU5J7O4KDZBQfvF
t72bFGO1AV9z/8oWcjcDaO7oZgIz8ZmR/WfvGlStYggWdwRZ1cMkWoGSEUOD/JDIRJZzTERxBIqn
qST4GwRBzMSGh6j1uWvdf3yCg7ivb/YrkzhIFneUdGqXJ7ed08Ab5rrAy9p3YPOz8gTpoCVIX/ci
why+Aqf2KRAywFuXnbEy80O7Rgl62mIH0EvElNzj34vRe6kUOZ3CpIpXNZBravUdE2ghzcSdkskZ
zboX8rsaUWc1H837VVGvU6qJa9gz+HBujRW7hqcwO79CLQBY+truEJx+9f5Tsr49JH1FE1id5F18
28J5Rk8eL/zUtGlNHvoIR0EOyU2XgCXd/ouQufOY8G6kELzbUfLvlUAAsm3WKO2Q53Dow06Se+II
Kgjc80QqFRx/0KCzHK5gwjoazEXMNhnLKDtk6zsuv45NDRzGIZb53S6SXXfSormfup9PR1mia+aL
AiH6XnvNwHsiKzjCvZiU+AuE1CQxENy4+zNopT84kfAd8YLBm2IiJBAAPVn79Awfcb910Q2KB+5e
B9vGGvqiZnKl2AdvGlJkRheqPWBFfSaS8OZUyMi4b9nlf0A5IUJ1l1TNtgNSRPt2jRqezyA6sCMj
9FV5xny1IwoHokkciAiZOCXU+dyv1ROBU7BGdutW4Wmxriy1TwXGuBQpne8THGAj2Vbz3LrAd2oA
yjYJAbPdNktrhWfWChsgXf50mSCVcBImSFXoKU2Z7GNCdbnyJ/DSnbOOGEPeIsoXaXsTg41H6gjA
ELO/MMcFwQ5CFK4cmS9Q2NFr85sAIVkjTM1YxE6NIeu+ovwZLgQp/i3K0hhD4wOVmhHcMp0xUQsC
/yQV72pE7UOrgQ6u/ZO9EiAYzsJV+rwDH9iq/VUO0/R95d/R8FsL81vpixCzNovZr9+yisZCiG9D
zNtkM3wfpAdmeuWwauFG1YbXzyMg8sZcG5fvtv9d93PJmqLbfZEkxUGk7MDfrA4Zu1BRBZOpNw2K
VxW4fDIX22uyqnLM8eHLbawwVsBh5GCVLO6Fr6ajFC7CxfGiUmUBurYLulwk+Yb49quR8CRkrloI
M5uSU8kflQxDqpP9g+eJWRTNjq1A4qBmx0ystARRrDMYBUlBeOIei0o6TmZtRSRUSAojhrxVuNxu
EEkIQfe6jBYFC0EHPN3XV49kiA8+rr9jw5cBHAfSTPr2lemskrVWZlFzcr3GFfTXt6clPptTvf1q
COabII8jhQHUKJvqEyYJ6rQPAsULzVpK9jURdqJ9hP9DDy2JQAeO6kd1flmHIormATJz7BK7RlvV
6IA6NNoS/OhGCF1M09jIutxC+98KoewedUnJcmeDNPRQ9qfmSu6CCGHYFjDi2yZOvjZoCFF1qMWn
iNCj2sjX+pEmbyMDa7yGvOLdMKObve27fo58nilhYRbK7kuZKYIvIISyd2RbMlwHnPG/+krn2UCy
wz4dRe/PfyNXHTWYyPEK/0sTMzBa2g8JQbJHF9CJMU0nk/BVxFfuH9T9VfuvsNYxM63D7FzEs178
ArBJPu+TGFyKQNBsw8ritb9igSeQ5RZ8vQc92xGHQtURB4I5VKZIQW7jP33+JBB2aePoOVhPETAj
G+DeKucA6rqO/XQj+uB89NrrjNyl2hA8sfwZXY/A5EhuaV0Kc2DAqi/o++NiszFvk5KC8pH6jyDo
QAULH7aT3Of1zGN7uFMnyU6oBM4KF3s5aS5wworDN4rQtu+PZNsL7e+6IQY99i6gU2MG/yhPicpI
9RmGz+tkqC8WYar9XGxbw2EM7zUh35UQJ+XGRZ7ed5EDaK9/HLj2b6r5R9SwzDRf091hsXtZhesn
UamMUsu1ha+rGSWg5tz3tGkHiH1YPtIDYxPF4VK8cWdPCpl3jmyAv4S46fersXGZCDwuVd2Gu4ZK
40zbdQd5tbch8vEP1yZo0doXp3awQQaEVcPUNt4+VRhvVPPxYj1kLzm+51mD7BS+KyxvaV4GjxGv
tgY8a1PKNd2GqJm48etibCcirmC2tqwtUv5+7q4vzv1iyP67hubOEh+epGGbBm1snDhAXg2QDSJ1
gagEvCMtCVUb3b7+G9b8QlK4ECmDyoAAhtvOqlXYKsckUIt1DEm+SBNrG6EOYfBDAJHQY8w+BbEi
ONGrG+Rzkoi/oKaKWbImoR2eDHXolj3f8U6on2SdWGxxDg16OdsiE7qwtYmHvyP9yC6rQ2QTDV+P
n6mcdeOHY2BJcoDXr/NSm9bYZN/uUYA0/TddAqnY3eg4f1iyBJElAPzaVOtrLD98KU8ja8L9Uy88
/OuJ4NztBcO0D7BBil4rkMmQnE6MJQ0R9lvt+rXFVBrjWC7k0QIjQ6ipznX9hhE7fGlNjHwEkbjI
nKflipTFelHdJOw2aypDFPJFvTCPyB2XWSg9aqQriR4RTc9ydAkFgBQMlEI5s9gdiSCryHOaeqDp
BI2q8MP8SmWFPKu1fppu16Rh/PDH9qjURFg5nxUfvT0cEUXb2ivh90lGHv/saC9RWe/rsgtYMZPm
4grjhPwNP+svg/+v4BnLJnYFW9xP2P9VC7uCHCzCC2oxUQ7cfxK4MDZ8du6emHZTLF5lJf8dkZ+o
hvysIY/1KwkfW1clEmGFUdUmfG5/CE0xFpADcCzgF1wevIK5OqAvXFY+hM2wcIin9DEPPx6VWZQF
39OwOG9DxFelwALzjzTDGxXWgCmmKDhyRMpVwtMciNxJ575rIxcreKf1+ibtYDErr5ehvTXtf1Az
sNiVOi5lxJE9AB/opWR65G+CGoPdvW8MP2cLftd2+3JOxLlYfhroRekAAdczHWh1pB+G00e9jQC6
nUShtzUjgA5euuUj2VDYxL92OqRLfhAH2IKCfx694Tfa2ixqsmjdQxntvDtSkq8OfsRLlLTlMqaS
hoKbjaS2DISlTqAtUlnHpBQ7bLB+W3NCajrdQ16QNW5XoKxTlSYrL2ptNf2ZOhCYHlt2eFRMDAh5
3YMw/EO73WKh4IdTfd/trsj9GpysEcXhbQUODLgLfCtUkio6rm4pAA3iQLLNNUrCOWX88WxTkEN7
3dNX//0YycUiy+Ra8s5Z+JakxKyj+FPGdacJO68r2Z1VPxM9t9QuMo3Izke9o5t2N4WgbiBd77e9
EVsnDcSuj2kkcTa5YYdIMacqUHGPKbtm150iXUxZcPi118jH/6IRQxrx5gtxAEc+Q21i9qBwVw0m
Y9m97vNpr+qJmjThah+5wXPbtpkhWKipZRna2+unIZmsvpNW1wTNjlFCmQ/137c4iKc/e39aJDR4
eFJ9KQuE0FyihP7mjNwm6gxKAqW7Ny/SNlZCQOUVhgy0ylnN8/F4NS9JovcEhjuO9RBDx3ZhiMwy
S3uVjMfsziKheGFWGr9XXXgamiAclrRWxWta4eRWKOiMVqWCTcCTC+6Hh8RswH++uqcSVP50ntZs
ptrnm6rcangquwG0KMmgl7iH25Dz2ZDExq8gWUZ/GwcZ55hYQO7URvFqMJY4S3jhX4woCpEGzbC0
rbP4wqgZm44iQYIhxm0oI8cciZ2omCDylWb1DevQUPHsYa+g6gThzOzEVi8oj0QvOS4YLOIN0Cbf
F9jyORvBe8oP0FzmxdEpLBjm+a6FI6FjTG/TC7FIaicvJrxxan6vhpZ+D49oTsNwNzoLKQjiTdxZ
xU682ZzA95hH4hAX5+AzOy3OmqqzVS78lHkedcL9hyAx7+FeYYWutMb+pnN5qS9O1n3HJuvfrTTF
SNeSDWtluIET9NvnCC5e3dmpA6v1AzEnpS8hCaEN415aZAyDEbwr8XU8qDwlAXbdDmJ71LYxU3+4
Dme5QtTKHpacDLfjesRQt+0N8ioORQCSxfH//p0WteKWGMI1zk2UC3nGOqsVXWcyCc2Db1fbKh7Z
gwALRwYgOmuukNyUlsKaOAyZqi7vX8NnI5jROSDxqdukq3WBWie0GdqnJqx82hMX4qhrSwkwfK/E
qUnuXCOCjMDrch/wJc3IEDiLlJg8TaFwzl3ha0jqx7Ff02Ece8U6qfHY7n4pUNUN8UTnKD02Ailk
gN3FboicaQILw1FyD7FWjANJ9OIwuZ17If4ehGznexg2pgGn/QkwZhM2Nt7IT6ng9dRJAUCS8Qwq
PBPXeKNFLtHRPvayqEGl2EqzhSG8aYX7d6bk6QYKR8JJVtGQkgjVlkOtYq42rim7ZfVEFFZZJP+U
N8c22rDbmLuudDDD9GNjc2nNEeER9qneWDPJJfDJqx7EEbMNLDUtPVD0L5NdIw6He7mwD9H73BQO
XFdHNpDbPVqXeunGt6UP3wEFTdQIi6WIyCIP+P2lhMtA//3vmgvif1BDlrGAAoKNbWxdhAIPDwrw
6L/5d1zCWoUDoepyykgXwvT+yy79/+6Dtj5IQUj5aEMKQI9nnlbHYIEjUSIH2eRUu8SdVYUbw8xE
/t59jv8y7rChE3Ch6jIm/iAyQ62R+Ib4Jjj7aoZVoeyWl12sSGzsccIPoKbrA2KAuJ1BM0VUT1mh
8ozHTWwHFZ9VsR42rM/ADL8CVbPIdfele03yTPCHk+U0Gapdb5A/U9YdjhSKwQJZlGHRr/dhz21n
PS+Y2cIZkzzVb+CUndajN7tlVOR/SGT2lbWQlzbTUZd4SEoXkcXrrV693gwfdF0tYCCkA1e6Dl71
BSKONHEsj1q/d7Y4kH8H0gYgdup76GufovsNlAJYJu6b3TfQCcbcBUfcq98piLZbkKu2gZgO7Ybk
oQtBbKlTFk8SDXl9OI+I3yJurIwrBFqdYQ9QvvOmn+XzP2pGel43WIr0jdUDAHrdkzQQ5PepTbwP
x30aPra6/31A/VY5uL6JtfAH7HOUrNxnWxIzb9QwXLhcYdos94xMOzmYsY6v0AWYsXo4O81KEVPw
l5nJNL3PyH1eoSaWKdhYYfd6BogwWzqfBSfod7oK0tNclP4EIQ3Ya85ye/wrxU7wKCtpLVPQvt2A
K0bCJwGwyzIvykC6b4kY47SG5MUKPkXpCzw5LiccolVluQFM5H3CwdPWwQsrTouhaLANVvMPDxct
P2oAPjZcxaFi0mGAusFjtIRG96ERuMYDVM3rm9ctZTaNF/amBJ7RxlT6tFi6Bpb+9qvEteLympFr
f2tBWAtJvgRutPycLhbgMS/Q2swDqWBB/XcSp2ww6jPYxMjMkzIFi0p7slBObhBDyL4+dd+BWDyl
k4kmJPSe+yXmbLAGCec+2cQC5yVqiOhwl+zgEfqQ5pdfxQGzqGt9yTdwrrJs5R9b3F5TbDCFfEIG
Xdg8X4yS0M3KhPfie5xK40/WSeh5bFmW/CHzR4syCGNPdzz0YmjxfBQZ8Lrs5GqieLRPy1+t9u6w
Im0cJYReb5XJAckcrRNLC9J/vh0K3qyjQERTjZ346xKJWjLHb/SCDA+chX6alJISmJy9BM4iMf9J
6/SxntXCr9j7HtBYn0lbHx013H8xrVBqz9o4VeWG22qh4risXZSqjEIp8T0vMIqV1K8Fc6dmYti3
9n3eInVm48zKsKy6gPQd9C6O7gVC4nGxbQZqxVmMvV8cgssW8Qx29R66w4P7JT2i9hMmPtxxx74D
SXXYZp6UBRKalNednKBmrd5NhvnVZ17IPaZbMENE3tyG/odNHHVrdXytQPapoldjt7iYyVeZ8Jca
RU/bAZS7TQOwxV0t9NqN64mE0aTYga9mOVVkwq6Yjje/deAuFsyy69xTfAfuHWQbWz2YqRRjaxMe
PQS3qNS1OUsXp6Fot7TWZroXY5pUqIFOBttGacQBY+EpyuOwUA2ESH3IllN8u7xHxUWHnUE8eBup
qt0fznGFTBpF3iY3eevZ6MfkQMFDg9YQkWFiW4tyrK6tSGUTeA4gryJaGvfvOylO+keLCMegx6dO
56CPJLNGVmnTDb64R7gSfovU+nafLz5NaBnliWtkAeozSaWbiwCoWiMpJKC46hwXMiWMQ5cR1Xxa
04NtK4kb87KtYTSXNjRyfVwDS2j0M+1+3TAlpGBEERVYuKQpnIIJdspiuMLnG1H+pX3HPxlcyHbl
WpZLiITo15oZXTjeyeowZqxyn0V5i8gFsMXG9B/yV7gB/GcmKhaVnpf4zEBtZoy5lJsW63bv1qLd
TRHDbm6Y/7MKT0Ouvc8LQ4RScrx/FoCIRzXUJrfKacZDRHxgxxsrVhtfBzWOkPU3LM6aZuiQJ0L6
27RaWhhxeR0mFNKI9XspBQmD/7qzpck8OfP1a3iFPc52wylZCGlEtcNT+idvz2MBzUFP3z0i2dxQ
/H0oVJQFVboJrLZfKFufNzuyWk4y7Ym3kv1sptFqfVL8CAZNwIQ5AUyZyoV4tsbLuE5SvsGa8gtL
81pxEkRdwPupKKMBg+f+qcHLUwkj/TEMlUvmOzkUL9WfPOZS3PQimbZgWzbwHdr4kN59H8Mx6B1t
u9CYN5k6ko+5DiTiusf0FYiE60g/ctxV9Tl2KOQRsXv7qiptI155CQ1SZTeUiMOIUdL+pj3v89yC
IIa7zpFLwtR3PwhpjrzlDJOzSR1R3yeb8V6Nt6SD848fB4QbafhRHSBvRgwyh+EyhPSmdTJLvj9Y
YvychSBsLQlNSWndhyvUFBeSuDJo8IY4tlkLOJZvP71PbG3ONflBJX42iqtR4HBdoJWueWQMVJK5
HIdN2j45U7CHPfmKt4VCL44hRD1kvMpcIbQfOobkWMQ2f7fcokP8/QsXuCASI1kUs+mecFp4esUr
/cznErMUwX+gfiwmM7IjREqvKxoB2NAE6oyqBqQJs34U/QNSkiwLv+VzyfvrtHJnWz343Ry4rln2
DU+XePHwsWWiWHiM+DVY1ntF0JFzEF4ZPcPdmq7pildC8FnzjA5nCqY2XlJ0XcwQxBB604ivO87k
r6twLgrQ2DppiSlzSTU3S+9b/vOshsNN8SFr3wPs43KxJzRhrZwwxw24njXMLafCue/VHzSLHRGM
+n1MmDw0Td5prpFNjDmqXXAZGtEl3alWkyJFNXtuwIKFmIFJ9TK5Cja0ncVAjfMRCXx0Kh055248
EX2sh53YNxjFXEn71rlg7L4OoINVJ2ALG/WhOYNAQmvlP1SJS5oScln1OUhCMaY/Rp0kF3ZpV55B
tfGTyfIXcf0lpwerW/L8P4dFpek0RQdU2PPK0vwWsJv2A0AoutRBOVIPjwOXQFETTYrUxdpmRxwP
9oL4gAia5eTvgWFkjXHZMHx3fvsRkXPj22G9Gaf9Nc/v4JILcuigUhUUgOel+G0pZPmqKedN+jzk
jkZhXYKahYtmauqLvYKCHmEwY40UuFpThLB/NNY5ihhQoYj2Bpj6R5FHOw7nnIEdMfwURbzJY2iT
M+HdfTuaLxXuDsgH9yWRqJ5+coDaF7myVS/C5MBzAaswrspYlJN0UvIj2QpZggFvTS4BEXP7BoN4
Fbjbb/weQrzi/cd1kDtKRs4kJnreaBojHAxWKegyngVspW9C0J9tovKs0pbPziKJoomCs2rZZ6sB
1iiNkPnoV3e3K8myrerjmDRRY8pg9TRU8yJU6i9026KIid7t688PTnb9DzVBwwu34Rn3jrOCE1xJ
AKfKlEuOqRIsxZ16SgCQgWI0KM+0E/8SXKFy+M/5zQa9eft7mKg54wFs2OYuZGtH7bvQHMjMYvZW
wWi1A04Pj2H+qbDMLePq4fjnFseFrKN0U7+xMq4/FZoWL3IyTEj/J/j+MnqFzDTPs6qt1hvRK1uA
PYatNLtU6KXqvg75NtzMTpOc/cyjm2r87q1qLnEBOXCO0RmgdypAaml/P65SiH0uLO5nD3RVjoN4
t9X9P9ZhLnebYBh9GIR6yF2xQ+F5Kp3TNgtT5EA/RQCEaOG7LAknt0QuO6nnkYjZuXSUZ7gVPioP
DEa7+ZriZVTcXbSXHDGEQl9uKcy6PxR1F+rF5NavOiSPve5VWXL5/gu0Kgq/B8jAMXLa/xdmLysF
l+dsB+pbaRlsK6IB4z9rLGLwAOwpTaWIvpesLGUvDfnlEP833qmbnHAfPBu00YvSng6KgvHfXNid
wMIrLvcBtGzrck2cq7jLg56lI/KdIUbw8XQcNVlBYr9+0VAJewvGZFb/i5UO/j4mKokPkMs4Da1r
bBLJBlq909sHIpCePTu5wcsyJxVlqEJQCfqyFFFj6HnIZ0zwS0WXq2bi84M9rhahSxdqptaA3yKc
ypmB5ABuguHcRlCBHhoFPkgVkqcj0RzOqA4dbooVY8GCgWtfx5ZZCvAQb9vVxeYxnjbHy3UZomL1
VNe36JyMEoozALg9kNKuDzdPNmaMuyHl4+F2JoEhyihfH39bbm/T4kH1mJW9J6lntWudv+jvcJRc
qY4zP6HIuEtmgBiteBs29Ifpv/Jt6K5DSX2vxau5zKsKjayptMSD6luYPL/Ru+QRhRo/OC7UD0c1
RBCDlTvopA6vvKDdarXQHDFQW5xrI5YyBCMqIiAU24BYRnxT9TTm7jdPWdyqSbQecciuGICeH5KA
lxDIuyzljaRBPU4t5jRxy4+Q1FhmqowP8nZVXzxfh/0dcAQuS5HUTWz+0MYMGb5Jmv6OhX5dsrnl
wyrZq9WJNqSPnY00gibw7XCsP2x/TLTE1OmzaPVJ53LeNyL7+YYP6GdA6mlV0kF/xsLsdShb02nC
q9nRRnQYms4uTbnp1wdzrcgIVeQ8YDhZsW/0nHPiG3cdRv8SX8gsy+MtnfrfLkBjOGPUHK7YZSZu
K4zGvSb1Q2hK9dbIkd8gjeaUaxspe2ozp0H0DwuEkL2bpIrDWXMx+X1hsAAroGmou6KgonGhs1vE
1keKETWkoaL92TdEurPiFLHnZUaSVOjS0tcMOyNDCN8/sk1r0tbmH4i+JU5cwC7By0lXPgWYW2Ws
t9e/2JR8U2dSqquIueUpJ9QV3zhmA09RX3VRd4ursfnaaqfOV5a/1xJ3Aag9EnDn6zXasw0eTsGR
2MrePnIYtWic4L3qRfFUWr9gn8cZLQm0HJ5jCfAX/a+kDzwpH/kPAySrLHkL3Zg7u9uRhnDlirSk
h0yednyL9d05faawU3BbJcGrfI6FIXGWiMgOy9ZxLzgjvZJ3LkXTLFWDcYCbJoQuA593ZYh3Cg/A
3Rh84ORieCGpRO25UiU0O7TkibS1UrSNEOBbEKLVbukq/LP7s8EtD246In5h4b96Dqx0G1QUneg9
Jdk11GJuK7bzpDYRts4w6Skl+CVRwJTEZU7fb0IGeozCGlyYipV825adPhYAbv2iU0MuiakV0TxJ
C8RigpPUrus+XQcta3ZBrGdL2GJdpWLgemIjdhY6S5OqRtNC/zekPp8tE+TGOzgg1YbTMEpG3wvG
5rGjglfcmmOlFJTW60fd6D7tnkwk3649WDqt9gBGcvSxNaFqPjQ3fpWhsnDS2Y5bchq/QKsD0sJn
OaC7l3oxgoBpYMmvPuTnoHfxrYQrLMYXjjf9RFEna8J8S5P4MfzUPSrjWqjyRTsghEJUM6wKEmkg
2sAOPbZVDlgviJ6c7XRYRK61zLVXsP+aFnv5nx0Z4GjTxN9H0v7gb+dggnemricZVlVAoO3uhhKj
VlABRL2n0wNJMgLr0dsTDtntcdOq9WfMpKPmK8C+OAi1WUzmY3ah3AGujA06+0Y+RDlSlYD3mVog
BZsigLsB8vIzw+SW082Zkt+fouXpw+o6fLpXjBjDaHTII4r5RmKIiaJrxVEVy04Fl/j9dCG5Zxk8
9D2yi/JKklanfHJwJZPhAuZ1nBv/UPVizMQGBTkweggshACc2GY8phgC3joFTKoaghLCX1cAr0t/
tYmP//mOzmLv5Kb+TmiRxFNLtW+qnPemV3sEeJaraVfl5sH+CjSwDDrIMy94of+Qcn213eO7uwKb
vIO/eV93z1GJyFezcma04dagSQXn2lZY9fI/SKyqtUVMHp0kzoQC25VK0t4ByB7yfg0g6wfklsB2
e7afuSSfNceL3S66KF+HUqsljugZv/YG2LfvpbEZJv0QRZXog2AGOIQ1UndfWBGve+nnqA6MplYi
GjK6V9UZ6BqwB9mMAf13UWLNSfPfFxFKB7etyI95YAFpPa2hVY53JaV8WK6MbUAm6xthaiZJoaMV
izmldaZEUGQnm+Vt3inyqCOg7Tx/ekG33il5U3d/xV/yVBwMj++B5tH8vprQrh6+gPS8gqFBc6+8
bx2XVOl25n2Dpy3/hYIfzHM47zRwjUugdd3cdaBhcUCKyVlIYpou8Huro1Ad3s1GUCN5WZPzV2Ak
vlfVnO7GJcnsJVDK0cw3v32C5f5Rqn9Nz8g0bHRzuZ6haO5ucjRJueBfexUH/2aDoJJbthjic/xg
DQX3sDUwBUTsFCVMRJRXMmO70D67tJeMIkfI9zcR6VUG1I2muh8XIIMm9+cZhqc5PwYlPunOdNGf
UP0GGx8leAL4E9e9Jj9gJ/pU7XoWVP0RpklPXdzh1RdXDoHjS6/A47ari+KUVNPj3RSpwXo86z62
C6fV6f72gube7+Uz/OmftPEhSqQHR4nu/E8panAILf8Uv19iE9gLm1hiI0RpK40oCNHKb15ahUc+
/QIrWY8Q7/CZFvhqu2y0+BIi6CWtb3T5W/KoF3MtbsjxLMfctPSWHY4qK+mvw2lx4lXG0MlNaRP+
JgDp02KXjyjB2HScjyNYUvuECmG8GURKAZ8JwVLx6UbK6k1Lh0gM82xZjeL+NjYA9J7O4wywyqBY
ljFbGe808bJ9NM4U5nJTqkPV232bPkZHdDc0IivchYQQNAgssnph5G7IsQ7CY6XfzbtfLGygi+l2
FjZ63Ic9/5B7IT1ADVVXIyaiTJ5dNyWD9J5NZ/JuCnKsjoaXIYCxaqo50lWUax+2LFjD8HWkwVHH
LTpsYA/GVNB2JZocbYXhnoDJHst41eOdoDr5CXueMPicZNZcr2ta2ORvRrxjiONv4Z0d/4su9oMi
dxR7aLxBQAG+VNaVZOPf1SQIPKkW0yyUFjgk90STpJwSRuxHaFZjBFPUr3aHq0EdMJnV7NGDTPxY
CLg/3l/QSziyh/VzpbN9LZqYF47gLBWeisyMTOzQNB9E+VWmBR7mbNRzP8fVQJmcafUl8oD0D8It
SZo/cf8CFgLoJWBApqmSON2/0neO4Co3Sz3r+JlAZmXq2b0/wJiMcb6dKJYchMZC2vUFKyKcJQcm
pw3r68b+qLEADvasS5LYfLwVESV7I9Ys7PfiQkFTtsJR3FxzgVDHrT/MyYFzNIpRSYPJoo6PG1sZ
4u/Qem9LeuL1xXXA0mdwvyIV3wwHL8jP8tUlN9+SM3FOku9cc+TWZG/3wFGyt+YcsE8C4y5NbDT3
rfG0HpV+0edvNkw5xk8Dsh1SrdpnFUeTXjDJOloFV9UGvs8u2wYqTKrWIIJmb7Zgtc/IuVhwQl4b
WFVhuPV1EottXdQ76ge/yMfv5AMVvtFY9gz6h7vg93rd97e26ttoW2qMNpPoNAWdNMBLIPwjNYaV
tgexcEJgL1embk4UMz9o61l/JaS/HRhCh8w0uEETf8UVCHd7uBbbS8MU7TBZqxkABzHzFAHyDqRT
FSNWCCpfxJpGlKE9C1LlyKvFiW2merqq2PlnJbWGV9x8N9ZfG3hZ1X79mOG0pxZtgAFSN99QmLmd
05Z9LrEBnuFhepqZfLRr91w4vIAgoKYAf14Dy9kvFK0c9/cVSbxEeT+aUGlUpqEgSAnbq8RhIdCW
yo0W2pLBgdvUi0zpz/AgzPp40r121vaW/MxyO6+fSd0++gLBGhrwKH02U2c2vW/JGRx5RLUGgfFt
xCoaPU8142FnPFbz5y7DjcNJxBWjemdCzvD8bNlqKvLLQ0mmmxmXJI15gNVGLaKaOo0gE7yiNnXU
0TUNSaSCJLSxG2XYeS/ZwJM5QkFXJvqBBVNgkm+WEZyzwq7HvIn0gn6xrTcY4jmDlHK+BYgpiG5x
s+mEDLOfp4vSV69aSglS0bMSQ/dud+pjiIt+7+txt5BbTAeczMwWp5H7XLsZ2kxiWl4nvH7a6lXO
sXL1fXx4Bc+C95qcStbvRNXFpBwCpjFDyRLBbU900Ipm17exH+v/PH8nBasIInEgUr6uSJUa/JAP
APaWrO5iLdRRxYA6GFhRnT1lx8TEmg28t3LW3Y6TXaTVsuFqgN2rRfDW1MaY82LDJ6TyNQEgcLy1
k3tIILxG3fxlVyNfmuz55F3MMKkxsq819NY0hUwjwBjWP/jYMtp0/2p5asL4zm3pLAjgETYlMMYm
x/h8pTSpXGwLyBEPG+iJYhUbYu2an8s40+3CMAjuSuhaOf3CsnK5Qa040ThW5FR7BGDYiW9fEkVt
N72LUVP5YpiTV2GhPPxZrHJ3s/z29bAgEdPrvlP3yKkgq93ZFjie7xEyb6e6yUdqMdDEyzT61DB/
thwEQB858AZwsfifdhB/MMRirqYXG/GzpmFJpCWL3+oazr/TbxvMUFJ3pg6NJE4NjSpxcgcGwE6l
3IVm1jSOdg4lwN3G7JQOojlpr669OV1V0YsJ63+geRDTPXoHiOGnAL1/fRDMyNsZjZonzYM3tcko
zTsDUqjywUK2wrEdHS4l08nQhmqDTOrRqt5WhzhTTmLmgosAjB3MNU5066B3FWFvkQZGLoyfyRK7
m41jytHorg8McmoseeA9VfZO3WU/JgD0FZ65brA9W3SecT+J4GcYcSvBNuYcqaN4QsJ4WSP5H3Ei
KAOpWVDCfB+3KutcmemvinSwAfDo9ay9siZQcycJQRfW0apvLeu9dSn5P3MO+sAhPeCaHtijGGEU
gLKu7rgu0AWaiXRW5KjpDtCzyHUcnV44zAnUjQB5T/G9G9axlvCrJL0BfrzMrIozwHWEwicEc7G9
oz9VSNenXeyxBw+EVMwjxpvcgXPrFG0ZjLdOMrH5nqLk0gOY27caILq67Q3rXmiI6MQE4fmSFTVK
OIxAjpWl/1qoMLUQCfZ4XpKj6EdzWzWd2IU09WpD0cPpnraGHdIJLlahOO1M701SjyYENAQpg54g
ve4a1QChGD00trTG1EmCUjTIt4//NF8UJyaFXc3o/S8h5G8Q0kik/oetEeaeUX69pKRKToTlFGYU
ZG5rOa4OhBObpxq62MNH6Pa7sa9Hf86/rxpzZ8Ylw138k4DZ3pgQNAGQrvR+gPxQuTMlT/tVw6eJ
H1Rj5E9H9MRZgmaQv5XKZqyW887gcXhTovQy7yIVnaIOJTWb6YLO1p0upXlEEeBu803VZc4gDomN
vAF/VjZt4Is2ibdjlWi4F/sH5Ek8t0WDDXGq/v90lmZ6wey5h0HiK2and3ooQB7LR29p0CD3gERz
jg3e6FeEbk7MAyKtPJDnwshteF4oNmntsudgvqxii7hNHqONjkRMplC/EKEuN632kNQ6XSlaD72/
lKGXRBuw0dvL/9f65OhYnh+rcqUFWPVjmgY7yUzWcQS06JhrTYn1NiimRARVsh5qKKlBNzBEN2tw
7nco5E+Y3jMTHQwW+9geHG7ZoJ774vxvZKBEF+STWGJgI78Os6IJ3nrp+MyPvSXGr/bIhwd0lAND
rUFbRZHVkHRIuXNAdbKCYWn8zAffojrm6DPosLZ+cyDcPLTaAKmI2NNGQ46OpQKLEQWEInvyU/1A
kfzPISN28VVdz5QrpQAgtMWNQUiJMW8bibV2j6BiTvBRQbipxHHL0RhFAhBOl+1XF7J2hjdIpBCq
e0ln20KGzZx6yMgbE9tLmcd8btVB44DyuOkPnKCaqyvs7YirSEwFqBzgWgxmBK3vZF1Pbd9TR4bv
NRal0KSeEedX5V37DEBA96+nlE3fOunKMQ5xkDFjD8Qne74FG7hw8EWS7YdZ/lkQXidcZcDV7ulv
cDt/YySS8OYUrvVptYUnxCenGIXIpKdPMlhc9KVyja7XazuZTZVBOPZ5lC5Oi4lh+GJ4HB/vWUfA
yjtfWAWDrog0mr2FVaIW5FiQknMCXobwdflVlQEfjjJ6doJ0q1CRiMbLbZ2gZdWie+0YYAu82Jsf
87bhIjje4hyxBkCQ1bHdI/8IUYeywUJFjcmiuKp1jTXkuz8yiTdPNMnIHohj7j2SmfmiWMzz7GTB
QxoOTX+IXDrSB0FYH0dDop6dxPyae4YYapVdmUCnXZrpmxCEFUqkUQcq3jVRZidxXNrsu6anIczp
6pvH5Jf9fybz8RmR+YNGxnoE/LbxVh2i0irl7W9iflYvMzlQe3e1BvGHzpdDW31ENcnZb8MuLMcI
NIR219phd0dWUMqc+QDvVt+t759bjkOD67/GS0Khkvs7Ll/wcn6G7M5l4yP0Dvr3SJwumZM4rZHl
EW/qTjG+KuWEZqNor2+FgZ0Ox+cvjgmIUlfV9fxEhQ++yYB1j1q8vsvYKcTe6TJnLhozBDJG63og
KLpBCTs9dlRASPwVOReiipoxwlaIrwKS0Vlx9/tUX50GEaJvf6d3WqRFFAV18QwOjD1ICL9k/DlU
V7qfaetJ7uwtDGWcTTPx9oR1R3/cS3EN4EXerM/XiDnXHP9NZPKZwzBIh6G5cqd+XFJ78VAQF8rS
8dLYJsAlDKt1O3aqvg1S9F+qCrhp5BxDWofNtDE7i6DqHGL2EoDdAceYskcTyYJnMoJBPrGDXLd3
AzH+XNTJeqs1exxbIdC0cwDwBDrlS80xaiKLfTPh7irxzcDxLhTZ2tJrW1diuOLuUiO+0/RK+Bi8
5dPHvLd/xgZ97d7LU2Tmxh7e6gMMj9E7Il3VqfWGAyO2qmXldFELJJgAXoVJSoFcfNCnyAlc9UA0
mRPmcWqQA5+V4jDIV7oXKznWDS/KahrYgC9+/ykxoBZBO/sDiWJSkiCiPAJDZ9Qbedfmwaw3RAr7
J7EJT5FIQmJJZoqZGZ8xavHmXr4x/a4tIIUENbAODpXfsfsT6AnraiJQ3hQdAwfC5b0iCQlKYmcW
798TQ41WcTTvV+N9LFsUYUxuWVZ9myuBj44smA7loHIUhiLpzuQEVflyuUptzQ0eV7MRiBpSWKxc
WVpHU3e9mPUDONV2ZOEmThE7u155H9t/n5A+Bw==
`protect end_protected
